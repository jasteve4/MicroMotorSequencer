magic
tech sky130B
magscale 1 2
timestamp 1662496270
<< metal1 >>
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 72970 700992 72976 701004
rect 8168 700964 72976 700992
rect 8168 700952 8174 700964
rect 72970 700952 72976 700964
rect 73028 700952 73034 701004
rect 397454 700952 397460 701004
rect 397512 700992 397518 701004
rect 462314 700992 462320 701004
rect 397512 700964 462320 700992
rect 397512 700952 397518 700964
rect 462314 700952 462320 700964
rect 462372 700992 462378 701004
rect 463602 700992 463608 701004
rect 462372 700964 463608 700992
rect 462372 700952 462378 700964
rect 463602 700952 463608 700964
rect 463660 700952 463666 701004
rect 22002 700340 22008 700392
rect 22060 700380 22066 700392
rect 89162 700380 89168 700392
rect 22060 700352 89168 700380
rect 22060 700340 22066 700352
rect 89162 700340 89168 700352
rect 89220 700340 89226 700392
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 198734 700380 198740 700392
rect 137888 700352 198740 700380
rect 137888 700340 137894 700352
rect 198734 700340 198740 700352
rect 198792 700340 198798 700392
rect 22186 700272 22192 700324
rect 22244 700312 22250 700324
rect 154114 700312 154120 700324
rect 22244 700284 154120 700312
rect 22244 700272 22250 700284
rect 154114 700272 154120 700284
rect 154172 700272 154178 700324
rect 302234 700272 302240 700324
rect 302292 700312 302298 700324
rect 413646 700312 413652 700324
rect 302292 700284 413652 700312
rect 302292 700272 302298 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 463602 700272 463608 700324
rect 463660 700312 463666 700324
rect 485774 700312 485780 700324
rect 463660 700284 485780 700312
rect 463660 700272 463666 700284
rect 485774 700272 485780 700284
rect 485832 700272 485838 700324
rect 198734 699796 198740 699848
rect 198792 699836 198798 699848
rect 200022 699836 200028 699848
rect 198792 699808 200028 699836
rect 198792 699796 198798 699808
rect 200022 699796 200028 699808
rect 200080 699836 200086 699848
rect 202782 699836 202788 699848
rect 200080 699808 202788 699836
rect 200080 699796 200086 699808
rect 202782 699796 202788 699808
rect 202840 699796 202846 699848
rect 22094 699660 22100 699712
rect 22152 699700 22158 699712
rect 24302 699700 24308 699712
rect 22152 699672 24308 699700
rect 22152 699660 22158 699672
rect 24302 699660 24308 699672
rect 24360 699660 24366 699712
rect 527174 697552 527180 697604
rect 527232 697592 527238 697604
rect 527818 697592 527824 697604
rect 527232 697564 527824 697592
rect 527232 697552 527238 697564
rect 527818 697552 527824 697564
rect 527876 697592 527882 697604
rect 580166 697592 580172 697604
rect 527876 697564 580172 697592
rect 527876 697552 527882 697564
rect 580166 697552 580172 697564
rect 580224 697552 580230 697604
rect 3418 671168 3424 671220
rect 3476 671208 3482 671220
rect 8938 671208 8944 671220
rect 3476 671180 8944 671208
rect 3476 671168 3482 671180
rect 8938 671168 8944 671180
rect 8996 671168 9002 671220
rect 92934 586440 92940 586492
rect 92992 586480 92998 586492
rect 96154 586480 96160 586492
rect 92992 586452 96160 586480
rect 92992 586440 92998 586452
rect 96154 586440 96160 586452
rect 96212 586440 96218 586492
rect 373258 586440 373264 586492
rect 373316 586480 373322 586492
rect 376478 586480 376484 586492
rect 373316 586452 376484 586480
rect 373316 586440 373322 586452
rect 376478 586440 376484 586452
rect 376536 586440 376542 586492
rect 21818 586168 21824 586220
rect 21876 586208 21882 586220
rect 34514 586208 34520 586220
rect 21876 586180 34520 586208
rect 21876 586168 21882 586180
rect 34514 586168 34520 586180
rect 34572 586168 34578 586220
rect 193122 586168 193128 586220
rect 193180 586208 193186 586220
rect 200206 586208 200212 586220
rect 193180 586180 200212 586208
rect 193180 586168 193186 586180
rect 200206 586168 200212 586180
rect 200264 586168 200270 586220
rect 301774 586168 301780 586220
rect 301832 586208 301838 586220
rect 310790 586208 310796 586220
rect 301832 586180 310796 586208
rect 301832 586168 301838 586180
rect 310790 586168 310796 586180
rect 310848 586168 310854 586220
rect 21634 586100 21640 586152
rect 21692 586140 21698 586152
rect 42058 586140 42064 586152
rect 21692 586112 42064 586140
rect 21692 586100 21698 586112
rect 42058 586100 42064 586112
rect 42116 586100 42122 586152
rect 185670 586100 185676 586152
rect 185728 586140 185734 586152
rect 200298 586140 200304 586152
rect 185728 586112 200304 586140
rect 185728 586100 185734 586112
rect 200298 586100 200304 586112
rect 200356 586100 200362 586152
rect 301866 586100 301872 586152
rect 301924 586140 301930 586152
rect 314654 586140 314660 586152
rect 301924 586112 314660 586140
rect 301924 586100 301930 586112
rect 314654 586100 314660 586112
rect 314712 586100 314718 586152
rect 372614 586100 372620 586152
rect 372672 586140 372678 586152
rect 373258 586140 373264 586152
rect 372672 586112 373264 586140
rect 372672 586100 372678 586112
rect 373258 586100 373264 586112
rect 373316 586100 373322 586152
rect 465350 586100 465356 586152
rect 465408 586140 465414 586152
rect 479058 586140 479064 586152
rect 465408 586112 479064 586140
rect 465408 586100 465414 586112
rect 479058 586100 479064 586112
rect 479116 586100 479122 586152
rect 22922 586032 22928 586084
rect 22980 586072 22986 586084
rect 45922 586072 45928 586084
rect 22980 586044 45928 586072
rect 22980 586032 22986 586044
rect 45922 586032 45928 586044
rect 45980 586032 45986 586084
rect 181806 586032 181812 586084
rect 181864 586072 181870 586084
rect 198090 586072 198096 586084
rect 181864 586044 198096 586072
rect 181864 586032 181870 586044
rect 198090 586032 198096 586044
rect 198148 586032 198154 586084
rect 302694 586032 302700 586084
rect 302752 586072 302758 586084
rect 318518 586072 318524 586084
rect 302752 586044 318524 586072
rect 302752 586032 302758 586044
rect 318518 586032 318524 586044
rect 318576 586032 318582 586084
rect 461486 586032 461492 586084
rect 461544 586072 461550 586084
rect 478138 586072 478144 586084
rect 461544 586044 478144 586072
rect 461544 586032 461550 586044
rect 478138 586032 478144 586044
rect 478196 586032 478202 586084
rect 20530 585964 20536 586016
rect 20588 586004 20594 586016
rect 49786 586004 49792 586016
rect 20588 585976 49792 586004
rect 20588 585964 20594 585976
rect 49786 585964 49792 585976
rect 49844 585964 49850 586016
rect 177942 585964 177948 586016
rect 178000 586004 178006 586016
rect 198918 586004 198924 586016
rect 178000 585976 198924 586004
rect 178000 585964 178006 585976
rect 198918 585964 198924 585976
rect 198976 585964 198982 586016
rect 302142 585964 302148 586016
rect 302200 586004 302206 586016
rect 322382 586004 322388 586016
rect 302200 585976 322388 586004
rect 302200 585964 302206 585976
rect 322382 585964 322388 585976
rect 322440 585964 322446 586016
rect 457622 585964 457628 586016
rect 457680 586004 457686 586016
rect 478966 586004 478972 586016
rect 457680 585976 478972 586004
rect 457680 585964 457686 585976
rect 478966 585964 478972 585976
rect 479024 585964 479030 586016
rect 21726 585896 21732 585948
rect 21784 585936 21790 585948
rect 53834 585936 53840 585948
rect 21784 585908 53840 585936
rect 21784 585896 21790 585908
rect 53834 585896 53840 585908
rect 53892 585896 53898 585948
rect 173802 585896 173808 585948
rect 173860 585936 173866 585948
rect 197998 585936 198004 585948
rect 173860 585908 198004 585936
rect 173860 585896 173866 585908
rect 197998 585896 198004 585908
rect 198056 585896 198062 585948
rect 302878 585896 302884 585948
rect 302936 585936 302942 585948
rect 326246 585936 326252 585948
rect 302936 585908 326252 585936
rect 302936 585896 302942 585908
rect 326246 585896 326252 585908
rect 326304 585896 326310 585948
rect 453758 585896 453764 585948
rect 453816 585936 453822 585948
rect 477954 585936 477960 585948
rect 453816 585908 477960 585936
rect 453816 585896 453822 585908
rect 477954 585896 477960 585908
rect 478012 585896 478018 585948
rect 21910 585828 21916 585880
rect 21968 585868 21974 585880
rect 30466 585868 30472 585880
rect 21968 585840 30472 585868
rect 21968 585828 21974 585840
rect 30466 585828 30472 585840
rect 30524 585828 30530 585880
rect 32398 585828 32404 585880
rect 32456 585868 32462 585880
rect 65242 585868 65248 585880
rect 32456 585840 65248 585868
rect 32456 585828 32462 585840
rect 65242 585828 65248 585840
rect 65300 585828 65306 585880
rect 170214 585828 170220 585880
rect 170272 585868 170278 585880
rect 198734 585868 198740 585880
rect 170272 585840 198740 585868
rect 170272 585828 170278 585840
rect 198734 585828 198740 585840
rect 198792 585828 198798 585880
rect 301958 585828 301964 585880
rect 302016 585868 302022 585880
rect 330110 585868 330116 585880
rect 302016 585840 330116 585868
rect 302016 585828 302022 585840
rect 330110 585828 330116 585840
rect 330168 585828 330174 585880
rect 449894 585828 449900 585880
rect 449952 585868 449958 585880
rect 479150 585868 479156 585880
rect 449952 585840 479156 585868
rect 449952 585828 449958 585840
rect 479150 585828 479156 585840
rect 479208 585828 479214 585880
rect 22830 585760 22836 585812
rect 22888 585800 22894 585812
rect 38194 585800 38200 585812
rect 22888 585772 38200 585800
rect 22888 585760 22894 585772
rect 38194 585760 38200 585772
rect 38252 585760 38258 585812
rect 39298 585760 39304 585812
rect 39356 585800 39362 585812
rect 88426 585800 88432 585812
rect 39356 585772 88432 585800
rect 39356 585760 39362 585772
rect 88426 585760 88432 585772
rect 88484 585760 88490 585812
rect 166350 585760 166356 585812
rect 166408 585800 166414 585812
rect 197906 585800 197912 585812
rect 166408 585772 197912 585800
rect 166408 585760 166414 585772
rect 197906 585760 197912 585772
rect 197964 585760 197970 585812
rect 302786 585760 302792 585812
rect 302844 585800 302850 585812
rect 333974 585800 333980 585812
rect 302844 585772 333980 585800
rect 302844 585760 302850 585772
rect 333974 585760 333980 585772
rect 334032 585760 334038 585812
rect 446030 585760 446036 585812
rect 446088 585800 446094 585812
rect 477862 585800 477868 585812
rect 446088 585772 477868 585800
rect 446088 585760 446094 585772
rect 477862 585760 477868 585772
rect 477920 585760 477926 585812
rect 473078 585148 473084 585200
rect 473136 585188 473142 585200
rect 478046 585188 478052 585200
rect 473136 585160 478052 585188
rect 473136 585148 473142 585160
rect 478046 585148 478052 585160
rect 478104 585148 478110 585200
rect 300670 583380 300676 583432
rect 300728 583420 300734 583432
rect 341702 583420 341708 583432
rect 300728 583392 341708 583420
rect 300728 583380 300734 583392
rect 341702 583380 341708 583392
rect 341760 583380 341766 583432
rect 442166 583380 442172 583432
rect 442224 583420 442230 583432
rect 481634 583420 481640 583432
rect 442224 583392 481640 583420
rect 442224 583380 442230 583392
rect 481634 583380 481640 583392
rect 481692 583380 481698 583432
rect 158622 583312 158628 583364
rect 158680 583352 158686 583364
rect 201586 583352 201592 583364
rect 158680 583324 201592 583352
rect 158680 583312 158686 583324
rect 201586 583312 201592 583324
rect 201644 583312 201650 583364
rect 299290 583312 299296 583364
rect 299348 583352 299354 583364
rect 353294 583352 353300 583364
rect 299348 583324 353300 583352
rect 299348 583312 299354 583324
rect 353294 583312 353300 583324
rect 353352 583312 353358 583364
rect 426710 583312 426716 583364
rect 426768 583352 426774 583364
rect 481818 583352 481824 583364
rect 426768 583324 481824 583352
rect 426768 583312 426774 583324
rect 481818 583312 481824 583324
rect 481876 583312 481882 583364
rect 150894 583244 150900 583296
rect 150952 583284 150958 583296
rect 198826 583284 198832 583296
rect 150952 583256 198832 583284
rect 150952 583244 150958 583256
rect 198826 583244 198832 583256
rect 198884 583244 198890 583296
rect 300762 583244 300768 583296
rect 300820 583284 300826 583296
rect 357158 583284 357164 583296
rect 300820 583256 357164 583284
rect 300820 583244 300826 583256
rect 357158 583244 357164 583256
rect 357216 583244 357222 583296
rect 422846 583244 422852 583296
rect 422904 583284 422910 583296
rect 480714 583284 480720 583296
rect 422904 583256 480720 583284
rect 422904 583244 422910 583256
rect 480714 583244 480720 583256
rect 480772 583244 480778 583296
rect 147030 583176 147036 583228
rect 147088 583216 147094 583228
rect 201494 583216 201500 583228
rect 147088 583188 201500 583216
rect 147088 583176 147094 583188
rect 201494 583176 201500 583188
rect 201552 583176 201558 583228
rect 300578 583176 300584 583228
rect 300636 583216 300642 583228
rect 361022 583216 361028 583228
rect 300636 583188 361028 583216
rect 300636 583176 300642 583188
rect 361022 583176 361028 583188
rect 361080 583176 361086 583228
rect 415118 583176 415124 583228
rect 415176 583216 415182 583228
rect 478874 583216 478880 583228
rect 415176 583188 478880 583216
rect 415176 583176 415182 583188
rect 478874 583176 478880 583188
rect 478932 583176 478938 583228
rect 143166 583108 143172 583160
rect 143224 583148 143230 583160
rect 200390 583148 200396 583160
rect 143224 583120 200396 583148
rect 143224 583108 143230 583120
rect 200390 583108 200396 583120
rect 200448 583108 200454 583160
rect 300486 583108 300492 583160
rect 300544 583148 300550 583160
rect 364886 583148 364892 583160
rect 300544 583120 364892 583148
rect 300544 583108 300550 583120
rect 364886 583108 364892 583120
rect 364944 583108 364950 583160
rect 411254 583108 411260 583160
rect 411312 583148 411318 583160
rect 484394 583148 484400 583160
rect 411312 583120 484400 583148
rect 411312 583108 411318 583120
rect 484394 583108 484400 583120
rect 484452 583108 484458 583160
rect 127710 583040 127716 583092
rect 127768 583080 127774 583092
rect 200114 583080 200120 583092
rect 127768 583052 200120 583080
rect 127768 583040 127774 583052
rect 200114 583040 200120 583052
rect 200172 583040 200178 583092
rect 297818 583040 297824 583092
rect 297876 583080 297882 583092
rect 368750 583080 368756 583092
rect 297876 583052 368756 583080
rect 297876 583040 297882 583052
rect 368750 583040 368756 583052
rect 368808 583040 368814 583092
rect 407390 583040 407396 583092
rect 407448 583080 407454 583092
rect 483014 583080 483020 583092
rect 407448 583052 483020 583080
rect 407448 583040 407454 583052
rect 483014 583040 483020 583052
rect 483072 583040 483078 583092
rect 20622 582972 20628 583024
rect 20680 583012 20686 583024
rect 73154 583012 73160 583024
rect 20680 582984 73160 583012
rect 20680 582972 20686 582984
rect 73154 582972 73160 582984
rect 73212 582972 73218 583024
rect 123846 582972 123852 583024
rect 123904 583012 123910 583024
rect 199378 583012 199384 583024
rect 123904 582984 199384 583012
rect 123904 582972 123910 582984
rect 199378 582972 199384 582984
rect 199436 582972 199442 583024
rect 298002 582972 298008 583024
rect 298060 583012 298066 583024
rect 380342 583012 380348 583024
rect 298060 582984 380348 583012
rect 298060 582972 298066 582984
rect 380342 582972 380348 582984
rect 380400 582972 380406 583024
rect 403526 582972 403532 583024
rect 403584 583012 403590 583024
rect 480254 583012 480260 583024
rect 403584 582984 480260 583012
rect 403584 582972 403590 582984
rect 480254 582972 480260 582984
rect 480312 582972 480318 583024
rect 297910 580320 297916 580372
rect 297968 580360 297974 580372
rect 384206 580360 384212 580372
rect 297968 580332 384212 580360
rect 297968 580320 297974 580332
rect 384206 580320 384212 580332
rect 384264 580320 384270 580372
rect 399662 580320 399668 580372
rect 399720 580360 399726 580372
rect 483106 580360 483112 580372
rect 399720 580332 483112 580360
rect 399720 580320 399726 580332
rect 483106 580320 483112 580332
rect 483164 580320 483170 580372
rect 299382 580252 299388 580304
rect 299440 580292 299446 580304
rect 388070 580292 388076 580304
rect 299440 580264 388076 580292
rect 299440 580252 299446 580264
rect 388070 580252 388076 580264
rect 388128 580252 388134 580304
rect 395798 580252 395804 580304
rect 395856 580292 395862 580304
rect 483198 580292 483204 580304
rect 395856 580264 483204 580292
rect 395856 580252 395862 580264
rect 483198 580252 483204 580264
rect 483256 580252 483262 580304
rect 577498 577260 577504 577312
rect 577556 577300 577562 577312
rect 579614 577300 579620 577312
rect 577556 577272 579620 577300
rect 577556 577260 577562 577272
rect 579614 577260 579620 577272
rect 579672 577260 579678 577312
rect 19150 572364 19156 572416
rect 19208 572404 19214 572416
rect 32398 572404 32404 572416
rect 19208 572376 32404 572404
rect 19208 572364 19214 572376
rect 32398 572364 32404 572376
rect 32456 572364 32462 572416
rect 161474 572364 161480 572416
rect 161532 572404 161538 572416
rect 201770 572404 201776 572416
rect 161532 572376 201776 572404
rect 161532 572364 161538 572376
rect 201770 572364 201776 572376
rect 201828 572364 201834 572416
rect 18874 572296 18880 572348
rect 18932 572336 18938 572348
rect 39298 572336 39304 572348
rect 18932 572308 39304 572336
rect 18932 572296 18938 572308
rect 39298 572296 39304 572308
rect 39356 572296 39362 572348
rect 153194 572296 153200 572348
rect 153252 572336 153258 572348
rect 201678 572336 201684 572348
rect 153252 572308 201684 572336
rect 153252 572296 153258 572308
rect 201678 572296 201684 572308
rect 201736 572296 201742 572348
rect 19058 572228 19064 572280
rect 19116 572268 19122 572280
rect 75914 572268 75920 572280
rect 19116 572240 75920 572268
rect 19116 572228 19122 572240
rect 75914 572228 75920 572240
rect 75972 572228 75978 572280
rect 131114 572228 131120 572280
rect 131172 572268 131178 572280
rect 202966 572268 202972 572280
rect 131172 572240 202972 572268
rect 131172 572228 131178 572240
rect 202966 572228 202972 572240
rect 203024 572228 203030 572280
rect 20346 572160 20352 572212
rect 20404 572200 20410 572212
rect 80054 572200 80060 572212
rect 20404 572172 80060 572200
rect 20404 572160 20410 572172
rect 80054 572160 80060 572172
rect 80112 572160 80118 572212
rect 118694 572160 118700 572212
rect 118752 572200 118758 572212
rect 202874 572200 202880 572212
rect 118752 572172 202880 572200
rect 118752 572160 118758 572172
rect 202874 572160 202880 572172
rect 202932 572160 202938 572212
rect 19978 572092 19984 572144
rect 20036 572132 20042 572144
rect 99374 572132 99380 572144
rect 20036 572104 99380 572132
rect 20036 572092 20042 572104
rect 99374 572092 99380 572104
rect 99432 572092 99438 572144
rect 114554 572092 114560 572144
rect 114612 572132 114618 572144
rect 203058 572132 203064 572144
rect 114612 572104 203064 572132
rect 114612 572092 114618 572104
rect 203058 572092 203064 572104
rect 203116 572092 203122 572144
rect 18966 572024 18972 572076
rect 19024 572064 19030 572076
rect 103514 572064 103520 572076
rect 19024 572036 103520 572064
rect 19024 572024 19030 572036
rect 103514 572024 103520 572036
rect 103572 572024 103578 572076
rect 189074 572024 189080 572076
rect 189132 572064 189138 572076
rect 298738 572064 298744 572076
rect 189132 572036 298744 572064
rect 189132 572024 189138 572036
rect 298738 572024 298744 572036
rect 298796 572024 298802 572076
rect 300394 572024 300400 572076
rect 300452 572064 300458 572076
rect 345014 572064 345020 572076
rect 300452 572036 345020 572064
rect 300452 572024 300458 572036
rect 345014 572024 345020 572036
rect 345072 572024 345078 572076
rect 437474 572024 437480 572076
rect 437532 572064 437538 572076
rect 480530 572064 480536 572076
rect 437532 572036 480536 572064
rect 437532 572024 437538 572036
rect 480530 572024 480536 572036
rect 480588 572024 480594 572076
rect 20438 571956 20444 572008
rect 20496 571996 20502 572008
rect 107654 571996 107660 572008
rect 20496 571968 107660 571996
rect 20496 571956 20502 571968
rect 107654 571956 107660 571968
rect 107712 571956 107718 572008
rect 138014 571956 138020 572008
rect 138072 571996 138078 572008
rect 245654 571996 245660 572008
rect 138072 571968 245660 571996
rect 138072 571956 138078 571968
rect 245654 571956 245660 571968
rect 245712 571956 245718 572008
rect 247034 571956 247040 572008
rect 247092 571996 247098 572008
rect 418154 571996 418160 572008
rect 247092 571968 418160 571996
rect 247092 571956 247098 571968
rect 418154 571956 418160 571968
rect 418212 571956 418218 572008
rect 433334 571956 433340 572008
rect 433392 571996 433398 572008
rect 481726 571996 481732 572008
rect 433392 571968 481732 571996
rect 433392 571956 433398 571968
rect 481726 571956 481732 571968
rect 481784 571956 481790 572008
rect 263594 570596 263600 570648
rect 263652 570636 263658 570648
rect 373258 570636 373264 570648
rect 263652 570608 373264 570636
rect 263652 570596 263658 570608
rect 373258 570596 373264 570608
rect 373316 570596 373322 570648
rect 2774 565904 2780 565956
rect 2832 565944 2838 565956
rect 4890 565944 4896 565956
rect 2832 565916 4896 565944
rect 2832 565904 2838 565916
rect 4890 565904 4896 565916
rect 4948 565904 4954 565956
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 7558 514808 7564 514820
rect 3476 514780 7564 514808
rect 3476 514768 3482 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 480898 470568 480904 470620
rect 480956 470608 480962 470620
rect 580166 470608 580172 470620
rect 480956 470580 580172 470608
rect 480956 470568 480962 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 20254 465740 20260 465792
rect 20312 465780 20318 465792
rect 20530 465780 20536 465792
rect 20312 465752 20536 465780
rect 20312 465740 20318 465752
rect 20530 465740 20536 465752
rect 20588 465740 20594 465792
rect 478782 462884 478788 462936
rect 478840 462924 478846 462936
rect 480438 462924 480444 462936
rect 478840 462896 480444 462924
rect 478840 462884 478846 462896
rect 480438 462884 480444 462896
rect 480496 462884 480502 462936
rect 22094 462612 22100 462664
rect 22152 462652 22158 462664
rect 23198 462652 23204 462664
rect 22152 462624 23204 462652
rect 22152 462612 22158 462624
rect 23198 462612 23204 462624
rect 23256 462612 23262 462664
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 199010 462340 199016 462392
rect 199068 462380 199074 462392
rect 199378 462380 199384 462392
rect 199068 462352 199384 462380
rect 199068 462340 199074 462352
rect 199378 462340 199384 462352
rect 199436 462380 199442 462392
rect 204254 462380 204260 462392
rect 199436 462352 204260 462380
rect 199436 462340 199442 462352
rect 204254 462340 204260 462352
rect 204312 462340 204318 462392
rect 392210 462340 392216 462392
rect 392268 462380 392274 462392
rect 478782 462380 478788 462392
rect 392268 462352 478788 462380
rect 392268 462340 392274 462352
rect 478782 462340 478788 462352
rect 478840 462340 478846 462392
rect 300302 462272 300308 462324
rect 300360 462312 300366 462324
rect 300486 462312 300492 462324
rect 300360 462284 300492 462312
rect 300360 462272 300366 462284
rect 300486 462272 300492 462284
rect 300544 462272 300550 462324
rect 479150 462272 479156 462324
rect 479208 462312 479214 462324
rect 479334 462312 479340 462324
rect 479208 462284 479340 462312
rect 479208 462272 479214 462284
rect 479334 462272 479340 462284
rect 479392 462272 479398 462324
rect 480622 462272 480628 462324
rect 480680 462312 480686 462324
rect 481634 462312 481640 462324
rect 480680 462284 481640 462312
rect 480680 462272 480686 462284
rect 481634 462272 481640 462284
rect 481692 462272 481698 462324
rect 20162 461524 20168 461576
rect 20220 461564 20226 461576
rect 20438 461564 20444 461576
rect 20220 461536 20444 461564
rect 20220 461524 20226 461536
rect 20438 461524 20444 461536
rect 20496 461524 20502 461576
rect 18598 461320 18604 461372
rect 18656 461360 18662 461372
rect 18966 461360 18972 461372
rect 18656 461332 18972 461360
rect 18656 461320 18662 461332
rect 18966 461320 18972 461332
rect 19024 461320 19030 461372
rect 18874 461116 18880 461168
rect 18932 461156 18938 461168
rect 88426 461156 88432 461168
rect 18932 461128 88432 461156
rect 18932 461116 18938 461128
rect 88426 461116 88432 461128
rect 88484 461116 88490 461168
rect 158622 461116 158628 461168
rect 158680 461156 158686 461168
rect 201586 461156 201592 461168
rect 158680 461128 201592 461156
rect 158680 461116 158686 461128
rect 201586 461116 201592 461128
rect 201644 461116 201650 461168
rect 300302 461116 300308 461168
rect 300360 461156 300366 461168
rect 364242 461156 364248 461168
rect 300360 461128 364248 461156
rect 300360 461116 300366 461128
rect 364242 461116 364248 461128
rect 364300 461116 364306 461168
rect 453942 461116 453948 461168
rect 454000 461156 454006 461168
rect 477954 461156 477960 461168
rect 454000 461128 477960 461156
rect 454000 461116 454006 461128
rect 477954 461116 477960 461128
rect 478012 461116 478018 461168
rect 17770 461048 17776 461100
rect 17828 461088 17834 461100
rect 19978 461088 19984 461100
rect 17828 461060 19984 461088
rect 17828 461048 17834 461060
rect 19978 461048 19984 461060
rect 20036 461088 20042 461100
rect 100340 461088 100346 461100
rect 20036 461060 100346 461088
rect 20036 461048 20042 461060
rect 100340 461048 100346 461060
rect 100398 461048 100404 461100
rect 146708 461048 146714 461100
rect 146766 461088 146772 461100
rect 201494 461088 201500 461100
rect 146766 461060 201500 461088
rect 146766 461048 146772 461060
rect 201494 461048 201500 461060
rect 201552 461048 201558 461100
rect 300762 461048 300768 461100
rect 300820 461088 300826 461100
rect 357158 461088 357164 461100
rect 300820 461060 357164 461088
rect 300820 461048 300826 461060
rect 357158 461048 357164 461060
rect 357216 461048 357222 461100
rect 449894 461048 449900 461100
rect 449952 461088 449958 461100
rect 479334 461088 479340 461100
rect 449952 461060 479340 461088
rect 449952 461048 449958 461060
rect 479334 461048 479340 461060
rect 479392 461048 479398 461100
rect 18966 460980 18972 461032
rect 19024 461020 19030 461032
rect 104204 461020 104210 461032
rect 19024 460992 104210 461020
rect 19024 460980 19030 460992
rect 104204 460980 104210 460992
rect 104262 460980 104268 461032
rect 142844 460980 142850 461032
rect 142902 461020 142908 461032
rect 200390 461020 200396 461032
rect 142902 460992 200396 461020
rect 142902 460980 142908 460992
rect 200390 460980 200396 460992
rect 200448 460980 200454 461032
rect 300578 460980 300584 461032
rect 300636 461020 300642 461032
rect 361022 461020 361028 461032
rect 300636 460992 361028 461020
rect 300636 460980 300642 460992
rect 361022 460980 361028 460992
rect 361080 460980 361086 461032
rect 446030 460980 446036 461032
rect 446088 461020 446094 461032
rect 477862 461020 477868 461032
rect 446088 460992 477868 461020
rect 446088 460980 446094 460992
rect 477862 460980 477868 460992
rect 477920 460980 477926 461032
rect 480622 461020 480628 461032
rect 480226 460992 480628 461020
rect 20162 460912 20168 460964
rect 20220 460952 20226 460964
rect 107746 460952 107752 460964
rect 20220 460924 107752 460952
rect 20220 460912 20226 460924
rect 107746 460912 107752 460924
rect 107804 460912 107810 460964
rect 123846 460912 123852 460964
rect 123904 460952 123910 460964
rect 199010 460952 199016 460964
rect 123904 460924 199016 460952
rect 123904 460912 123910 460924
rect 199010 460912 199016 460924
rect 199068 460912 199074 460964
rect 297910 460912 297916 460964
rect 297968 460952 297974 460964
rect 384206 460952 384212 460964
rect 297968 460924 384212 460952
rect 297968 460912 297974 460924
rect 384206 460912 384212 460924
rect 384264 460912 384270 460964
rect 442166 460912 442172 460964
rect 442224 460952 442230 460964
rect 480226 460952 480254 460992
rect 480622 460980 480628 460992
rect 480680 460980 480686 461032
rect 442224 460924 480254 460952
rect 442224 460912 442230 460924
rect 177942 460844 177948 460896
rect 178000 460884 178006 460896
rect 198918 460884 198924 460896
rect 178000 460856 198924 460884
rect 178000 460844 178006 460856
rect 198918 460844 198924 460856
rect 198976 460844 198982 460896
rect 473078 460844 473084 460896
rect 473136 460884 473142 460896
rect 478046 460884 478052 460896
rect 473136 460856 478052 460884
rect 473136 460844 473142 460856
rect 478046 460844 478052 460856
rect 478104 460844 478110 460896
rect 22002 459484 22008 459536
rect 22060 459524 22066 459536
rect 26602 459524 26608 459536
rect 22060 459496 26608 459524
rect 22060 459484 22066 459496
rect 26602 459484 26608 459496
rect 26660 459484 26666 459536
rect 92934 459484 92940 459536
rect 92992 459524 92998 459536
rect 95878 459524 95884 459536
rect 92992 459496 95884 459524
rect 92992 459484 92998 459496
rect 95878 459484 95884 459496
rect 95936 459484 95942 459536
rect 115842 459484 115848 459536
rect 115900 459524 115906 459536
rect 203242 459524 203248 459536
rect 115900 459496 203248 459524
rect 115900 459484 115906 459496
rect 203242 459484 203248 459496
rect 203300 459484 203306 459536
rect 372614 459484 372620 459536
rect 372672 459524 372678 459536
rect 373258 459524 373264 459536
rect 372672 459496 373264 459524
rect 372672 459484 372678 459496
rect 373258 459484 373264 459496
rect 373316 459524 373322 459536
rect 376478 459524 376484 459536
rect 373316 459496 376484 459524
rect 373316 459484 373322 459496
rect 376478 459484 376484 459496
rect 376536 459484 376542 459536
rect 415118 459484 415124 459536
rect 415176 459524 415182 459536
rect 418706 459524 418712 459536
rect 415176 459496 418712 459524
rect 415176 459484 415182 459496
rect 418706 459484 418712 459496
rect 418764 459484 418770 459536
rect 457622 459484 457628 459536
rect 457680 459524 457686 459536
rect 461486 459524 461492 459536
rect 457680 459496 461492 459524
rect 457680 459484 457686 459496
rect 461486 459484 461492 459496
rect 461544 459484 461550 459536
rect 461578 459484 461584 459536
rect 461636 459524 461642 459536
rect 463786 459524 463792 459536
rect 461636 459496 463792 459524
rect 461636 459484 461642 459496
rect 463786 459484 463792 459496
rect 463844 459484 463850 459536
rect 465350 459484 465356 459536
rect 465408 459524 465414 459536
rect 469306 459524 469312 459536
rect 465408 459496 469312 459524
rect 465408 459484 465414 459496
rect 469306 459484 469312 459496
rect 469364 459484 469370 459536
rect 18966 459416 18972 459468
rect 19024 459456 19030 459468
rect 76834 459456 76840 459468
rect 19024 459428 76840 459456
rect 19024 459416 19030 459428
rect 76834 459416 76840 459428
rect 76892 459416 76898 459468
rect 131574 459416 131580 459468
rect 131632 459456 131638 459468
rect 202966 459456 202972 459468
rect 131632 459428 202972 459456
rect 131632 459416 131638 459428
rect 202966 459416 202972 459428
rect 203024 459416 203030 459468
rect 298002 459416 298008 459468
rect 298060 459456 298066 459468
rect 380342 459456 380348 459468
rect 298060 459428 380348 459456
rect 298060 459416 298066 459428
rect 380342 459416 380348 459428
rect 380400 459416 380406 459468
rect 407390 459416 407396 459468
rect 407448 459456 407454 459468
rect 483014 459456 483020 459468
rect 407448 459428 483020 459456
rect 407448 459416 407454 459428
rect 483014 459416 483020 459428
rect 483072 459416 483078 459468
rect 19242 459348 19248 459400
rect 19300 459388 19306 459400
rect 61378 459388 61384 459400
rect 19300 459360 61384 459388
rect 19300 459348 19306 459360
rect 61378 459348 61384 459360
rect 61436 459348 61442 459400
rect 135162 459348 135168 459400
rect 135220 459388 135226 459400
rect 197354 459388 197360 459400
rect 135220 459360 197360 459388
rect 135220 459348 135226 459360
rect 197354 459348 197360 459360
rect 197412 459348 197418 459400
rect 297818 459348 297824 459400
rect 297876 459388 297882 459400
rect 368750 459388 368756 459400
rect 297876 459360 368756 459388
rect 297876 459348 297882 459360
rect 368750 459348 368756 459360
rect 368808 459348 368814 459400
rect 411254 459348 411260 459400
rect 411312 459388 411318 459400
rect 484394 459388 484400 459400
rect 411312 459360 484400 459388
rect 411312 459348 411318 459360
rect 484394 459348 484400 459360
rect 484452 459348 484458 459400
rect 20346 459280 20352 459332
rect 20404 459320 20410 459332
rect 80698 459320 80704 459332
rect 20404 459292 80704 459320
rect 20404 459280 20410 459292
rect 80698 459280 80704 459292
rect 80756 459280 80762 459332
rect 162486 459280 162492 459332
rect 162544 459320 162550 459332
rect 201862 459320 201868 459332
rect 162544 459292 201868 459320
rect 162544 459280 162550 459292
rect 201862 459280 201868 459292
rect 201920 459280 201926 459332
rect 299290 459280 299296 459332
rect 299348 459320 299354 459332
rect 353294 459320 353300 459332
rect 299348 459292 353300 459320
rect 299348 459280 299354 459292
rect 353294 459280 353300 459292
rect 353352 459280 353358 459332
rect 430574 459280 430580 459332
rect 430632 459320 430638 459332
rect 479150 459320 479156 459332
rect 430632 459292 479156 459320
rect 430632 459280 430638 459292
rect 479150 459280 479156 459292
rect 479208 459280 479214 459332
rect 300486 459212 300492 459264
rect 300544 459252 300550 459264
rect 345566 459252 345572 459264
rect 300544 459224 345572 459252
rect 300544 459212 300550 459224
rect 345566 459212 345572 459224
rect 345624 459212 345630 459264
rect 438302 459212 438308 459264
rect 438360 459252 438366 459264
rect 480530 459252 480536 459264
rect 438360 459224 480536 459252
rect 438360 459212 438366 459224
rect 480530 459212 480536 459224
rect 480588 459212 480594 459264
rect 300670 459144 300676 459196
rect 300728 459184 300734 459196
rect 341702 459184 341708 459196
rect 300728 459156 341708 459184
rect 300728 459144 300734 459156
rect 341702 459144 341708 459156
rect 341760 459144 341766 459196
rect 403526 459144 403532 459196
rect 403584 459184 403590 459196
rect 480254 459184 480260 459196
rect 403584 459156 480260 459184
rect 403584 459144 403590 459156
rect 480254 459144 480260 459156
rect 480312 459184 480318 459196
rect 482094 459184 482100 459196
rect 480312 459156 482100 459184
rect 480312 459144 480318 459156
rect 482094 459144 482100 459156
rect 482152 459144 482158 459196
rect 299382 459076 299388 459128
rect 299440 459116 299446 459128
rect 388070 459116 388076 459128
rect 299440 459088 388076 459116
rect 299440 459076 299446 459088
rect 388070 459076 388076 459088
rect 388128 459076 388134 459128
rect 19150 459008 19156 459060
rect 19208 459048 19214 459060
rect 20438 459048 20444 459060
rect 19208 459020 20444 459048
rect 19208 459008 19214 459020
rect 20438 459008 20444 459020
rect 20496 459008 20502 459060
rect 42794 459008 42800 459060
rect 42852 459048 42858 459060
rect 45922 459048 45928 459060
rect 42852 459020 45928 459048
rect 42852 459008 42858 459020
rect 45922 459008 45928 459020
rect 45980 459008 45986 459060
rect 20622 458940 20628 458992
rect 20680 458980 20686 458992
rect 21450 458980 21456 458992
rect 20680 458952 21456 458980
rect 20680 458940 20686 458952
rect 21450 458940 21456 458952
rect 21508 458940 21514 458992
rect 22738 458940 22744 458992
rect 22796 458980 22802 458992
rect 30466 458980 30472 458992
rect 22796 458952 30472 458980
rect 22796 458940 22802 458952
rect 30466 458940 30472 458952
rect 30524 458940 30530 458992
rect 154482 458940 154488 458992
rect 154540 458980 154546 458992
rect 200390 458980 200396 458992
rect 154540 458952 200396 458980
rect 154540 458940 154546 458952
rect 200390 458940 200396 458952
rect 200448 458980 200454 458992
rect 201678 458980 201684 458992
rect 200448 458952 201684 458980
rect 200448 458940 200454 458952
rect 201678 458940 201684 458952
rect 201736 458940 201742 458992
rect 20438 458872 20444 458924
rect 20496 458912 20502 458924
rect 65242 458912 65248 458924
rect 20496 458884 65248 458912
rect 20496 458872 20502 458884
rect 65242 458872 65248 458884
rect 65300 458872 65306 458924
rect 119982 458872 119988 458924
rect 120040 458912 120046 458924
rect 197170 458912 197176 458924
rect 120040 458884 197176 458912
rect 120040 458872 120046 458884
rect 197170 458872 197176 458884
rect 197228 458912 197234 458924
rect 202874 458912 202880 458924
rect 197228 458884 202880 458912
rect 197228 458872 197234 458884
rect 202874 458872 202880 458884
rect 202932 458872 202938 458924
rect 469214 458872 469220 458924
rect 469272 458912 469278 458924
rect 481634 458912 481640 458924
rect 469272 458884 481640 458912
rect 469272 458872 469278 458884
rect 481634 458872 481640 458884
rect 481692 458872 481698 458924
rect 21450 458804 21456 458856
rect 21508 458844 21514 458856
rect 73154 458844 73160 458856
rect 21508 458816 73160 458844
rect 21508 458804 21514 458816
rect 73154 458804 73160 458816
rect 73212 458804 73218 458856
rect 139302 458804 139308 458856
rect 139360 458844 139366 458856
rect 244274 458844 244280 458856
rect 139360 458816 244280 458844
rect 139360 458804 139366 458816
rect 244274 458804 244280 458816
rect 244332 458804 244338 458856
rect 283558 458804 283564 458856
rect 283616 458844 283622 458856
rect 418982 458844 418988 458856
rect 283616 458816 418988 458844
rect 283616 458804 283622 458816
rect 418982 458804 418988 458816
rect 419040 458804 419046 458856
rect 434438 458804 434444 458856
rect 434496 458844 434502 458856
rect 480346 458844 480352 458856
rect 434496 458816 480352 458844
rect 434496 458804 434502 458816
rect 480346 458804 480352 458816
rect 480404 458844 480410 458856
rect 481726 458844 481732 458856
rect 480404 458816 481732 458844
rect 480404 458804 480410 458816
rect 481726 458804 481732 458816
rect 481784 458804 481790 458856
rect 30374 458464 30380 458516
rect 30432 458504 30438 458516
rect 34514 458504 34520 458516
rect 30432 458476 34520 458504
rect 30432 458464 30438 458476
rect 34514 458464 34520 458476
rect 34572 458464 34578 458516
rect 18782 458192 18788 458244
rect 18840 458232 18846 458244
rect 19242 458232 19248 458244
rect 18840 458204 19248 458232
rect 18840 458192 18846 458204
rect 19242 458192 19248 458204
rect 19300 458192 19306 458244
rect 483014 458192 483020 458244
rect 483072 458232 483078 458244
rect 484486 458232 484492 458244
rect 483072 458204 484492 458232
rect 483072 458192 483078 458204
rect 484486 458192 484492 458204
rect 484544 458192 484550 458244
rect 150894 458124 150900 458176
rect 150952 458164 150958 458176
rect 198826 458164 198832 458176
rect 150952 458136 198832 458164
rect 150952 458124 150958 458136
rect 198826 458124 198832 458136
rect 198884 458124 198890 458176
rect 302786 458124 302792 458176
rect 302844 458164 302850 458176
rect 333974 458164 333980 458176
rect 302844 458136 333980 458164
rect 302844 458124 302850 458136
rect 333974 458124 333980 458136
rect 334032 458124 334038 458176
rect 395798 458124 395804 458176
rect 395856 458164 395862 458176
rect 483290 458164 483296 458176
rect 395856 458136 483296 458164
rect 395856 458124 395862 458136
rect 483290 458124 483296 458136
rect 483348 458124 483354 458176
rect 20254 458056 20260 458108
rect 20312 458096 20318 458108
rect 49786 458096 49792 458108
rect 20312 458068 49792 458096
rect 20312 458056 20318 458068
rect 49786 458056 49792 458068
rect 49844 458056 49850 458108
rect 166350 458056 166356 458108
rect 166408 458096 166414 458108
rect 197906 458096 197912 458108
rect 166408 458068 197912 458096
rect 166408 458056 166414 458068
rect 197906 458056 197912 458068
rect 197964 458056 197970 458108
rect 301958 458056 301964 458108
rect 302016 458096 302022 458108
rect 330110 458096 330116 458108
rect 302016 458068 330116 458096
rect 302016 458056 302022 458068
rect 330110 458056 330116 458068
rect 330168 458056 330174 458108
rect 399662 458056 399668 458108
rect 399720 458096 399726 458108
rect 483106 458096 483112 458108
rect 399720 458068 483112 458096
rect 399720 458056 399726 458068
rect 483106 458056 483112 458068
rect 483164 458056 483170 458108
rect 21910 457988 21916 458040
rect 21968 458028 21974 458040
rect 22738 458028 22744 458040
rect 21968 458000 22744 458028
rect 21968 457988 21974 458000
rect 22738 457988 22744 458000
rect 22796 457988 22802 458040
rect 22922 457988 22928 458040
rect 22980 458028 22986 458040
rect 42794 458028 42800 458040
rect 22980 458000 42800 458028
rect 22980 457988 22986 458000
rect 42794 457988 42800 458000
rect 42852 457988 42858 458040
rect 170214 457988 170220 458040
rect 170272 458028 170278 458040
rect 198734 458028 198740 458040
rect 170272 458000 198740 458028
rect 170272 457988 170278 458000
rect 198734 457988 198740 458000
rect 198792 457988 198798 458040
rect 302878 457988 302884 458040
rect 302936 458028 302942 458040
rect 326246 458028 326252 458040
rect 302936 458000 326252 458028
rect 302936 457988 302942 458000
rect 326246 457988 326252 458000
rect 326304 457988 326310 458040
rect 418706 457988 418712 458040
rect 418764 458028 418770 458040
rect 478874 458028 478880 458040
rect 418764 458000 478880 458028
rect 418764 457988 418770 458000
rect 478874 457988 478880 458000
rect 478932 457988 478938 458040
rect 21726 457920 21732 457972
rect 21784 457960 21790 457972
rect 53834 457960 53840 457972
rect 21784 457932 53840 457960
rect 21784 457920 21790 457932
rect 53834 457920 53840 457932
rect 53892 457920 53898 457972
rect 422846 457920 422852 457972
rect 422904 457960 422910 457972
rect 480714 457960 480720 457972
rect 422904 457932 480720 457960
rect 422904 457920 422910 457932
rect 480714 457920 480720 457932
rect 480772 457960 480778 457972
rect 483198 457960 483204 457972
rect 480772 457932 483204 457960
rect 480772 457920 480778 457932
rect 483198 457920 483204 457932
rect 483256 457920 483262 457972
rect 426710 457852 426716 457904
rect 426768 457892 426774 457904
rect 481818 457892 481824 457904
rect 426768 457864 481824 457892
rect 426768 457852 426774 457864
rect 481818 457852 481824 457864
rect 481876 457852 481882 457904
rect 21818 457444 21824 457496
rect 21876 457484 21882 457496
rect 22830 457484 22836 457496
rect 21876 457456 22836 457484
rect 21876 457444 21882 457456
rect 22830 457444 22836 457456
rect 22888 457484 22894 457496
rect 30374 457484 30380 457496
rect 22888 457456 30380 457484
rect 22888 457444 22894 457456
rect 30374 457444 30380 457456
rect 30432 457444 30438 457496
rect 20530 456764 20536 456816
rect 20588 456804 20594 456816
rect 22922 456804 22928 456816
rect 20588 456776 22928 456804
rect 20588 456764 20594 456776
rect 22922 456764 22928 456776
rect 22980 456764 22986 456816
rect 197906 456764 197912 456816
rect 197964 456804 197970 456816
rect 198090 456804 198096 456816
rect 197964 456776 198096 456804
rect 197964 456764 197970 456776
rect 198090 456764 198096 456776
rect 198148 456764 198154 456816
rect 198826 456764 198832 456816
rect 198884 456804 198890 456816
rect 199010 456804 199016 456816
rect 198884 456776 199016 456804
rect 198884 456764 198890 456776
rect 199010 456764 199016 456776
rect 199068 456764 199074 456816
rect 302602 456764 302608 456816
rect 302660 456804 302666 456816
rect 302786 456804 302792 456816
rect 302660 456776 302792 456804
rect 302660 456764 302666 456776
rect 302786 456764 302792 456776
rect 302844 456764 302850 456816
rect 478782 456696 478788 456748
rect 478840 456736 478846 456748
rect 480438 456736 480444 456748
rect 478840 456708 480444 456736
rect 478840 456696 478846 456708
rect 480438 456696 480444 456708
rect 480496 456696 480502 456748
rect 264974 445000 264980 445052
rect 265032 445040 265038 445052
rect 373258 445040 373264 445052
rect 265032 445012 373264 445040
rect 265032 445000 265038 445012
rect 373258 445000 373264 445012
rect 373316 445000 373322 445052
rect 126974 444320 126980 444372
rect 127032 444360 127038 444372
rect 200114 444360 200120 444372
rect 127032 444332 200120 444360
rect 127032 444320 127038 444332
rect 200114 444320 200120 444332
rect 200172 444360 200178 444372
rect 201770 444360 201776 444372
rect 200172 444332 201776 444360
rect 200172 444320 200178 444332
rect 201770 444320 201776 444332
rect 201828 444320 201834 444372
rect 21542 443912 21548 443964
rect 21600 443952 21606 443964
rect 23474 443952 23480 443964
rect 21600 443924 23480 443952
rect 21600 443912 21606 443924
rect 23474 443912 23480 443924
rect 23532 443912 23538 443964
rect 197262 443708 197268 443760
rect 197320 443748 197326 443760
rect 204346 443748 204352 443760
rect 197320 443720 204352 443748
rect 197320 443708 197326 443720
rect 204346 443708 204352 443720
rect 204404 443708 204410 443760
rect 95878 443640 95884 443692
rect 95936 443680 95942 443692
rect 260834 443680 260840 443692
rect 95936 443652 260840 443680
rect 95936 443640 95942 443652
rect 260834 443640 260840 443652
rect 260892 443640 260898 443692
rect 2866 410184 2872 410236
rect 2924 410224 2930 410236
rect 4982 410224 4988 410236
rect 2924 410196 4988 410224
rect 2924 410184 2930 410196
rect 4982 410184 4988 410196
rect 5040 410184 5046 410236
rect 479518 364352 479524 364404
rect 479576 364392 479582 364404
rect 580166 364392 580172 364404
rect 479576 364364 580172 364392
rect 479576 364352 479582 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 20898 345080 20904 345092
rect 3384 345052 20904 345080
rect 3384 345040 3390 345052
rect 20898 345040 20904 345052
rect 20956 345040 20962 345092
rect 200482 335248 200488 335300
rect 200540 335288 200546 335300
rect 200540 335260 200620 335288
rect 200540 335248 200546 335260
rect 200592 335096 200620 335260
rect 200574 335044 200580 335096
rect 200632 335044 200638 335096
rect 21450 334636 21456 334688
rect 21508 334676 21514 334688
rect 72970 334676 72976 334688
rect 21508 334648 72976 334676
rect 21508 334636 21514 334648
rect 72970 334636 72976 334648
rect 73028 334636 73034 334688
rect 18598 334568 18604 334620
rect 18656 334608 18662 334620
rect 103882 334608 103888 334620
rect 18656 334580 103888 334608
rect 18656 334568 18662 334580
rect 103882 334568 103888 334580
rect 103940 334568 103946 334620
rect 17954 334092 17960 334144
rect 18012 334132 18018 334144
rect 18598 334132 18604 334144
rect 18012 334104 18604 334132
rect 18012 334092 18018 334104
rect 18598 334092 18604 334104
rect 18656 334092 18662 334144
rect 19242 334024 19248 334076
rect 19300 334064 19306 334076
rect 19300 334036 26234 334064
rect 19300 334024 19306 334036
rect 19150 333956 19156 334008
rect 19208 333996 19214 334008
rect 21450 333996 21456 334008
rect 19208 333968 21456 333996
rect 19208 333956 19214 333968
rect 21450 333956 21456 333968
rect 21508 333956 21514 334008
rect 26206 333996 26234 334036
rect 76834 333996 76840 334008
rect 26206 333968 76840 333996
rect 76834 333956 76840 333968
rect 76892 333956 76898 334008
rect 442442 333956 442448 334008
rect 442500 333996 442506 334008
rect 480622 333996 480628 334008
rect 442500 333968 480628 333996
rect 442500 333956 442506 333968
rect 480622 333956 480628 333968
rect 480680 333956 480686 334008
rect 478414 333276 478420 333328
rect 478472 333316 478478 333328
rect 479150 333316 479156 333328
rect 478472 333288 479156 333316
rect 478472 333276 478478 333288
rect 479150 333276 479156 333288
rect 479208 333276 479214 333328
rect 438854 333208 438860 333260
rect 438912 333248 438918 333260
rect 480530 333248 480536 333260
rect 438912 333220 480536 333248
rect 438912 333208 438918 333220
rect 480530 333208 480536 333220
rect 480588 333248 480594 333260
rect 482002 333248 482008 333260
rect 480588 333220 482008 333248
rect 480588 333208 480594 333220
rect 482002 333208 482008 333220
rect 482060 333208 482066 333260
rect 162486 332936 162492 332988
rect 162544 332976 162550 332988
rect 201678 332976 201684 332988
rect 162544 332948 201684 332976
rect 162544 332936 162550 332948
rect 201678 332936 201684 332948
rect 201736 332976 201742 332988
rect 201862 332976 201868 332988
rect 201736 332948 201868 332976
rect 201736 332936 201742 332948
rect 201862 332936 201868 332948
rect 201920 332936 201926 332988
rect 158714 332868 158720 332920
rect 158772 332908 158778 332920
rect 201586 332908 201592 332920
rect 158772 332880 201592 332908
rect 158772 332868 158778 332880
rect 201586 332868 201592 332880
rect 201644 332908 201650 332920
rect 201954 332908 201960 332920
rect 201644 332880 201960 332908
rect 201644 332868 201650 332880
rect 201954 332868 201960 332880
rect 202012 332868 202018 332920
rect 299290 332868 299296 332920
rect 299348 332908 299354 332920
rect 300118 332908 300124 332920
rect 299348 332880 300124 332908
rect 299348 332868 299354 332880
rect 300118 332868 300124 332880
rect 300176 332908 300182 332920
rect 350534 332908 350540 332920
rect 300176 332880 350540 332908
rect 300176 332868 300182 332880
rect 350534 332868 350540 332880
rect 350592 332868 350598 332920
rect 8938 332800 8944 332852
rect 8996 332840 9002 332852
rect 26602 332840 26608 332852
rect 8996 332812 26608 332840
rect 8996 332800 9002 332812
rect 26602 332800 26608 332812
rect 26660 332800 26666 332852
rect 154758 332800 154764 332852
rect 154816 332840 154822 332852
rect 200298 332840 200304 332852
rect 154816 332812 200304 332840
rect 154816 332800 154822 332812
rect 200298 332800 200304 332812
rect 200356 332800 200362 332852
rect 302878 332800 302884 332852
rect 302936 332840 302942 332852
rect 361574 332840 361580 332852
rect 302936 332812 361580 332840
rect 302936 332800 302942 332812
rect 361574 332800 361580 332812
rect 361632 332800 361638 332852
rect 20346 332732 20352 332784
rect 20404 332772 20410 332784
rect 80698 332772 80704 332784
rect 20404 332744 80704 332772
rect 20404 332732 20410 332744
rect 80698 332732 80704 332744
rect 80756 332732 80762 332784
rect 137922 332732 137928 332784
rect 137980 332772 137986 332784
rect 197354 332772 197360 332784
rect 137980 332744 197360 332772
rect 137980 332732 137986 332744
rect 197354 332732 197360 332744
rect 197412 332732 197418 332784
rect 297726 332732 297732 332784
rect 297784 332772 297790 332784
rect 368750 332772 368756 332784
rect 297784 332744 368756 332772
rect 297784 332732 297790 332744
rect 368750 332732 368756 332744
rect 368808 332732 368814 332784
rect 433242 332732 433248 332784
rect 433300 332772 433306 332784
rect 478414 332772 478420 332784
rect 433300 332744 478420 332772
rect 433300 332732 433306 332744
rect 478414 332732 478420 332744
rect 478472 332732 478478 332784
rect 16482 332664 16488 332716
rect 16540 332704 16546 332716
rect 17770 332704 17776 332716
rect 16540 332676 17776 332704
rect 16540 332664 16546 332676
rect 17770 332664 17776 332676
rect 17828 332704 17834 332716
rect 100018 332704 100024 332716
rect 17828 332676 100024 332704
rect 17828 332664 17834 332676
rect 100018 332664 100024 332676
rect 100076 332664 100082 332716
rect 143166 332664 143172 332716
rect 143224 332704 143230 332716
rect 200390 332704 200396 332716
rect 143224 332676 200396 332704
rect 143224 332664 143230 332676
rect 200390 332664 200396 332676
rect 200448 332704 200454 332716
rect 202046 332704 202052 332716
rect 200448 332676 202052 332704
rect 200448 332664 200454 332676
rect 202046 332664 202052 332676
rect 202104 332664 202110 332716
rect 297910 332664 297916 332716
rect 297968 332704 297974 332716
rect 384206 332704 384212 332716
rect 297968 332676 384212 332704
rect 297968 332664 297974 332676
rect 384206 332664 384212 332676
rect 384264 332664 384270 332716
rect 395798 332664 395804 332716
rect 395856 332704 395862 332716
rect 483198 332704 483204 332716
rect 395856 332676 483204 332704
rect 395856 332664 395862 332676
rect 483198 332664 483204 332676
rect 483256 332664 483262 332716
rect 20070 332596 20076 332648
rect 20128 332636 20134 332648
rect 107746 332636 107752 332648
rect 20128 332608 107752 332636
rect 20128 332596 20134 332608
rect 107746 332596 107752 332608
rect 107804 332596 107810 332648
rect 123846 332596 123852 332648
rect 123904 332636 123910 332648
rect 199930 332636 199936 332648
rect 123904 332608 199936 332636
rect 123904 332596 123910 332608
rect 199930 332596 199936 332608
rect 199988 332636 199994 332648
rect 199988 332608 200114 332636
rect 199988 332596 199994 332608
rect 3602 332528 3608 332580
rect 3660 332568 3666 332580
rect 22922 332568 22928 332580
rect 3660 332540 22928 332568
rect 3660 332528 3666 332540
rect 22922 332528 22928 332540
rect 22980 332528 22986 332580
rect 92934 332528 92940 332580
rect 92992 332568 92998 332580
rect 96430 332568 96436 332580
rect 92992 332540 96436 332568
rect 92992 332528 92998 332540
rect 96430 332528 96436 332540
rect 96488 332528 96494 332580
rect 135070 332528 135076 332580
rect 135128 332568 135134 332580
rect 137922 332568 137928 332580
rect 135128 332540 137928 332568
rect 135128 332528 135134 332540
rect 137922 332528 137928 332540
rect 137980 332528 137986 332580
rect 166350 332528 166356 332580
rect 166408 332568 166414 332580
rect 198090 332568 198096 332580
rect 166408 332540 198096 332568
rect 166408 332528 166414 332540
rect 198090 332528 198096 332540
rect 198148 332528 198154 332580
rect 200086 332568 200114 332608
rect 306926 332596 306932 332648
rect 306984 332636 306990 332648
rect 577498 332636 577504 332648
rect 306984 332608 577504 332636
rect 306984 332596 306990 332608
rect 577498 332596 577504 332608
rect 577556 332596 577562 332648
rect 204254 332568 204260 332580
rect 200086 332540 204260 332568
rect 204254 332528 204260 332540
rect 204312 332528 204318 332580
rect 300486 332528 300492 332580
rect 300544 332568 300550 332580
rect 345566 332568 345572 332580
rect 300544 332540 345572 332568
rect 300544 332528 300550 332540
rect 345566 332528 345572 332540
rect 345624 332528 345630 332580
rect 350534 332528 350540 332580
rect 350592 332568 350598 332580
rect 353294 332568 353300 332580
rect 350592 332540 353300 332568
rect 350592 332528 350598 332540
rect 353294 332528 353300 332540
rect 353352 332528 353358 332580
rect 361574 332528 361580 332580
rect 361632 332568 361638 332580
rect 364886 332568 364892 332580
rect 361632 332540 364892 332568
rect 361632 332528 361638 332540
rect 364886 332528 364892 332540
rect 364944 332528 364950 332580
rect 372614 332528 372620 332580
rect 372672 332568 372678 332580
rect 376478 332568 376484 332580
rect 372672 332540 376484 332568
rect 372672 332528 372678 332540
rect 376478 332528 376484 332540
rect 376536 332528 376542 332580
rect 430574 332528 430580 332580
rect 430632 332568 430638 332580
rect 433242 332568 433248 332580
rect 430632 332540 433248 332568
rect 430632 332528 430638 332540
rect 433242 332528 433248 332540
rect 433300 332528 433306 332580
rect 473078 332528 473084 332580
rect 473136 332568 473142 332580
rect 478046 332568 478052 332580
rect 473136 332540 478052 332568
rect 473136 332528 473142 332540
rect 478046 332528 478052 332540
rect 478104 332568 478110 332580
rect 478104 332540 480254 332568
rect 478104 332528 478110 332540
rect 20162 332460 20168 332512
rect 20220 332500 20226 332512
rect 49786 332500 49792 332512
rect 20220 332472 49792 332500
rect 20220 332460 20226 332472
rect 49786 332460 49792 332472
rect 49844 332460 49850 332512
rect 170214 332460 170220 332512
rect 170272 332500 170278 332512
rect 198826 332500 198832 332512
rect 170272 332472 198832 332500
rect 170272 332460 170278 332472
rect 198826 332460 198832 332472
rect 198884 332460 198890 332512
rect 301958 332460 301964 332512
rect 302016 332500 302022 332512
rect 330110 332500 330116 332512
rect 302016 332472 330116 332500
rect 302016 332460 302022 332472
rect 330110 332460 330116 332472
rect 330168 332460 330174 332512
rect 449894 332460 449900 332512
rect 449952 332500 449958 332512
rect 479334 332500 479340 332512
rect 449952 332472 479340 332500
rect 449952 332460 449958 332472
rect 479334 332460 479340 332472
rect 479392 332460 479398 332512
rect 20530 332392 20536 332444
rect 20588 332432 20594 332444
rect 45922 332432 45928 332444
rect 20588 332404 45928 332432
rect 20588 332392 20594 332404
rect 45922 332392 45928 332404
rect 45980 332392 45986 332444
rect 173710 332392 173716 332444
rect 173768 332432 173774 332444
rect 197998 332432 198004 332444
rect 173768 332404 198004 332432
rect 173768 332392 173774 332404
rect 197998 332392 198004 332404
rect 198056 332392 198062 332444
rect 302786 332392 302792 332444
rect 302844 332432 302850 332444
rect 326246 332432 326252 332444
rect 302844 332404 326252 332432
rect 302844 332392 302850 332404
rect 326246 332392 326252 332404
rect 326304 332392 326310 332444
rect 453758 332392 453764 332444
rect 453816 332432 453822 332444
rect 477954 332432 477960 332444
rect 453816 332404 477960 332432
rect 453816 332392 453822 332404
rect 477954 332392 477960 332404
rect 478012 332392 478018 332444
rect 480226 332432 480254 332540
rect 481910 332432 481916 332444
rect 480226 332404 481916 332432
rect 481910 332392 481916 332404
rect 481968 332392 481974 332444
rect 22554 332324 22560 332376
rect 22612 332364 22618 332376
rect 38194 332364 38200 332376
rect 22612 332336 38200 332364
rect 22612 332324 22618 332336
rect 38194 332324 38200 332336
rect 38252 332324 38258 332376
rect 177942 332324 177948 332376
rect 178000 332364 178006 332376
rect 198918 332364 198924 332376
rect 178000 332336 198924 332364
rect 178000 332324 178006 332336
rect 198918 332324 198924 332336
rect 198976 332324 198982 332376
rect 301866 332324 301872 332376
rect 301924 332364 301930 332376
rect 322382 332364 322388 332376
rect 301924 332336 322388 332364
rect 301924 332324 301930 332336
rect 322382 332324 322388 332336
rect 322440 332324 322446 332376
rect 457622 332324 457628 332376
rect 457680 332364 457686 332376
rect 478966 332364 478972 332376
rect 457680 332336 478972 332364
rect 457680 332324 457686 332336
rect 478966 332324 478972 332336
rect 479024 332324 479030 332376
rect 22830 332256 22836 332308
rect 22888 332296 22894 332308
rect 34514 332296 34520 332308
rect 22888 332268 34520 332296
rect 22888 332256 22894 332268
rect 34514 332256 34520 332268
rect 34572 332256 34578 332308
rect 181806 332256 181812 332308
rect 181864 332296 181870 332308
rect 198182 332296 198188 332308
rect 181864 332268 198188 332296
rect 181864 332256 181870 332268
rect 198182 332256 198188 332268
rect 198240 332256 198246 332308
rect 302694 332256 302700 332308
rect 302752 332296 302758 332308
rect 318518 332296 318524 332308
rect 302752 332268 318524 332296
rect 302752 332256 302758 332268
rect 318518 332256 318524 332268
rect 318576 332256 318582 332308
rect 461486 332256 461492 332308
rect 461544 332296 461550 332308
rect 478138 332296 478144 332308
rect 461544 332268 478144 332296
rect 461544 332256 461550 332268
rect 478138 332256 478144 332268
rect 478196 332256 478202 332308
rect 22646 332188 22652 332240
rect 22704 332228 22710 332240
rect 30466 332228 30472 332240
rect 22704 332200 30472 332228
rect 22704 332188 22710 332200
rect 30466 332188 30472 332200
rect 30524 332188 30530 332240
rect 185670 332188 185676 332240
rect 185728 332228 185734 332240
rect 200206 332228 200212 332240
rect 185728 332200 200212 332228
rect 185728 332188 185734 332200
rect 200206 332188 200212 332200
rect 200264 332228 200270 332240
rect 200666 332228 200672 332240
rect 200264 332200 200672 332228
rect 200264 332188 200270 332200
rect 200666 332188 200672 332200
rect 200724 332188 200730 332240
rect 301498 332188 301504 332240
rect 301556 332228 301562 332240
rect 314654 332228 314660 332240
rect 301556 332200 314660 332228
rect 301556 332188 301562 332200
rect 314654 332188 314660 332200
rect 314712 332188 314718 332240
rect 465350 332188 465356 332240
rect 465408 332228 465414 332240
rect 479058 332228 479064 332240
rect 465408 332200 479064 332228
rect 465408 332188 465414 332200
rect 479058 332188 479064 332200
rect 479116 332188 479122 332240
rect 21910 332120 21916 332172
rect 21968 332160 21974 332172
rect 53834 332160 53840 332172
rect 21968 332132 53840 332160
rect 21968 332120 21974 332132
rect 53834 332120 53840 332132
rect 53892 332120 53898 332172
rect 193030 332120 193036 332172
rect 193088 332160 193094 332172
rect 200574 332160 200580 332172
rect 193088 332132 200580 332160
rect 193088 332120 193094 332132
rect 200574 332120 200580 332132
rect 200632 332120 200638 332172
rect 302050 332120 302056 332172
rect 302108 332160 302114 332172
rect 310790 332160 310796 332172
rect 302108 332132 310796 332160
rect 302108 332120 302114 332132
rect 310790 332120 310796 332132
rect 310848 332120 310854 332172
rect 446030 332120 446036 332172
rect 446088 332160 446094 332172
rect 477862 332160 477868 332172
rect 446088 332132 477868 332160
rect 446088 332120 446094 332132
rect 477862 332120 477868 332132
rect 477920 332120 477926 332172
rect 22186 331848 22192 331900
rect 22244 331888 22250 331900
rect 42058 331888 42064 331900
rect 22244 331860 42064 331888
rect 22244 331848 22250 331860
rect 42058 331848 42064 331860
rect 42116 331848 42122 331900
rect 301682 331780 301688 331832
rect 301740 331820 301746 331832
rect 302050 331820 302056 331832
rect 301740 331792 302056 331820
rect 301740 331780 301746 331792
rect 302050 331780 302056 331792
rect 302108 331780 302114 331832
rect 22002 331440 22008 331492
rect 22060 331480 22066 331492
rect 22554 331480 22560 331492
rect 22060 331452 22560 331480
rect 22060 331440 22066 331452
rect 22554 331440 22560 331452
rect 22612 331440 22618 331492
rect 17770 331236 17776 331288
rect 17828 331276 17834 331288
rect 21542 331276 21548 331288
rect 17828 331248 21548 331276
rect 17828 331236 17834 331248
rect 21542 331236 21548 331248
rect 21600 331236 21606 331288
rect 22646 331236 22652 331288
rect 22704 331276 22710 331288
rect 22922 331276 22928 331288
rect 22704 331248 22928 331276
rect 22704 331236 22710 331248
rect 22922 331236 22928 331248
rect 22980 331236 22986 331288
rect 84562 331276 84568 331288
rect 84166 331248 84568 331276
rect 21560 331140 21588 331236
rect 84166 331140 84194 331248
rect 84562 331236 84568 331248
rect 84620 331236 84626 331288
rect 197906 331236 197912 331288
rect 197964 331276 197970 331288
rect 198090 331276 198096 331288
rect 197964 331248 198096 331276
rect 197964 331236 197970 331248
rect 198090 331236 198096 331248
rect 198148 331236 198154 331288
rect 301498 331236 301504 331288
rect 301556 331276 301562 331288
rect 301774 331276 301780 331288
rect 301556 331248 301780 331276
rect 301556 331236 301562 331248
rect 301774 331236 301780 331248
rect 301832 331236 301838 331288
rect 399662 331236 399668 331288
rect 399720 331276 399726 331288
rect 400858 331276 400864 331288
rect 399720 331248 400864 331276
rect 399720 331236 399726 331248
rect 400858 331236 400864 331248
rect 400916 331236 400922 331288
rect 403526 331236 403532 331288
rect 403584 331276 403590 331288
rect 404998 331276 405004 331288
rect 403584 331248 405004 331276
rect 403584 331236 403590 331248
rect 404998 331236 405004 331248
rect 405056 331236 405062 331288
rect 415118 331236 415124 331288
rect 415176 331276 415182 331288
rect 415176 331248 418108 331276
rect 415176 331236 415182 331248
rect 127710 331168 127716 331220
rect 127768 331208 127774 331220
rect 418080 331208 418108 331248
rect 477862 331236 477868 331288
rect 477920 331276 477926 331288
rect 478322 331276 478328 331288
rect 477920 331248 478328 331276
rect 477920 331236 477926 331248
rect 478322 331236 478328 331248
rect 478380 331236 478386 331288
rect 478874 331236 478880 331288
rect 478932 331276 478938 331288
rect 479058 331276 479064 331288
rect 478932 331248 479064 331276
rect 478932 331236 478938 331248
rect 479058 331236 479064 331248
rect 479116 331236 479122 331288
rect 418614 331208 418620 331220
rect 127768 331180 180794 331208
rect 418080 331180 418620 331208
rect 127768 331168 127774 331180
rect 21560 331112 84194 331140
rect 180766 331140 180794 331180
rect 418614 331168 418620 331180
rect 418672 331168 418678 331220
rect 201862 331140 201868 331152
rect 180766 331112 201868 331140
rect 201862 331100 201868 331112
rect 201920 331100 201926 331152
rect 18874 331032 18880 331084
rect 18932 331072 18938 331084
rect 88426 331072 88432 331084
rect 18932 331044 88432 331072
rect 18932 331032 18938 331044
rect 88426 331032 88432 331044
rect 88484 331032 88490 331084
rect 21634 330964 21640 331016
rect 21692 331004 21698 331016
rect 22186 331004 22192 331016
rect 21692 330976 22192 331004
rect 21692 330964 21698 330976
rect 22186 330964 22192 330976
rect 22244 330964 22250 331016
rect 147030 330556 147036 330608
rect 147088 330596 147094 330608
rect 200390 330596 200396 330608
rect 147088 330568 200396 330596
rect 147088 330556 147094 330568
rect 200390 330556 200396 330568
rect 200448 330596 200454 330608
rect 201494 330596 201500 330608
rect 200448 330568 201500 330596
rect 200448 330556 200454 330568
rect 201494 330556 201500 330568
rect 201552 330556 201558 330608
rect 119982 330488 119988 330540
rect 120040 330528 120046 330540
rect 203058 330528 203064 330540
rect 120040 330500 203064 330528
rect 120040 330488 120046 330500
rect 203058 330488 203064 330500
rect 203116 330528 203122 330540
rect 204346 330528 204352 330540
rect 203116 330500 204352 330528
rect 203116 330488 203122 330500
rect 204346 330488 204352 330500
rect 204404 330488 204410 330540
rect 18782 329740 18788 329792
rect 18840 329780 18846 329792
rect 18966 329780 18972 329792
rect 18840 329752 18972 329780
rect 18840 329740 18846 329752
rect 18966 329740 18972 329752
rect 19024 329740 19030 329792
rect 20254 329740 20260 329792
rect 20312 329780 20318 329792
rect 20438 329780 20444 329792
rect 20312 329752 20444 329780
rect 20312 329740 20318 329752
rect 20438 329740 20444 329752
rect 20496 329780 20502 329792
rect 65242 329780 65248 329792
rect 20496 329752 65248 329780
rect 20496 329740 20502 329752
rect 65242 329740 65248 329752
rect 65300 329740 65306 329792
rect 131022 329740 131028 329792
rect 131080 329780 131086 329792
rect 202966 329780 202972 329792
rect 131080 329752 202972 329780
rect 131080 329740 131086 329752
rect 202966 329740 202972 329752
rect 203024 329780 203030 329792
rect 203150 329780 203156 329792
rect 203024 329752 203156 329780
rect 203024 329740 203030 329752
rect 203150 329740 203156 329752
rect 203208 329740 203214 329792
rect 407390 329740 407396 329792
rect 407448 329780 407454 329792
rect 484486 329780 484492 329792
rect 407448 329752 484492 329780
rect 407448 329740 407454 329752
rect 484486 329740 484492 329752
rect 484544 329740 484550 329792
rect 18984 329712 19012 329740
rect 61378 329712 61384 329724
rect 18984 329684 61384 329712
rect 61378 329672 61384 329684
rect 61436 329672 61442 329724
rect 411254 329672 411260 329724
rect 411312 329712 411318 329724
rect 484394 329712 484400 329724
rect 411312 329684 484400 329712
rect 411312 329672 411318 329684
rect 484394 329672 484400 329684
rect 484452 329672 484458 329724
rect 418614 329604 418620 329656
rect 418672 329644 418678 329656
rect 477494 329644 477500 329656
rect 418672 329616 477500 329644
rect 418672 329604 418678 329616
rect 477494 329604 477500 329616
rect 477552 329604 477558 329656
rect 484394 329400 484400 329452
rect 484452 329440 484458 329452
rect 484578 329440 484584 329452
rect 484452 329412 484584 329440
rect 484452 329400 484458 329412
rect 484578 329400 484584 329412
rect 484636 329400 484642 329452
rect 3602 318792 3608 318844
rect 3660 318832 3666 318844
rect 21450 318832 21456 318844
rect 3660 318804 21456 318832
rect 3660 318792 3666 318804
rect 21450 318792 21456 318804
rect 21508 318792 21514 318844
rect 249794 318044 249800 318096
rect 249852 318084 249858 318096
rect 418154 318084 418160 318096
rect 249852 318056 418160 318084
rect 249852 318044 249858 318056
rect 418154 318044 418160 318056
rect 418212 318044 418218 318096
rect 138014 316684 138020 316736
rect 138072 316724 138078 316736
rect 241514 316724 241520 316736
rect 138072 316696 241520 316724
rect 138072 316684 138078 316696
rect 241514 316684 241520 316696
rect 241572 316684 241578 316736
rect 114554 315936 114560 315988
rect 114612 315976 114618 315988
rect 203242 315976 203248 315988
rect 114612 315948 203248 315976
rect 114612 315936 114618 315948
rect 203242 315936 203248 315948
rect 203300 315936 203306 315988
rect 298002 315936 298008 315988
rect 298060 315976 298066 315988
rect 379514 315976 379520 315988
rect 298060 315948 379520 315976
rect 298060 315936 298066 315948
rect 379514 315936 379520 315948
rect 379572 315936 379578 315988
rect 391934 315936 391940 315988
rect 391992 315976 391998 315988
rect 480438 315976 480444 315988
rect 391992 315948 480444 315976
rect 391992 315936 391998 315948
rect 480438 315936 480444 315948
rect 480496 315936 480502 315988
rect 150342 315868 150348 315920
rect 150400 315908 150406 315920
rect 199010 315908 199016 315920
rect 150400 315880 199016 315908
rect 150400 315868 150406 315880
rect 199010 315868 199016 315880
rect 199068 315868 199074 315920
rect 300578 315868 300584 315920
rect 300636 315908 300642 315920
rect 360194 315908 360200 315920
rect 300636 315880 360200 315908
rect 300636 315868 300642 315880
rect 360194 315868 360200 315880
rect 360252 315868 360258 315920
rect 404998 315868 405004 315920
rect 405056 315908 405062 315920
rect 482094 315908 482100 315920
rect 405056 315880 482100 315908
rect 405056 315868 405062 315880
rect 482094 315868 482100 315880
rect 482152 315868 482158 315920
rect 300762 315800 300768 315852
rect 300820 315840 300826 315852
rect 356054 315840 356060 315852
rect 300820 315812 356060 315840
rect 300820 315800 300826 315812
rect 356054 315800 356060 315812
rect 356112 315800 356118 315852
rect 400858 315800 400864 315852
rect 400916 315840 400922 315852
rect 476114 315840 476120 315852
rect 400916 315812 476120 315840
rect 400916 315800 400922 315812
rect 476114 315800 476120 315812
rect 476172 315800 476178 315852
rect 302142 315732 302148 315784
rect 302200 315772 302206 315784
rect 349154 315772 349160 315784
rect 302200 315744 349160 315772
rect 302200 315732 302206 315744
rect 349154 315732 349160 315744
rect 349212 315732 349218 315784
rect 422294 315732 422300 315784
rect 422352 315772 422358 315784
rect 483106 315772 483112 315784
rect 422352 315744 483112 315772
rect 422352 315732 422358 315744
rect 483106 315732 483112 315744
rect 483164 315732 483170 315784
rect 300670 315664 300676 315716
rect 300728 315704 300734 315716
rect 340874 315704 340880 315716
rect 300728 315676 340880 315704
rect 300728 315664 300734 315676
rect 340874 315664 340880 315676
rect 340932 315664 340938 315716
rect 426434 315664 426440 315716
rect 426492 315704 426498 315716
rect 481818 315704 481824 315716
rect 426492 315676 481824 315704
rect 426492 315664 426498 315676
rect 481818 315664 481824 315676
rect 481876 315664 481882 315716
rect 303522 315596 303528 315648
rect 303580 315636 303586 315648
rect 336734 315636 336740 315648
rect 303580 315608 336740 315636
rect 303580 315596 303586 315608
rect 336734 315596 336740 315608
rect 336792 315596 336798 315648
rect 433334 315596 433340 315648
rect 433392 315636 433398 315648
rect 480346 315636 480352 315648
rect 433392 315608 480352 315636
rect 433392 315596 433398 315608
rect 480346 315596 480352 315608
rect 480404 315596 480410 315648
rect 302602 315528 302608 315580
rect 302660 315568 302666 315580
rect 333974 315568 333980 315580
rect 302660 315540 333980 315568
rect 302660 315528 302666 315540
rect 333974 315528 333980 315540
rect 334032 315528 334038 315580
rect 111794 315324 111800 315376
rect 111852 315364 111858 315376
rect 200482 315364 200488 315376
rect 111852 315336 200488 315364
rect 111852 315324 111858 315336
rect 200482 315324 200488 315336
rect 200540 315324 200546 315376
rect 301590 315324 301596 315376
rect 301648 315364 301654 315376
rect 302142 315364 302148 315376
rect 301648 315336 302148 315364
rect 301648 315324 301654 315336
rect 302142 315324 302148 315336
rect 302200 315324 302206 315376
rect 195974 315256 195980 315308
rect 196032 315296 196038 315308
rect 298830 315296 298836 315308
rect 196032 315268 298836 315296
rect 196032 315256 196038 315268
rect 298830 315256 298836 315268
rect 298888 315256 298894 315308
rect 481726 315188 481732 315240
rect 481784 315228 481790 315240
rect 482094 315228 482100 315240
rect 481784 315200 482100 315228
rect 481784 315188 481790 315200
rect 482094 315188 482100 315200
rect 482152 315188 482158 315240
rect 302602 314780 302608 314832
rect 302660 314820 302666 314832
rect 302878 314820 302884 314832
rect 302660 314792 302884 314820
rect 302660 314780 302666 314792
rect 302878 314780 302884 314792
rect 302936 314780 302942 314832
rect 198734 314644 198740 314696
rect 198792 314684 198798 314696
rect 199010 314684 199016 314696
rect 198792 314656 199016 314684
rect 198792 314644 198798 314656
rect 199010 314644 199016 314656
rect 199068 314644 199074 314696
rect 202966 314644 202972 314696
rect 203024 314684 203030 314696
rect 203242 314684 203248 314696
rect 203024 314656 203248 314684
rect 203024 314644 203030 314656
rect 203242 314644 203248 314656
rect 203300 314644 203306 314696
rect 300578 314644 300584 314696
rect 300636 314684 300642 314696
rect 300762 314684 300768 314696
rect 300636 314656 300768 314684
rect 300636 314644 300642 314656
rect 300762 314644 300768 314656
rect 300820 314644 300826 314696
rect 481818 314644 481824 314696
rect 481876 314684 481882 314696
rect 483382 314684 483388 314696
rect 481876 314656 483388 314684
rect 481876 314644 481882 314656
rect 483382 314644 483388 314656
rect 483440 314644 483446 314696
rect 299382 314236 299388 314288
rect 299440 314276 299446 314288
rect 300210 314276 300216 314288
rect 299440 314248 300216 314276
rect 299440 314236 299446 314248
rect 300210 314236 300216 314248
rect 300268 314236 300274 314288
rect 2774 292612 2780 292664
rect 2832 292652 2838 292664
rect 5074 292652 5080 292664
rect 2832 292624 5080 292652
rect 2832 292612 2838 292624
rect 5074 292612 5080 292624
rect 5132 292612 5138 292664
rect 3326 240116 3332 240168
rect 3384 240156 3390 240168
rect 17218 240156 17224 240168
rect 3384 240128 17224 240156
rect 3384 240116 3390 240128
rect 17218 240116 17224 240128
rect 17276 240116 17282 240168
rect 481174 207000 481180 207052
rect 481232 207040 481238 207052
rect 483014 207040 483020 207052
rect 481232 207012 483020 207040
rect 481232 207000 481238 207012
rect 483014 207000 483020 207012
rect 483072 207000 483078 207052
rect 476114 206524 476120 206576
rect 476172 206564 476178 206576
rect 480438 206564 480444 206576
rect 476172 206536 480444 206564
rect 476172 206524 476178 206536
rect 480438 206524 480444 206536
rect 480496 206524 480502 206576
rect 297910 206320 297916 206372
rect 297968 206360 297974 206372
rect 313274 206360 313280 206372
rect 297968 206332 313280 206360
rect 297968 206320 297974 206332
rect 313274 206320 313280 206332
rect 313332 206320 313338 206372
rect 16390 206252 16396 206304
rect 16448 206292 16454 206304
rect 17862 206292 17868 206304
rect 16448 206264 17868 206292
rect 16448 206252 16454 206264
rect 17862 206252 17868 206264
rect 17920 206292 17926 206304
rect 103882 206292 103888 206304
rect 17920 206264 103888 206292
rect 17920 206252 17926 206264
rect 103882 206252 103888 206264
rect 103940 206252 103946 206304
rect 300210 206252 300216 206304
rect 300268 206292 300274 206304
rect 387794 206292 387800 206304
rect 300268 206264 387800 206292
rect 300268 206252 300274 206264
rect 387794 206252 387800 206264
rect 387852 206252 387858 206304
rect 162486 205844 162492 205896
rect 162544 205884 162550 205896
rect 201494 205884 201500 205896
rect 162544 205856 201500 205884
rect 162544 205844 162550 205856
rect 201494 205844 201500 205856
rect 201552 205844 201558 205896
rect 158622 205776 158628 205828
rect 158680 205816 158686 205828
rect 201770 205816 201776 205828
rect 158680 205788 201776 205816
rect 158680 205776 158686 205788
rect 201770 205776 201776 205788
rect 201828 205816 201834 205828
rect 201954 205816 201960 205828
rect 201828 205788 201960 205816
rect 201828 205776 201834 205788
rect 201954 205776 201960 205788
rect 202012 205776 202018 205828
rect 154574 205708 154580 205760
rect 154632 205748 154638 205760
rect 200114 205748 200120 205760
rect 154632 205720 200120 205748
rect 154632 205708 154638 205720
rect 200114 205708 200120 205720
rect 200172 205748 200178 205760
rect 200298 205748 200304 205760
rect 200172 205720 200304 205748
rect 200172 205708 200178 205720
rect 200298 205708 200304 205720
rect 200356 205708 200362 205760
rect 438578 205708 438584 205760
rect 438636 205748 438642 205760
rect 480714 205748 480720 205760
rect 438636 205720 480720 205748
rect 438636 205708 438642 205720
rect 480714 205708 480720 205720
rect 480772 205748 480778 205760
rect 482002 205748 482008 205760
rect 480772 205720 482008 205748
rect 480772 205708 480778 205720
rect 482002 205708 482008 205720
rect 482060 205708 482066 205760
rect 20346 205640 20352 205692
rect 20404 205680 20410 205692
rect 28902 205680 28908 205692
rect 20404 205652 28908 205680
rect 20404 205640 20410 205652
rect 28902 205640 28908 205652
rect 28960 205640 28966 205692
rect 143166 205640 143172 205692
rect 143224 205680 143230 205692
rect 201586 205680 201592 205692
rect 143224 205652 201592 205680
rect 143224 205640 143230 205652
rect 201586 205640 201592 205652
rect 201644 205680 201650 205692
rect 202046 205680 202052 205692
rect 201644 205652 202052 205680
rect 201644 205640 201650 205652
rect 202046 205640 202052 205652
rect 202104 205640 202110 205692
rect 392210 205640 392216 205692
rect 392268 205680 392274 205692
rect 476114 205680 476120 205692
rect 392268 205652 476120 205680
rect 392268 205640 392274 205652
rect 476114 205640 476120 205652
rect 476172 205640 476178 205692
rect 299382 204892 299388 204944
rect 299440 204932 299446 204944
rect 300118 204932 300124 204944
rect 299440 204904 300124 204932
rect 299440 204892 299446 204904
rect 300118 204892 300124 204904
rect 300176 204932 300182 204944
rect 349246 204932 349252 204944
rect 300176 204904 349252 204932
rect 300176 204892 300182 204904
rect 349246 204892 349252 204904
rect 349304 204892 349310 204944
rect 434714 204688 434720 204740
rect 434772 204728 434778 204740
rect 480346 204728 480352 204740
rect 434772 204700 480352 204728
rect 434772 204688 434778 204700
rect 480346 204688 480352 204700
rect 480404 204688 480410 204740
rect 300670 204620 300676 204672
rect 300728 204660 300734 204672
rect 341334 204660 341340 204672
rect 300728 204632 341340 204660
rect 300728 204620 300734 204632
rect 341334 204620 341340 204632
rect 341392 204620 341398 204672
rect 418706 204620 418712 204672
rect 418764 204660 418770 204672
rect 479058 204660 479064 204672
rect 418764 204632 479064 204660
rect 418764 204620 418770 204632
rect 479058 204620 479064 204632
rect 479116 204620 479122 204672
rect 302878 204552 302884 204604
rect 302936 204592 302942 204604
rect 333974 204592 333980 204604
rect 302936 204564 333980 204592
rect 302936 204552 302942 204564
rect 333974 204552 333980 204564
rect 334032 204552 334038 204604
rect 407022 204552 407028 204604
rect 407080 204592 407086 204604
rect 481726 204592 481732 204604
rect 407080 204564 481732 204592
rect 407080 204552 407086 204564
rect 481726 204552 481732 204564
rect 481784 204552 481790 204604
rect 300578 204484 300584 204536
rect 300636 204524 300642 204536
rect 357158 204524 357164 204536
rect 300636 204496 357164 204524
rect 300636 204484 300642 204496
rect 357158 204484 357164 204496
rect 357216 204484 357222 204536
rect 426710 204484 426716 204536
rect 426768 204524 426774 204536
rect 483382 204524 483388 204536
rect 426768 204496 483388 204524
rect 426768 204484 426774 204496
rect 483382 204484 483388 204496
rect 483440 204484 483446 204536
rect 296622 204416 296628 204468
rect 296680 204456 296686 204468
rect 298002 204456 298008 204468
rect 296680 204428 298008 204456
rect 296680 204416 296686 204428
rect 298002 204416 298008 204428
rect 298060 204456 298066 204468
rect 380342 204456 380348 204468
rect 298060 204428 380348 204456
rect 298060 204416 298066 204428
rect 380342 204416 380348 204428
rect 380400 204416 380406 204468
rect 422846 204416 422852 204468
rect 422904 204456 422910 204468
rect 483106 204456 483112 204468
rect 422904 204428 483112 204456
rect 422904 204416 422910 204428
rect 483106 204416 483112 204428
rect 483164 204416 483170 204468
rect 306926 204348 306932 204400
rect 306984 204388 306990 204400
rect 480898 204388 480904 204400
rect 306984 204360 480904 204388
rect 306984 204348 306990 204360
rect 480898 204348 480904 204360
rect 480956 204348 480962 204400
rect 23014 204320 23020 204332
rect 22848 204292 23020 204320
rect 7558 204212 7564 204264
rect 7616 204252 7622 204264
rect 22848 204252 22876 204292
rect 23014 204280 23020 204292
rect 23072 204280 23078 204332
rect 147030 204280 147036 204332
rect 147088 204320 147094 204332
rect 197354 204320 197360 204332
rect 147088 204292 197360 204320
rect 147088 204280 147094 204292
rect 197354 204280 197360 204292
rect 197412 204280 197418 204332
rect 202874 204320 202880 204332
rect 200086 204292 202880 204320
rect 7616 204224 22876 204252
rect 7616 204212 7622 204224
rect 22922 204212 22928 204264
rect 22980 204252 22986 204264
rect 30466 204252 30472 204264
rect 22980 204224 30472 204252
rect 22980 204212 22986 204224
rect 30466 204212 30472 204224
rect 30524 204212 30530 204264
rect 92934 204212 92940 204264
rect 92992 204252 92998 204264
rect 95878 204252 95884 204264
rect 92992 204224 95884 204252
rect 92992 204212 92998 204224
rect 95878 204212 95884 204224
rect 95936 204252 95942 204264
rect 96154 204252 96160 204264
rect 95936 204224 96160 204252
rect 95936 204212 95942 204224
rect 96154 204212 96160 204224
rect 96212 204212 96218 204264
rect 177942 204212 177948 204264
rect 178000 204252 178006 204264
rect 179874 204252 179880 204264
rect 178000 204224 179880 204252
rect 178000 204212 178006 204224
rect 179874 204212 179880 204224
rect 179932 204212 179938 204264
rect 199930 204252 199936 204264
rect 180766 204224 199936 204252
rect 19058 204144 19064 204196
rect 19116 204184 19122 204196
rect 19242 204184 19248 204196
rect 19116 204156 19248 204184
rect 19116 204144 19122 204156
rect 19242 204144 19248 204156
rect 19300 204184 19306 204196
rect 76834 204184 76840 204196
rect 19300 204156 76840 204184
rect 19300 204144 19306 204156
rect 76834 204144 76840 204156
rect 76892 204144 76898 204196
rect 123846 204144 123852 204196
rect 123904 204184 123910 204196
rect 180766 204184 180794 204224
rect 199930 204212 199936 204224
rect 199988 204252 199994 204264
rect 200086 204252 200114 204292
rect 202874 204280 202880 204292
rect 202932 204280 202938 204332
rect 303062 204280 303068 204332
rect 303120 204320 303126 204332
rect 580534 204320 580540 204332
rect 303120 204292 580540 204320
rect 303120 204280 303126 204292
rect 580534 204280 580540 204292
rect 580592 204280 580598 204332
rect 199988 204224 200114 204252
rect 199988 204212 199994 204224
rect 302694 204212 302700 204264
rect 302752 204252 302758 204264
rect 318518 204252 318524 204264
rect 302752 204224 318524 204252
rect 302752 204212 302758 204224
rect 318518 204212 318524 204224
rect 318576 204212 318582 204264
rect 349246 204212 349252 204264
rect 349304 204252 349310 204264
rect 353294 204252 353300 204264
rect 349304 204224 353300 204252
rect 349304 204212 349310 204224
rect 353294 204212 353300 204224
rect 353352 204212 353358 204264
rect 372614 204212 372620 204264
rect 372672 204252 372678 204264
rect 376478 204252 376484 204264
rect 372672 204224 376484 204252
rect 372672 204212 372678 204224
rect 376478 204212 376484 204224
rect 376536 204212 376542 204264
rect 403526 204212 403532 204264
rect 403584 204252 403590 204264
rect 407022 204252 407028 204264
rect 403584 204224 407028 204252
rect 403584 204212 403590 204224
rect 407022 204212 407028 204224
rect 407080 204212 407086 204264
rect 415118 204212 415124 204264
rect 415176 204252 415182 204264
rect 418706 204252 418712 204264
rect 415176 204224 418712 204252
rect 415176 204212 415182 204224
rect 418706 204212 418712 204224
rect 418764 204212 418770 204264
rect 475470 204212 475476 204264
rect 475528 204252 475534 204264
rect 477862 204252 477868 204264
rect 475528 204224 477868 204252
rect 475528 204212 475534 204224
rect 477862 204212 477868 204224
rect 477920 204252 477926 204264
rect 478138 204252 478144 204264
rect 477920 204224 478144 204252
rect 477920 204212 477926 204224
rect 478138 204212 478144 204224
rect 478196 204212 478202 204264
rect 123904 204156 180794 204184
rect 123904 204144 123910 204156
rect 197354 204144 197360 204196
rect 197412 204184 197418 204196
rect 197814 204184 197820 204196
rect 197412 204156 197820 204184
rect 197412 204144 197418 204156
rect 197814 204144 197820 204156
rect 197872 204184 197878 204196
rect 200390 204184 200396 204196
rect 197872 204156 200396 204184
rect 197872 204144 197878 204156
rect 200390 204144 200396 204156
rect 200448 204144 200454 204196
rect 301958 204144 301964 204196
rect 302016 204184 302022 204196
rect 330110 204184 330116 204196
rect 302016 204156 330116 204184
rect 302016 204144 302022 204156
rect 330110 204144 330116 204156
rect 330168 204144 330174 204196
rect 453758 204144 453764 204196
rect 453816 204184 453822 204196
rect 478046 204184 478052 204196
rect 453816 204156 478052 204184
rect 453816 204144 453822 204156
rect 478046 204144 478052 204156
rect 478104 204144 478110 204196
rect 19150 204076 19156 204128
rect 19208 204116 19214 204128
rect 73154 204116 73160 204128
rect 19208 204088 73160 204116
rect 19208 204076 19214 204088
rect 73154 204076 73160 204088
rect 73212 204076 73218 204128
rect 150894 204076 150900 204128
rect 150952 204116 150958 204128
rect 150952 204088 190454 204116
rect 150952 204076 150958 204088
rect 18966 204008 18972 204060
rect 19024 204048 19030 204060
rect 19242 204048 19248 204060
rect 19024 204020 19248 204048
rect 19024 204008 19030 204020
rect 19242 204008 19248 204020
rect 19300 204008 19306 204060
rect 30466 204008 30472 204060
rect 30524 204048 30530 204060
rect 34514 204048 34520 204060
rect 30524 204020 34520 204048
rect 30524 204008 30530 204020
rect 34514 204008 34520 204020
rect 34572 204008 34578 204060
rect 34606 204008 34612 204060
rect 34664 204048 34670 204060
rect 80698 204048 80704 204060
rect 34664 204020 80704 204048
rect 34664 204008 34670 204020
rect 80698 204008 80704 204020
rect 80756 204008 80762 204060
rect 173710 204008 173716 204060
rect 173768 204048 173774 204060
rect 183462 204048 183468 204060
rect 173768 204020 183468 204048
rect 173768 204008 173774 204020
rect 183462 204008 183468 204020
rect 183520 204008 183526 204060
rect 190426 204048 190454 204088
rect 193030 204076 193036 204128
rect 193088 204116 193094 204128
rect 195882 204116 195888 204128
rect 193088 204088 195888 204116
rect 193088 204076 193094 204088
rect 195882 204076 195888 204088
rect 195940 204076 195946 204128
rect 198734 204076 198740 204128
rect 198792 204116 198798 204128
rect 199010 204116 199016 204128
rect 198792 204088 199016 204116
rect 198792 204076 198798 204088
rect 199010 204076 199016 204088
rect 199068 204076 199074 204128
rect 302786 204076 302792 204128
rect 302844 204116 302850 204128
rect 326246 204116 326252 204128
rect 302844 204088 326252 204116
rect 302844 204076 302850 204088
rect 326246 204076 326252 204088
rect 326304 204076 326310 204128
rect 411254 204076 411260 204128
rect 411312 204116 411318 204128
rect 413922 204116 413928 204128
rect 411312 204088 413928 204116
rect 411312 204076 411318 204088
rect 413922 204076 413928 204088
rect 413980 204076 413986 204128
rect 457622 204076 457628 204128
rect 457680 204116 457686 204128
rect 457680 204088 476160 204116
rect 457680 204076 457686 204088
rect 198752 204048 198780 204076
rect 190426 204020 198780 204048
rect 301866 204008 301872 204060
rect 301924 204048 301930 204060
rect 322382 204048 322388 204060
rect 301924 204020 322388 204048
rect 301924 204008 301930 204020
rect 322382 204008 322388 204020
rect 322440 204008 322446 204060
rect 461486 204008 461492 204060
rect 461544 204048 461550 204060
rect 475470 204048 475476 204060
rect 461544 204020 475476 204048
rect 461544 204008 461550 204020
rect 475470 204008 475476 204020
rect 475528 204008 475534 204060
rect 20438 203940 20444 203992
rect 20496 203980 20502 203992
rect 65242 203980 65248 203992
rect 20496 203952 65248 203980
rect 20496 203940 20502 203952
rect 65242 203940 65248 203952
rect 65300 203940 65306 203992
rect 112254 203940 112260 203992
rect 112312 203980 112318 203992
rect 200298 203980 200304 203992
rect 112312 203952 200304 203980
rect 112312 203940 112318 203952
rect 200298 203940 200304 203952
rect 200356 203980 200362 203992
rect 200482 203980 200488 203992
rect 200356 203952 200488 203980
rect 200356 203940 200362 203952
rect 200482 203940 200488 203952
rect 200540 203940 200546 203992
rect 301774 203940 301780 203992
rect 301832 203980 301838 203992
rect 314654 203980 314660 203992
rect 301832 203952 314660 203980
rect 301832 203940 301838 203952
rect 314654 203940 314660 203952
rect 314712 203940 314718 203992
rect 465350 203940 465356 203992
rect 465408 203980 465414 203992
rect 465408 203952 473032 203980
rect 465408 203940 465414 203952
rect 19242 203872 19248 203924
rect 19300 203912 19306 203924
rect 61378 203912 61384 203924
rect 19300 203884 61384 203912
rect 19300 203872 19306 203884
rect 61378 203872 61384 203884
rect 61436 203872 61442 203924
rect 302050 203872 302056 203924
rect 302108 203912 302114 203924
rect 310790 203912 310796 203924
rect 302108 203884 310796 203912
rect 302108 203872 302114 203884
rect 310790 203872 310796 203884
rect 310848 203872 310854 203924
rect 312538 203872 312544 203924
rect 312596 203912 312602 203924
rect 313274 203912 313280 203924
rect 312596 203884 313280 203912
rect 312596 203872 312602 203884
rect 313274 203872 313280 203884
rect 313332 203912 313338 203924
rect 384206 203912 384212 203924
rect 313332 203884 384212 203912
rect 313332 203872 313338 203884
rect 384206 203872 384212 203884
rect 384264 203872 384270 203924
rect 449894 203872 449900 203924
rect 449952 203912 449958 203924
rect 473004 203912 473032 203952
rect 473078 203940 473084 203992
rect 473136 203980 473142 203992
rect 476022 203980 476028 203992
rect 473136 203952 476028 203980
rect 473136 203940 473142 203952
rect 476022 203940 476028 203952
rect 476080 203940 476086 203992
rect 476132 203980 476160 204088
rect 476942 204076 476948 204128
rect 477000 204116 477006 204128
rect 480530 204116 480536 204128
rect 477000 204088 480536 204116
rect 477000 204076 477006 204088
rect 480530 204076 480536 204088
rect 480588 204076 480594 204128
rect 478966 203980 478972 203992
rect 476132 203952 478972 203980
rect 478966 203940 478972 203952
rect 479024 203940 479030 203992
rect 478874 203912 478880 203924
rect 449952 203884 470594 203912
rect 473004 203884 478880 203912
rect 449952 203872 449958 203884
rect 17862 203804 17868 203856
rect 17920 203844 17926 203856
rect 84562 203844 84568 203856
rect 17920 203816 84568 203844
rect 17920 203804 17926 203816
rect 84562 203804 84568 203816
rect 84620 203804 84626 203856
rect 181806 203804 181812 203856
rect 181864 203844 181870 203856
rect 187878 203844 187884 203856
rect 181864 203816 187884 203844
rect 181864 203804 181870 203816
rect 187878 203804 187884 203816
rect 187936 203804 187942 203856
rect 470566 203844 470594 203884
rect 478874 203872 478880 203884
rect 478932 203872 478938 203924
rect 479150 203844 479156 203856
rect 470566 203816 479156 203844
rect 479150 203804 479156 203816
rect 479208 203804 479214 203856
rect 28902 203736 28908 203788
rect 28960 203776 28966 203788
rect 34606 203776 34612 203788
rect 28960 203748 34612 203776
rect 28960 203736 28966 203748
rect 34606 203736 34612 203748
rect 34664 203736 34670 203788
rect 34698 203736 34704 203788
rect 34756 203776 34762 203788
rect 38194 203776 38200 203788
rect 34756 203748 38200 203776
rect 34756 203736 34762 203748
rect 38194 203736 38200 203748
rect 38252 203736 38258 203788
rect 127710 203668 127716 203720
rect 127768 203708 127774 203720
rect 200758 203708 200764 203720
rect 127768 203680 200764 203708
rect 127768 203668 127774 203680
rect 200758 203668 200764 203680
rect 200816 203708 200822 203720
rect 201862 203708 201868 203720
rect 200816 203680 201868 203708
rect 200816 203668 200822 203680
rect 201862 203668 201868 203680
rect 201920 203668 201926 203720
rect 139302 203600 139308 203652
rect 139360 203640 139366 203652
rect 240134 203640 240140 203652
rect 139360 203612 240140 203640
rect 139360 203600 139366 203612
rect 240134 203600 240140 203612
rect 240192 203600 240198 203652
rect 269114 203600 269120 203652
rect 269172 203640 269178 203652
rect 372614 203640 372620 203652
rect 269172 203612 372620 203640
rect 269172 203600 269178 203612
rect 372614 203600 372620 203612
rect 372672 203600 372678 203652
rect 189534 203532 189540 203584
rect 189592 203572 189598 203584
rect 300118 203572 300124 203584
rect 189592 203544 300124 203572
rect 189592 203532 189598 203544
rect 300118 203532 300124 203544
rect 300176 203532 300182 203584
rect 469214 203532 469220 203584
rect 469272 203572 469278 203584
rect 481910 203572 481916 203584
rect 469272 203544 481916 203572
rect 469272 203532 469278 203544
rect 481910 203532 481916 203544
rect 481968 203532 481974 203584
rect 185670 203192 185676 203244
rect 185728 203232 185734 203244
rect 188798 203232 188804 203244
rect 185728 203204 188804 203232
rect 185728 203192 185734 203204
rect 188798 203192 188804 203204
rect 188856 203192 188862 203244
rect 17770 202852 17776 202904
rect 17828 202892 17834 202904
rect 22370 202892 22376 202904
rect 17828 202864 22376 202892
rect 17828 202852 17834 202864
rect 22370 202852 22376 202864
rect 22428 202852 22434 202904
rect 39022 202852 39028 202904
rect 39080 202892 39086 202904
rect 42058 202892 42064 202904
rect 39080 202864 42064 202892
rect 39080 202852 39086 202864
rect 42058 202852 42064 202864
rect 42116 202852 42122 202904
rect 399662 202852 399668 202904
rect 399720 202892 399726 202904
rect 399720 202864 402974 202892
rect 399720 202852 399726 202864
rect 22002 202784 22008 202836
rect 22060 202824 22066 202836
rect 22738 202824 22744 202836
rect 22060 202796 22744 202824
rect 22060 202784 22066 202796
rect 22738 202784 22744 202796
rect 22796 202784 22802 202836
rect 53834 202824 53840 202836
rect 23676 202796 53840 202824
rect 21910 202716 21916 202768
rect 21968 202756 21974 202768
rect 23676 202756 23704 202796
rect 53834 202784 53840 202796
rect 53892 202784 53898 202836
rect 166350 202784 166356 202836
rect 166408 202824 166414 202836
rect 197906 202824 197912 202836
rect 166408 202796 197912 202824
rect 166408 202784 166414 202796
rect 197906 202784 197912 202796
rect 197964 202784 197970 202836
rect 402946 202824 402974 202864
rect 407390 202852 407396 202904
rect 407448 202892 407454 202904
rect 410794 202892 410800 202904
rect 407448 202864 410800 202892
rect 407448 202852 407454 202864
rect 410794 202852 410800 202864
rect 410852 202852 410858 202904
rect 477494 202824 477500 202836
rect 402946 202796 477500 202824
rect 477494 202784 477500 202796
rect 477552 202784 477558 202836
rect 21968 202728 23704 202756
rect 21968 202716 21974 202728
rect 23750 202716 23756 202768
rect 23808 202756 23814 202768
rect 49786 202756 49792 202768
rect 23808 202728 49792 202756
rect 23808 202716 23814 202728
rect 49786 202716 49792 202728
rect 49844 202716 49850 202768
rect 170214 202716 170220 202768
rect 170272 202756 170278 202768
rect 198826 202756 198832 202768
rect 170272 202728 198832 202756
rect 170272 202716 170278 202728
rect 198826 202716 198832 202728
rect 198884 202716 198890 202768
rect 20530 202648 20536 202700
rect 20588 202688 20594 202700
rect 45922 202688 45928 202700
rect 20588 202660 45928 202688
rect 20588 202648 20594 202660
rect 45922 202648 45928 202660
rect 45980 202648 45986 202700
rect 187878 202648 187884 202700
rect 187936 202688 187942 202700
rect 197354 202688 197360 202700
rect 187936 202660 197360 202688
rect 187936 202648 187942 202660
rect 197354 202648 197360 202660
rect 197412 202648 197418 202700
rect 20622 202580 20628 202632
rect 20680 202620 20686 202632
rect 22186 202620 22192 202632
rect 20680 202592 22192 202620
rect 20680 202580 20686 202592
rect 22186 202580 22192 202592
rect 22244 202620 22250 202632
rect 39022 202620 39028 202632
rect 22244 202592 39028 202620
rect 22244 202580 22250 202592
rect 39022 202580 39028 202592
rect 39080 202580 39086 202632
rect 20162 202512 20168 202564
rect 20220 202552 20226 202564
rect 23750 202552 23756 202564
rect 20220 202524 23756 202552
rect 20220 202512 20226 202524
rect 23750 202512 23756 202524
rect 23808 202512 23814 202564
rect 198090 202240 198096 202292
rect 198148 202240 198154 202292
rect 197354 202172 197360 202224
rect 197412 202212 197418 202224
rect 198108 202212 198136 202240
rect 200482 202212 200488 202224
rect 197412 202184 200488 202212
rect 197412 202172 197418 202184
rect 200482 202172 200488 202184
rect 200540 202172 200546 202224
rect 188798 202104 188804 202156
rect 188856 202144 188862 202156
rect 198090 202144 198096 202156
rect 188856 202116 198096 202144
rect 188856 202104 188862 202116
rect 198090 202104 198096 202116
rect 198148 202144 198154 202156
rect 200206 202144 200212 202156
rect 198148 202116 200212 202144
rect 198148 202104 198154 202116
rect 200206 202104 200212 202116
rect 200264 202104 200270 202156
rect 22738 202036 22744 202088
rect 22796 202076 22802 202088
rect 34698 202076 34704 202088
rect 22796 202048 34704 202076
rect 22796 202036 22802 202048
rect 34698 202036 34704 202048
rect 34756 202036 34762 202088
rect 135070 201492 135076 201544
rect 135128 201532 135134 201544
rect 135128 201504 137968 201532
rect 135128 201492 135134 201504
rect 137940 201464 137968 201504
rect 198642 201464 198648 201476
rect 137940 201436 198648 201464
rect 198642 201424 198648 201436
rect 198700 201424 198706 201476
rect 297726 201424 297732 201476
rect 297784 201464 297790 201476
rect 368750 201464 368756 201476
rect 297784 201436 368756 201464
rect 297784 201424 297790 201436
rect 368750 201424 368756 201436
rect 368808 201424 368814 201476
rect 395798 201424 395804 201476
rect 395856 201464 395862 201476
rect 483198 201464 483204 201476
rect 395856 201436 483204 201464
rect 395856 201424 395862 201436
rect 483198 201424 483204 201436
rect 483256 201424 483262 201476
rect 410794 201356 410800 201408
rect 410852 201396 410858 201408
rect 484394 201396 484400 201408
rect 410852 201368 484400 201396
rect 410852 201356 410858 201368
rect 484394 201356 484400 201368
rect 484452 201356 484458 201408
rect 413922 201288 413928 201340
rect 413980 201328 413986 201340
rect 484578 201328 484584 201340
rect 413980 201300 484584 201328
rect 413980 201288 413986 201300
rect 484578 201288 484584 201300
rect 484636 201288 484642 201340
rect 484578 200744 484584 200796
rect 484636 200784 484642 200796
rect 485866 200784 485872 200796
rect 484636 200756 485872 200784
rect 484636 200744 484642 200756
rect 485866 200744 485872 200756
rect 485924 200744 485930 200796
rect 483198 200608 483204 200660
rect 483256 200648 483262 200660
rect 484486 200648 484492 200660
rect 483256 200620 484492 200648
rect 483256 200608 483262 200620
rect 484486 200608 484492 200620
rect 484544 200608 484550 200660
rect 296530 200132 296536 200184
rect 296588 200172 296594 200184
rect 297726 200172 297732 200184
rect 296588 200144 297732 200172
rect 296588 200132 296594 200144
rect 297726 200132 297732 200144
rect 297784 200132 297790 200184
rect 20070 200064 20076 200116
rect 20128 200104 20134 200116
rect 107654 200104 107660 200116
rect 20128 200076 107660 200104
rect 20128 200064 20134 200076
rect 107654 200064 107660 200076
rect 107712 200064 107718 200116
rect 16482 199384 16488 199436
rect 16540 199424 16546 199436
rect 17678 199424 17684 199436
rect 16540 199396 17684 199424
rect 16540 199384 16546 199396
rect 17678 199384 17684 199396
rect 17736 199424 17742 199436
rect 99374 199424 99380 199436
rect 17736 199396 99380 199424
rect 17736 199384 17742 199396
rect 99374 199384 99380 199396
rect 99432 199384 99438 199436
rect 18874 198704 18880 198756
rect 18932 198744 18938 198756
rect 20070 198744 20076 198756
rect 18932 198716 20076 198744
rect 18932 198704 18938 198716
rect 20070 198704 20076 198716
rect 20128 198704 20134 198756
rect 252554 189728 252560 189780
rect 252612 189768 252618 189780
rect 418154 189768 418160 189780
rect 252612 189740 418160 189768
rect 252612 189728 252618 189740
rect 418154 189728 418160 189740
rect 418212 189728 418218 189780
rect 118694 188980 118700 189032
rect 118752 189020 118758 189032
rect 203058 189020 203064 189032
rect 118752 188992 203064 189020
rect 118752 188980 118758 188992
rect 203058 188980 203064 188992
rect 203116 188980 203122 189032
rect 131114 188300 131120 188352
rect 131172 188340 131178 188352
rect 202138 188340 202144 188352
rect 131172 188312 202144 188340
rect 131172 188300 131178 188312
rect 202138 188300 202144 188312
rect 202196 188340 202202 188352
rect 203150 188340 203156 188352
rect 202196 188312 203156 188340
rect 202196 188300 202202 188312
rect 203150 188300 203156 188312
rect 203208 188300 203214 188352
rect 2774 187960 2780 188012
rect 2832 188000 2838 188012
rect 4890 188000 4896 188012
rect 2832 187972 4896 188000
rect 2832 187960 2838 187972
rect 4890 187960 4896 187972
rect 4948 187960 4954 188012
rect 299290 187620 299296 187672
rect 299348 187660 299354 187672
rect 360194 187660 360200 187672
rect 299348 187632 360200 187660
rect 299348 187620 299354 187632
rect 360194 187620 360200 187632
rect 360252 187620 360258 187672
rect 302142 187552 302148 187604
rect 302200 187592 302206 187604
rect 349154 187592 349160 187604
rect 302200 187564 349160 187592
rect 302200 187552 302206 187564
rect 349154 187552 349160 187564
rect 349212 187552 349218 187604
rect 195974 187008 195980 187060
rect 196032 187048 196038 187060
rect 300210 187048 300216 187060
rect 196032 187020 300216 187048
rect 196032 187008 196038 187020
rect 300210 187008 300216 187020
rect 300268 187008 300274 187060
rect 95878 186940 95884 186992
rect 95936 186980 95942 186992
rect 256694 186980 256700 186992
rect 95936 186952 256700 186980
rect 95936 186940 95942 186952
rect 256694 186940 256700 186952
rect 256752 186940 256758 186992
rect 298002 186940 298008 186992
rect 298060 186980 298066 186992
rect 312538 186980 312544 186992
rect 298060 186952 312544 186980
rect 298060 186940 298066 186952
rect 312538 186940 312544 186952
rect 312596 186940 312602 186992
rect 3326 149336 3332 149388
rect 3384 149376 3390 149388
rect 8938 149376 8944 149388
rect 3384 149348 8944 149376
rect 3384 149336 3390 149348
rect 8938 149336 8944 149348
rect 8996 149336 9002 149388
rect 2774 136688 2780 136740
rect 2832 136728 2838 136740
rect 5166 136728 5172 136740
rect 2832 136700 5172 136728
rect 2832 136688 2838 136700
rect 5166 136688 5172 136700
rect 5224 136688 5230 136740
rect 3326 110440 3332 110492
rect 3384 110480 3390 110492
rect 20898 110480 20904 110492
rect 3384 110452 20904 110480
rect 3384 110440 3390 110452
rect 20898 110440 20904 110452
rect 20956 110440 20962 110492
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 20898 84232 20904 84244
rect 3384 84204 20904 84232
rect 3384 84192 3390 84204
rect 20898 84192 20904 84204
rect 20956 84192 20962 84244
rect 20898 79296 20904 79348
rect 20956 79336 20962 79348
rect 21634 79336 21640 79348
rect 20956 79308 21640 79336
rect 20956 79296 20962 79308
rect 21634 79296 21640 79308
rect 21692 79296 21698 79348
rect 301774 78344 301780 78396
rect 301832 78384 301838 78396
rect 314746 78384 314752 78396
rect 301832 78356 314752 78384
rect 301832 78344 301838 78356
rect 314746 78344 314752 78356
rect 314804 78344 314810 78396
rect 302694 78276 302700 78328
rect 302752 78316 302758 78328
rect 317414 78316 317420 78328
rect 302752 78288 317420 78316
rect 302752 78276 302758 78288
rect 317414 78276 317420 78288
rect 317472 78316 317478 78328
rect 318150 78316 318156 78328
rect 317472 78288 318156 78316
rect 317472 78276 317478 78288
rect 318150 78276 318156 78288
rect 318208 78276 318214 78328
rect 301866 78208 301872 78260
rect 301924 78248 301930 78260
rect 316770 78248 316776 78260
rect 301924 78220 316776 78248
rect 301924 78208 301930 78220
rect 316770 78208 316776 78220
rect 316828 78208 316834 78260
rect 302786 78140 302792 78192
rect 302844 78180 302850 78192
rect 318794 78180 318800 78192
rect 302844 78152 318800 78180
rect 302844 78140 302850 78152
rect 318794 78140 318800 78152
rect 318852 78140 318858 78192
rect 430666 78140 430672 78192
rect 430724 78180 430730 78192
rect 478230 78180 478236 78192
rect 430724 78152 478236 78180
rect 430724 78140 430730 78152
rect 478230 78140 478236 78152
rect 478288 78140 478294 78192
rect 301958 78072 301964 78124
rect 302016 78112 302022 78124
rect 329834 78112 329840 78124
rect 302016 78084 329840 78112
rect 302016 78072 302022 78084
rect 329834 78072 329840 78084
rect 329892 78072 329898 78124
rect 394694 78072 394700 78124
rect 394752 78112 394758 78124
rect 480530 78112 480536 78124
rect 394752 78084 480536 78112
rect 394752 78072 394758 78084
rect 480530 78072 480536 78084
rect 480588 78072 480594 78124
rect 18782 78004 18788 78056
rect 18840 78044 18846 78056
rect 88426 78044 88432 78056
rect 18840 78016 88432 78044
rect 18840 78004 18846 78016
rect 88426 78004 88432 78016
rect 88484 78004 88490 78056
rect 191834 78004 191840 78056
rect 191892 78044 191898 78056
rect 192938 78044 192944 78056
rect 191892 78016 192944 78044
rect 191892 78004 191898 78016
rect 192938 78004 192944 78016
rect 192996 78044 193002 78056
rect 200390 78044 200396 78056
rect 192996 78016 200396 78044
rect 192996 78004 193002 78016
rect 200390 78004 200396 78016
rect 200448 78004 200454 78056
rect 307202 78004 307208 78056
rect 307260 78044 307266 78056
rect 479518 78044 479524 78056
rect 307260 78016 479524 78044
rect 307260 78004 307266 78016
rect 479518 78004 479524 78016
rect 479576 78004 479582 78056
rect 16390 77936 16396 77988
rect 16448 77976 16454 77988
rect 103974 77976 103980 77988
rect 16448 77948 103980 77976
rect 16448 77936 16454 77948
rect 103974 77936 103980 77948
rect 104032 77936 104038 77988
rect 185670 77936 185676 77988
rect 185728 77976 185734 77988
rect 198090 77976 198096 77988
rect 185728 77948 198096 77976
rect 185728 77936 185734 77948
rect 198090 77936 198096 77948
rect 198148 77936 198154 77988
rect 302050 77936 302056 77988
rect 302108 77976 302114 77988
rect 310514 77976 310520 77988
rect 302108 77948 310520 77976
rect 302108 77936 302114 77948
rect 310514 77936 310520 77948
rect 310572 77936 310578 77988
rect 311158 77936 311164 77988
rect 311216 77976 311222 77988
rect 579614 77976 579620 77988
rect 311216 77948 579620 77976
rect 311216 77936 311222 77948
rect 579614 77936 579620 77948
rect 579672 77936 579678 77988
rect 372706 77256 372712 77308
rect 372764 77296 372770 77308
rect 480254 77296 480260 77308
rect 372764 77268 480260 77296
rect 372764 77256 372770 77268
rect 480254 77256 480260 77268
rect 480312 77256 480318 77308
rect 99374 77052 99380 77104
rect 99432 77092 99438 77104
rect 100340 77092 100346 77104
rect 99432 77064 100346 77092
rect 99432 77052 99438 77064
rect 100340 77052 100346 77064
rect 100398 77052 100404 77104
rect 283834 76508 283840 76560
rect 283892 76548 283898 76560
rect 369854 76548 369860 76560
rect 283892 76520 369860 76548
rect 283892 76508 283898 76520
rect 369854 76508 369860 76520
rect 369912 76508 369918 76560
rect 17678 75964 17684 76016
rect 17736 76004 17742 76016
rect 99374 76004 99380 76016
rect 17736 75976 99380 76004
rect 17736 75964 17742 75976
rect 99374 75964 99380 75976
rect 99432 75964 99438 76016
rect 18874 75896 18880 75948
rect 18932 75936 18938 75948
rect 108298 75936 108304 75948
rect 18932 75908 108304 75936
rect 18932 75896 18938 75908
rect 108298 75896 108304 75908
rect 108356 75896 108362 75948
rect 422846 75896 422852 75948
rect 422904 75936 422910 75948
rect 483290 75936 483296 75948
rect 422904 75908 483296 75936
rect 422904 75896 422910 75908
rect 483290 75896 483296 75908
rect 483348 75896 483354 75948
rect 19058 75828 19064 75880
rect 19116 75868 19122 75880
rect 76834 75868 76840 75880
rect 19116 75840 76840 75868
rect 19116 75828 19122 75840
rect 76834 75828 76840 75840
rect 76892 75828 76898 75880
rect 92934 75828 92940 75880
rect 92992 75868 92998 75880
rect 96430 75868 96436 75880
rect 92992 75840 96436 75868
rect 92992 75828 92998 75840
rect 96430 75828 96436 75840
rect 96488 75828 96494 75880
rect 150894 75828 150900 75880
rect 150952 75868 150958 75880
rect 199010 75868 199016 75880
rect 150952 75840 199016 75868
rect 150952 75828 150958 75840
rect 199010 75828 199016 75840
rect 199068 75828 199074 75880
rect 300670 75828 300676 75880
rect 300728 75868 300734 75880
rect 340966 75868 340972 75880
rect 300728 75840 340972 75868
rect 300728 75828 300734 75840
rect 340966 75828 340972 75840
rect 341024 75828 341030 75880
rect 372614 75828 372620 75880
rect 372672 75868 372678 75880
rect 376478 75868 376484 75880
rect 372672 75840 376484 75868
rect 372672 75828 372678 75840
rect 376478 75828 376484 75840
rect 376536 75828 376542 75880
rect 19150 75760 19156 75812
rect 19208 75800 19214 75812
rect 73338 75800 73344 75812
rect 19208 75772 73344 75800
rect 19208 75760 19214 75772
rect 73338 75760 73344 75772
rect 73396 75760 73402 75812
rect 158622 75760 158628 75812
rect 158680 75800 158686 75812
rect 201770 75800 201776 75812
rect 158680 75772 201776 75800
rect 158680 75760 158686 75772
rect 201770 75760 201776 75772
rect 201828 75800 201834 75812
rect 202782 75800 202788 75812
rect 201828 75772 202788 75800
rect 201828 75760 201834 75772
rect 202782 75760 202788 75772
rect 202840 75760 202846 75812
rect 316770 75760 316776 75812
rect 316828 75800 316834 75812
rect 316954 75800 316960 75812
rect 316828 75772 316960 75800
rect 316828 75760 316834 75772
rect 316954 75760 316960 75772
rect 317012 75800 317018 75812
rect 322382 75800 322388 75812
rect 317012 75772 322388 75800
rect 317012 75760 317018 75772
rect 322382 75760 322388 75772
rect 322440 75760 322446 75812
rect 326246 75800 326252 75812
rect 325666 75772 326252 75800
rect 17770 75692 17776 75744
rect 17828 75732 17834 75744
rect 69566 75732 69572 75744
rect 17828 75704 69572 75732
rect 17828 75692 17834 75704
rect 69566 75692 69572 75704
rect 69624 75692 69630 75744
rect 177942 75692 177948 75744
rect 178000 75732 178006 75744
rect 198918 75732 198924 75744
rect 178000 75704 198924 75732
rect 178000 75692 178006 75704
rect 198918 75692 198924 75704
rect 198976 75692 198982 75744
rect 318794 75692 318800 75744
rect 318852 75732 318858 75744
rect 325666 75732 325694 75772
rect 326246 75760 326252 75772
rect 326304 75760 326310 75812
rect 433978 75760 433984 75812
rect 434036 75800 434042 75812
rect 434438 75800 434444 75812
rect 434036 75772 434444 75800
rect 434036 75760 434042 75772
rect 434438 75760 434444 75772
rect 434496 75800 434502 75812
rect 480438 75800 480444 75812
rect 434496 75772 480444 75800
rect 434496 75760 434502 75772
rect 480438 75760 480444 75772
rect 480496 75760 480502 75812
rect 318852 75704 325694 75732
rect 318852 75692 318858 75704
rect 438302 75692 438308 75744
rect 438360 75732 438366 75744
rect 480714 75732 480720 75744
rect 438360 75704 480720 75732
rect 438360 75692 438366 75704
rect 480714 75692 480720 75704
rect 480772 75692 480778 75744
rect 20438 75624 20444 75676
rect 20496 75664 20502 75676
rect 65334 75664 65340 75676
rect 20496 75636 65340 75664
rect 20496 75624 20502 75636
rect 65334 75624 65340 75636
rect 65392 75624 65398 75676
rect 442258 75624 442264 75676
rect 442316 75664 442322 75676
rect 483014 75664 483020 75676
rect 442316 75636 483020 75664
rect 442316 75624 442322 75636
rect 483014 75624 483020 75636
rect 483072 75624 483078 75676
rect 19242 75556 19248 75608
rect 19300 75596 19306 75608
rect 61378 75596 61384 75608
rect 19300 75568 61384 75596
rect 19300 75556 19306 75568
rect 61378 75556 61384 75568
rect 61436 75556 61442 75608
rect 449894 75556 449900 75608
rect 449952 75596 449958 75608
rect 479150 75596 479156 75608
rect 449952 75568 479156 75596
rect 449952 75556 449958 75568
rect 479150 75556 479156 75568
rect 479208 75556 479214 75608
rect 20346 75488 20352 75540
rect 20404 75528 20410 75540
rect 50338 75528 50344 75540
rect 20404 75500 50344 75528
rect 20404 75488 20410 75500
rect 50338 75488 50344 75500
rect 50396 75488 50402 75540
rect 414658 75488 414664 75540
rect 414716 75528 414722 75540
rect 415118 75528 415124 75540
rect 414716 75500 415124 75528
rect 414716 75488 414722 75500
rect 415118 75488 415124 75500
rect 415176 75528 415182 75540
rect 479058 75528 479064 75540
rect 415176 75500 479064 75528
rect 415176 75488 415182 75500
rect 479058 75488 479064 75500
rect 479116 75488 479122 75540
rect 4982 75420 4988 75472
rect 5040 75460 5046 75472
rect 23014 75460 23020 75472
rect 5040 75432 23020 75460
rect 5040 75420 5046 75432
rect 23014 75420 23020 75432
rect 23072 75420 23078 75472
rect 189534 75352 189540 75404
rect 189592 75392 189598 75404
rect 229738 75392 229744 75404
rect 189592 75364 229744 75392
rect 189592 75352 189598 75364
rect 229738 75352 229744 75364
rect 229796 75352 229802 75404
rect 322198 75352 322204 75404
rect 322256 75392 322262 75404
rect 333974 75392 333980 75404
rect 322256 75364 333980 75392
rect 322256 75352 322262 75364
rect 333974 75352 333980 75364
rect 334032 75352 334038 75404
rect 375374 75352 375380 75404
rect 375432 75392 375438 75404
rect 449894 75392 449900 75404
rect 375432 75364 449900 75392
rect 375432 75352 375438 75364
rect 449894 75352 449900 75364
rect 449952 75352 449958 75404
rect 96430 75284 96436 75336
rect 96488 75324 96494 75336
rect 112438 75324 112444 75336
rect 96488 75296 112444 75324
rect 96488 75284 96494 75296
rect 112438 75284 112444 75296
rect 112496 75284 112502 75336
rect 199010 75284 199016 75336
rect 199068 75324 199074 75336
rect 255958 75324 255964 75336
rect 199068 75296 255964 75324
rect 199068 75284 199074 75296
rect 255958 75284 255964 75296
rect 256016 75284 256022 75336
rect 327074 75284 327080 75336
rect 327132 75324 327138 75336
rect 345566 75324 345572 75336
rect 327132 75296 345572 75324
rect 327132 75284 327138 75296
rect 345566 75284 345572 75296
rect 345624 75284 345630 75336
rect 376754 75284 376760 75336
rect 376812 75324 376818 75336
rect 480346 75324 480352 75336
rect 376812 75296 480352 75324
rect 376812 75284 376818 75296
rect 480346 75284 480352 75296
rect 480404 75284 480410 75336
rect 112254 75216 112260 75268
rect 112312 75256 112318 75268
rect 139210 75256 139216 75268
rect 112312 75228 139216 75256
rect 112312 75216 112318 75228
rect 139210 75216 139216 75228
rect 139268 75216 139274 75268
rect 147030 75216 147036 75268
rect 147088 75256 147094 75268
rect 156598 75256 156604 75268
rect 147088 75228 156604 75256
rect 147088 75216 147094 75228
rect 156598 75216 156604 75228
rect 156656 75216 156662 75268
rect 202782 75216 202788 75268
rect 202840 75256 202846 75268
rect 288434 75256 288440 75268
rect 202840 75228 288440 75256
rect 202840 75216 202846 75228
rect 288434 75216 288440 75228
rect 288492 75216 288498 75268
rect 300578 75216 300584 75268
rect 300636 75256 300642 75268
rect 331214 75256 331220 75268
rect 300636 75228 331220 75256
rect 300636 75216 300642 75228
rect 331214 75216 331220 75228
rect 331272 75256 331278 75268
rect 357158 75256 357164 75268
rect 331272 75228 357164 75256
rect 331272 75216 331278 75228
rect 357158 75216 357164 75228
rect 357216 75216 357222 75268
rect 378134 75216 378140 75268
rect 378192 75256 378198 75268
rect 481910 75256 481916 75268
rect 378192 75228 481916 75256
rect 378192 75216 378198 75228
rect 481910 75216 481916 75228
rect 481968 75216 481974 75268
rect 69566 75148 69572 75200
rect 69624 75188 69630 75200
rect 122098 75188 122104 75200
rect 69624 75160 122104 75188
rect 69624 75148 69630 75160
rect 122098 75148 122104 75160
rect 122156 75148 122162 75200
rect 139302 75148 139308 75200
rect 139360 75188 139366 75200
rect 238754 75188 238760 75200
rect 139360 75160 238760 75188
rect 139360 75148 139366 75160
rect 238754 75148 238760 75160
rect 238812 75148 238818 75200
rect 278774 75148 278780 75200
rect 278832 75188 278838 75200
rect 438302 75188 438308 75200
rect 278832 75160 438308 75188
rect 278832 75148 278838 75160
rect 438302 75148 438308 75160
rect 438360 75148 438366 75200
rect 271874 74604 271880 74656
rect 271932 74644 271938 74656
rect 422846 74644 422852 74656
rect 271932 74616 422852 74644
rect 271932 74604 271938 74616
rect 422846 74604 422852 74616
rect 422904 74604 422910 74656
rect 274634 74536 274640 74588
rect 274692 74576 274698 74588
rect 430574 74576 430580 74588
rect 274692 74548 430580 74576
rect 274692 74536 274698 74548
rect 430574 74536 430580 74548
rect 430632 74536 430638 74588
rect 17862 74468 17868 74520
rect 17920 74508 17926 74520
rect 84930 74508 84936 74520
rect 17920 74480 84936 74508
rect 17920 74468 17926 74480
rect 84930 74468 84936 74480
rect 84988 74468 84994 74520
rect 139210 74468 139216 74520
rect 139268 74508 139274 74520
rect 200298 74508 200304 74520
rect 139268 74480 200304 74508
rect 139268 74468 139274 74480
rect 200298 74468 200304 74480
rect 200356 74508 200362 74520
rect 201402 74508 201408 74520
rect 200356 74480 201408 74508
rect 200356 74468 200362 74480
rect 201402 74468 201408 74480
rect 201460 74468 201466 74520
rect 427078 74468 427084 74520
rect 427136 74508 427142 74520
rect 483382 74508 483388 74520
rect 427136 74480 483388 74508
rect 427136 74468 427142 74480
rect 483382 74468 483388 74480
rect 483440 74468 483446 74520
rect 21910 74400 21916 74452
rect 21968 74440 21974 74452
rect 54478 74440 54484 74452
rect 21968 74412 54484 74440
rect 21968 74400 21974 74412
rect 54478 74400 54484 74412
rect 54536 74400 54542 74452
rect 446398 74400 446404 74452
rect 446456 74440 446462 74452
rect 477954 74440 477960 74452
rect 446456 74412 477960 74440
rect 446456 74400 446462 74412
rect 477954 74400 477960 74412
rect 478012 74400 478018 74452
rect 20530 74332 20536 74384
rect 20588 74372 20594 74384
rect 46198 74372 46204 74384
rect 20588 74344 46204 74372
rect 20588 74332 20594 74344
rect 46198 74332 46204 74344
rect 46256 74332 46262 74384
rect 453758 74332 453764 74384
rect 453816 74372 453822 74384
rect 478046 74372 478052 74384
rect 453816 74344 478052 74372
rect 453816 74332 453822 74344
rect 478046 74332 478052 74344
rect 478104 74332 478110 74384
rect 20622 74264 20628 74316
rect 20680 74304 20686 74316
rect 42058 74304 42064 74316
rect 20680 74276 42064 74304
rect 20680 74264 20686 74276
rect 42058 74264 42064 74276
rect 42116 74264 42122 74316
rect 457622 74264 457628 74316
rect 457680 74304 457686 74316
rect 478966 74304 478972 74316
rect 457680 74276 478972 74304
rect 457680 74264 457686 74276
rect 478966 74264 478972 74276
rect 479024 74264 479030 74316
rect 22738 74196 22744 74248
rect 22796 74236 22802 74248
rect 38102 74236 38108 74248
rect 22796 74208 38108 74236
rect 22796 74196 22802 74208
rect 38102 74196 38108 74208
rect 38160 74196 38166 74248
rect 461486 74196 461492 74248
rect 461544 74236 461550 74248
rect 477862 74236 477868 74248
rect 461544 74208 477868 74236
rect 461544 74196 461550 74208
rect 477862 74196 477868 74208
rect 477920 74196 477926 74248
rect 22830 74128 22836 74180
rect 22888 74168 22894 74180
rect 35158 74168 35164 74180
rect 22888 74140 35164 74168
rect 22888 74128 22894 74140
rect 35158 74128 35164 74140
rect 35216 74128 35222 74180
rect 465718 74128 465724 74180
rect 465776 74168 465782 74180
rect 478874 74168 478880 74180
rect 465776 74140 478880 74168
rect 465776 74128 465782 74140
rect 478874 74128 478880 74140
rect 478932 74128 478938 74180
rect 22922 74060 22928 74112
rect 22980 74100 22986 74112
rect 31018 74100 31024 74112
rect 22980 74072 31024 74100
rect 22980 74060 22986 74072
rect 31018 74060 31024 74072
rect 31076 74060 31082 74112
rect 473078 74060 473084 74112
rect 473136 74100 473142 74112
rect 481818 74100 481824 74112
rect 473136 74072 481824 74100
rect 473136 74060 473142 74072
rect 481818 74060 481824 74072
rect 481876 74060 481882 74112
rect 198918 73992 198924 74044
rect 198976 74032 198982 74044
rect 307018 74032 307024 74044
rect 198976 74004 307024 74032
rect 198976 73992 198982 74004
rect 307018 73992 307024 74004
rect 307076 73992 307082 74044
rect 311158 73992 311164 74044
rect 311216 74032 311222 74044
rect 427078 74032 427084 74044
rect 311216 74004 427084 74032
rect 311216 73992 311222 74004
rect 427078 73992 427084 74004
rect 427136 73992 427142 74044
rect 201402 73924 201408 73976
rect 201460 73964 201466 73976
rect 227714 73964 227720 73976
rect 201460 73936 227720 73964
rect 201460 73924 201466 73936
rect 227714 73924 227720 73936
rect 227772 73924 227778 73976
rect 298646 73924 298652 73976
rect 298704 73964 298710 73976
rect 461486 73964 461492 73976
rect 298704 73936 461492 73964
rect 298704 73924 298710 73936
rect 461486 73924 461492 73936
rect 461544 73924 461550 73976
rect 212626 73856 212632 73908
rect 212684 73896 212690 73908
rect 395798 73896 395804 73908
rect 212684 73868 395804 73896
rect 212684 73856 212690 73868
rect 395798 73856 395804 73868
rect 395856 73856 395862 73908
rect 73338 73788 73344 73840
rect 73396 73828 73402 73840
rect 356698 73828 356704 73840
rect 73396 73800 356704 73828
rect 73396 73788 73402 73800
rect 356698 73788 356704 73800
rect 356756 73788 356762 73840
rect 119890 73108 119896 73160
rect 119948 73148 119954 73160
rect 203058 73148 203064 73160
rect 119948 73120 203064 73148
rect 119948 73108 119954 73120
rect 203058 73108 203064 73120
rect 203116 73108 203122 73160
rect 403618 73108 403624 73160
rect 403676 73148 403682 73160
rect 481726 73148 481732 73160
rect 403676 73120 481732 73148
rect 403676 73108 403682 73120
rect 481726 73108 481732 73120
rect 481784 73108 481790 73160
rect 173802 73040 173808 73092
rect 173860 73080 173866 73092
rect 197998 73080 198004 73092
rect 173860 73052 198004 73080
rect 173860 73040 173866 73052
rect 197998 73040 198004 73052
rect 198056 73040 198062 73092
rect 407758 73040 407764 73092
rect 407816 73080 407822 73092
rect 484394 73080 484400 73092
rect 407816 73052 484400 73080
rect 407816 73040 407822 73052
rect 484394 73040 484400 73052
rect 484452 73040 484458 73092
rect 411254 72972 411260 73024
rect 411312 73012 411318 73024
rect 411898 73012 411904 73024
rect 411312 72984 411904 73012
rect 411312 72972 411318 72984
rect 411898 72972 411904 72984
rect 411956 73012 411962 73024
rect 485866 73012 485872 73024
rect 411956 72984 485872 73012
rect 411956 72972 411962 72984
rect 485866 72972 485872 72984
rect 485924 72972 485930 73024
rect 203058 72632 203064 72684
rect 203116 72672 203122 72684
rect 230842 72672 230848 72684
rect 203116 72644 230848 72672
rect 203116 72632 203122 72644
rect 230842 72632 230848 72644
rect 230900 72632 230906 72684
rect 293954 72632 293960 72684
rect 294012 72672 294018 72684
rect 375374 72672 375380 72684
rect 294012 72644 375380 72672
rect 294012 72632 294018 72644
rect 375374 72632 375380 72644
rect 375432 72632 375438 72684
rect 197998 72564 198004 72616
rect 198056 72604 198062 72616
rect 305362 72604 305368 72616
rect 198056 72576 305368 72604
rect 198056 72564 198062 72576
rect 305362 72564 305368 72576
rect 305420 72564 305426 72616
rect 330294 72564 330300 72616
rect 330352 72604 330358 72616
rect 353294 72604 353300 72616
rect 330352 72576 353300 72604
rect 330352 72564 330358 72576
rect 353294 72564 353300 72576
rect 353352 72564 353358 72616
rect 104434 72496 104440 72548
rect 104492 72536 104498 72548
rect 224218 72536 224224 72548
rect 104492 72508 224224 72536
rect 104492 72496 104498 72508
rect 224218 72496 224224 72508
rect 224276 72496 224282 72548
rect 254026 72496 254032 72548
rect 254084 72536 254090 72548
rect 418982 72536 418988 72548
rect 254084 72508 418988 72536
rect 254084 72496 254090 72508
rect 418982 72496 418988 72508
rect 419040 72496 419046 72548
rect 38102 72428 38108 72480
rect 38160 72468 38166 72480
rect 340874 72468 340880 72480
rect 38160 72440 340880 72468
rect 38160 72428 38166 72440
rect 340874 72428 340880 72440
rect 340932 72428 340938 72480
rect 131482 71680 131488 71732
rect 131540 71720 131546 71732
rect 202138 71720 202144 71732
rect 131540 71692 202144 71720
rect 131540 71680 131546 71692
rect 202138 71680 202144 71692
rect 202196 71720 202202 71732
rect 202782 71720 202788 71732
rect 202196 71692 202788 71720
rect 202196 71680 202202 71692
rect 202782 71680 202788 71692
rect 202840 71680 202846 71732
rect 299382 71680 299388 71732
rect 299440 71720 299446 71732
rect 329834 71720 329840 71732
rect 299440 71692 329840 71720
rect 299440 71680 299446 71692
rect 329834 71680 329840 71692
rect 329892 71720 329898 71732
rect 330294 71720 330300 71732
rect 329892 71692 330300 71720
rect 329892 71680 329898 71692
rect 330294 71680 330300 71692
rect 330352 71680 330358 71732
rect 202782 71204 202788 71256
rect 202840 71244 202846 71256
rect 235994 71244 236000 71256
rect 202840 71216 236000 71244
rect 202840 71204 202846 71216
rect 235994 71204 236000 71216
rect 236052 71204 236058 71256
rect 270586 71204 270592 71256
rect 270644 71244 270650 71256
rect 372614 71244 372620 71256
rect 270644 71216 372620 71244
rect 270644 71204 270650 71216
rect 372614 71204 372620 71216
rect 372672 71204 372678 71256
rect 203058 71136 203064 71188
rect 203116 71176 203122 71188
rect 473078 71176 473084 71188
rect 203116 71148 473084 71176
rect 203116 71136 203122 71148
rect 473078 71136 473084 71148
rect 473136 71136 473142 71188
rect 88978 71068 88984 71120
rect 89036 71108 89042 71120
rect 363322 71108 363328 71120
rect 89036 71080 363328 71108
rect 89036 71068 89042 71080
rect 363322 71068 363328 71080
rect 363380 71068 363386 71120
rect 81250 71000 81256 71052
rect 81308 71040 81314 71052
rect 360194 71040 360200 71052
rect 81308 71012 360200 71040
rect 81308 71000 81314 71012
rect 360194 71000 360200 71012
rect 360252 71000 360258 71052
rect 127618 70320 127624 70372
rect 127676 70360 127682 70372
rect 200758 70360 200764 70372
rect 127676 70332 200764 70360
rect 127676 70320 127682 70332
rect 200758 70320 200764 70332
rect 200816 70360 200822 70372
rect 201402 70360 201408 70372
rect 200816 70332 201408 70360
rect 200816 70320 200822 70332
rect 201402 70320 201408 70332
rect 201460 70320 201466 70372
rect 170122 70252 170128 70304
rect 170180 70292 170186 70304
rect 198826 70292 198832 70304
rect 170180 70264 198832 70292
rect 170180 70252 170186 70264
rect 198826 70252 198832 70264
rect 198884 70292 198890 70304
rect 199378 70292 199384 70304
rect 198884 70264 199384 70292
rect 198884 70252 198890 70264
rect 199378 70252 199384 70264
rect 199436 70252 199442 70304
rect 199378 69776 199384 69828
rect 199436 69816 199442 69828
rect 303706 69816 303712 69828
rect 199436 69788 303712 69816
rect 199436 69776 199442 69788
rect 303706 69776 303712 69788
rect 303764 69776 303770 69828
rect 201402 69708 201408 69760
rect 201460 69748 201466 69760
rect 234154 69748 234160 69760
rect 201460 69720 234160 69748
rect 201460 69708 201466 69720
rect 234154 69708 234160 69720
rect 234212 69708 234218 69760
rect 297082 69708 297088 69760
rect 297140 69748 297146 69760
rect 457622 69748 457628 69760
rect 297140 69720 457628 69748
rect 297140 69708 297146 69720
rect 457622 69708 457628 69720
rect 457680 69708 457686 69760
rect 76834 69640 76840 69692
rect 76892 69680 76898 69692
rect 358354 69680 358360 69692
rect 76892 69652 358360 69680
rect 76892 69640 76898 69652
rect 358354 69640 358360 69652
rect 358412 69640 358418 69692
rect 135162 68960 135168 69012
rect 135220 69000 135226 69012
rect 198734 69000 198740 69012
rect 135220 68972 198740 69000
rect 135220 68960 135226 68972
rect 198734 68960 198740 68972
rect 198792 68960 198798 69012
rect 300762 68960 300768 69012
rect 300820 69000 300826 69012
rect 327074 69000 327080 69012
rect 300820 68972 327080 69000
rect 300820 68960 300826 68972
rect 327074 68960 327080 68972
rect 327132 68960 327138 69012
rect 166258 68892 166264 68944
rect 166316 68932 166322 68944
rect 197354 68932 197360 68944
rect 166316 68904 197360 68932
rect 166316 68892 166322 68904
rect 197354 68892 197360 68904
rect 197412 68892 197418 68944
rect 198734 68552 198740 68604
rect 198792 68592 198798 68604
rect 237466 68592 237472 68604
rect 198792 68564 237472 68592
rect 198792 68552 198798 68564
rect 237466 68552 237472 68564
rect 237524 68552 237530 68604
rect 197354 68484 197360 68536
rect 197412 68524 197418 68536
rect 197906 68524 197912 68536
rect 197412 68496 197912 68524
rect 197412 68484 197418 68496
rect 197906 68484 197912 68496
rect 197964 68524 197970 68536
rect 302234 68524 302240 68536
rect 197964 68496 302240 68524
rect 197964 68484 197970 68496
rect 302234 68484 302240 68496
rect 302292 68484 302298 68536
rect 233878 68416 233884 68468
rect 233936 68456 233942 68468
rect 368566 68456 368572 68468
rect 233936 68428 368572 68456
rect 233936 68416 233942 68428
rect 368566 68416 368572 68428
rect 368624 68416 368630 68468
rect 108298 68348 108304 68400
rect 108356 68388 108362 68400
rect 225874 68388 225880 68400
rect 108356 68360 225880 68388
rect 108356 68348 108362 68360
rect 225874 68348 225880 68360
rect 225932 68348 225938 68400
rect 295426 68348 295432 68400
rect 295484 68388 295490 68400
rect 453758 68388 453764 68400
rect 295484 68360 453764 68388
rect 295484 68348 295490 68360
rect 453758 68348 453764 68360
rect 453816 68348 453822 68400
rect 84930 68280 84936 68332
rect 84988 68320 84994 68332
rect 361666 68320 361672 68332
rect 84988 68292 361672 68320
rect 84988 68280 84994 68292
rect 361666 68280 361672 68292
rect 361724 68280 361730 68332
rect 302878 67532 302884 67584
rect 302936 67572 302942 67584
rect 322198 67572 322204 67584
rect 302936 67544 322204 67572
rect 302936 67532 302942 67544
rect 322198 67532 322204 67544
rect 322256 67532 322262 67584
rect 112438 66988 112444 67040
rect 112496 67028 112502 67040
rect 255682 67028 255688 67040
rect 112496 67000 255688 67028
rect 112496 66988 112502 67000
rect 255682 66988 255688 67000
rect 255740 66988 255746 67040
rect 255958 66988 255964 67040
rect 256016 67028 256022 67040
rect 285674 67028 285680 67040
rect 256016 67000 285680 67028
rect 256016 66988 256022 67000
rect 285674 66988 285680 67000
rect 285732 66988 285738 67040
rect 302142 66988 302148 67040
rect 302200 67028 302206 67040
rect 328546 67028 328552 67040
rect 302200 67000 328552 67028
rect 302200 66988 302206 67000
rect 328546 66988 328552 67000
rect 328604 67028 328610 67040
rect 349154 67028 349160 67040
rect 328604 67000 349160 67028
rect 328604 66988 328610 67000
rect 349154 66988 349160 67000
rect 349212 66988 349218 67040
rect 122098 66920 122104 66972
rect 122156 66960 122162 66972
rect 355042 66960 355048 66972
rect 122156 66932 355048 66960
rect 122156 66920 122162 66932
rect 355042 66920 355048 66932
rect 355100 66920 355106 66972
rect 54478 66852 54484 66904
rect 54536 66892 54542 66904
rect 348418 66892 348424 66904
rect 54536 66864 348424 66892
rect 54536 66852 54542 66864
rect 348418 66852 348424 66864
rect 348476 66852 348482 66904
rect 142154 66172 142160 66224
rect 142212 66212 142218 66224
rect 201586 66212 201592 66224
rect 142212 66184 201592 66212
rect 142212 66172 142218 66184
rect 201586 66172 201592 66184
rect 201644 66212 201650 66224
rect 202782 66212 202788 66224
rect 201644 66184 202788 66212
rect 201644 66172 201650 66184
rect 202782 66172 202788 66184
rect 202840 66172 202846 66224
rect 202782 65696 202788 65748
rect 202840 65736 202846 65748
rect 282178 65736 282184 65748
rect 202840 65708 282184 65736
rect 202840 65696 202846 65708
rect 282178 65696 282184 65708
rect 282236 65696 282242 65748
rect 292114 65696 292120 65748
rect 292172 65736 292178 65748
rect 446398 65736 446404 65748
rect 292172 65708 446404 65736
rect 292172 65696 292178 65708
rect 446398 65696 446404 65708
rect 446456 65696 446462 65748
rect 220906 65628 220912 65680
rect 220964 65668 220970 65680
rect 414658 65668 414664 65680
rect 220964 65640 414664 65668
rect 220964 65628 220970 65640
rect 414658 65628 414664 65640
rect 414716 65628 414722 65680
rect 46198 65560 46204 65612
rect 46256 65600 46262 65612
rect 345106 65600 345112 65612
rect 46256 65572 345112 65600
rect 46256 65560 46262 65572
rect 345106 65560 345112 65572
rect 345164 65560 345170 65612
rect 31018 65492 31024 65544
rect 31076 65532 31082 65544
rect 338482 65532 338488 65544
rect 31076 65504 338488 65532
rect 31076 65492 31082 65504
rect 338482 65492 338488 65504
rect 338540 65492 338546 65544
rect 300026 64812 300032 64864
rect 300084 64852 300090 64864
rect 387794 64852 387800 64864
rect 300084 64824 387800 64852
rect 300084 64812 300090 64824
rect 387794 64812 387800 64824
rect 387852 64812 387858 64864
rect 299290 64336 299296 64388
rect 299348 64376 299354 64388
rect 333514 64376 333520 64388
rect 299348 64348 333520 64376
rect 299348 64336 299354 64348
rect 333514 64336 333520 64348
rect 333572 64376 333578 64388
rect 360286 64376 360292 64388
rect 333572 64348 360292 64376
rect 333572 64336 333578 64348
rect 360286 64336 360292 64348
rect 360344 64336 360350 64388
rect 57238 64268 57244 64320
rect 57296 64308 57302 64320
rect 332594 64308 332600 64320
rect 57296 64280 332600 64308
rect 57296 64268 57302 64280
rect 332594 64268 332600 64280
rect 332652 64268 332658 64320
rect 65518 64200 65524 64252
rect 65576 64240 65582 64252
rect 353386 64240 353392 64252
rect 65576 64212 353392 64240
rect 65576 64200 65582 64212
rect 353386 64200 353392 64212
rect 353444 64200 353450 64252
rect 61378 64132 61384 64184
rect 61436 64172 61442 64184
rect 351914 64172 351920 64184
rect 61436 64144 351920 64172
rect 61436 64132 61442 64144
rect 351914 64132 351920 64144
rect 351972 64132 351978 64184
rect 209314 63520 209320 63572
rect 209372 63560 209378 63572
rect 300026 63560 300032 63572
rect 209372 63532 300032 63560
rect 209372 63520 209378 63532
rect 300026 63520 300032 63532
rect 300084 63520 300090 63572
rect 156598 63452 156604 63504
rect 156656 63492 156662 63504
rect 197814 63492 197820 63504
rect 156656 63464 197820 63492
rect 156656 63452 156662 63464
rect 197814 63452 197820 63464
rect 197872 63452 197878 63504
rect 336826 63452 336832 63504
rect 336884 63492 336890 63504
rect 364334 63492 364340 63504
rect 336884 63464 364340 63492
rect 336884 63452 336890 63464
rect 364334 63452 364340 63464
rect 364392 63452 364398 63504
rect 99374 62976 99380 63028
rect 99432 63016 99438 63028
rect 222562 63016 222568 63028
rect 99432 62988 222568 63016
rect 99432 62976 99438 62988
rect 222562 62976 222568 62988
rect 222620 62976 222626 63028
rect 320266 62976 320272 63028
rect 320324 63016 320330 63028
rect 329926 63016 329932 63028
rect 320324 62988 329932 63016
rect 320324 62976 320330 62988
rect 329926 62976 329932 62988
rect 329984 62976 329990 63028
rect 219434 62908 219440 62960
rect 219492 62948 219498 62960
rect 411898 62948 411904 62960
rect 219492 62920 411904 62948
rect 219492 62908 219498 62920
rect 411898 62908 411904 62920
rect 411956 62908 411962 62960
rect 42058 62840 42064 62892
rect 42116 62880 42122 62892
rect 343634 62880 343640 62892
rect 42116 62852 343640 62880
rect 42116 62840 42122 62852
rect 343634 62840 343640 62852
rect 343692 62840 343698 62892
rect 35158 62772 35164 62824
rect 35216 62812 35222 62824
rect 340138 62812 340144 62824
rect 35216 62784 340144 62812
rect 35216 62772 35222 62784
rect 340138 62772 340144 62784
rect 340196 62772 340202 62824
rect 341058 62772 341064 62824
rect 341116 62812 341122 62824
rect 433978 62812 433984 62824
rect 341116 62784 433984 62812
rect 341116 62772 341122 62784
rect 433978 62772 433984 62784
rect 434036 62772 434042 62824
rect 197814 62092 197820 62144
rect 197872 62132 197878 62144
rect 283834 62132 283840 62144
rect 197872 62104 283840 62132
rect 197872 62092 197878 62104
rect 283834 62092 283840 62104
rect 283892 62092 283898 62144
rect 335354 62092 335360 62144
rect 335412 62132 335418 62144
rect 336826 62132 336832 62144
rect 335412 62104 336832 62132
rect 335412 62092 335418 62104
rect 336826 62092 336832 62104
rect 336884 62092 336890 62144
rect 5166 62024 5172 62076
rect 5224 62064 5230 62076
rect 57054 62064 57060 62076
rect 5224 62036 57060 62064
rect 5224 62024 5230 62036
rect 57054 62024 57060 62036
rect 57112 62024 57118 62076
rect 298002 62024 298008 62076
rect 298060 62064 298066 62076
rect 383654 62064 383660 62076
rect 298060 62036 383660 62064
rect 298060 62024 298066 62036
rect 383654 62024 383660 62036
rect 383712 62024 383718 62076
rect 207658 61548 207664 61600
rect 207716 61588 207722 61600
rect 298002 61588 298008 61600
rect 207716 61560 298008 61588
rect 207716 61548 207722 61560
rect 298002 61548 298008 61560
rect 298060 61548 298066 61600
rect 211154 61480 211160 61532
rect 211212 61520 211218 61532
rect 392578 61520 392584 61532
rect 211212 61492 392584 61520
rect 211212 61480 211218 61492
rect 392578 61480 392584 61492
rect 392636 61480 392642 61532
rect 214282 61412 214288 61464
rect 214340 61452 214346 61464
rect 399478 61452 399484 61464
rect 214340 61424 399484 61452
rect 214340 61412 214346 61424
rect 399478 61412 399484 61424
rect 399536 61412 399542 61464
rect 217594 61344 217600 61396
rect 217652 61384 217658 61396
rect 407758 61384 407764 61396
rect 217652 61356 407764 61384
rect 217652 61344 217658 61356
rect 407758 61344 407764 61356
rect 407816 61344 407822 61396
rect 114554 60664 114560 60716
rect 114612 60704 114618 60716
rect 202966 60704 202972 60716
rect 114612 60676 202972 60704
rect 114612 60664 114618 60676
rect 202966 60664 202972 60676
rect 203024 60704 203030 60716
rect 204070 60704 204076 60716
rect 203024 60676 204076 60704
rect 203024 60664 203030 60676
rect 204070 60664 204076 60676
rect 204128 60664 204134 60716
rect 295334 60664 295340 60716
rect 295392 60704 295398 60716
rect 296622 60704 296628 60716
rect 295392 60676 296628 60704
rect 295392 60664 295398 60676
rect 296622 60664 296628 60676
rect 296680 60704 296686 60716
rect 379514 60704 379520 60716
rect 296680 60676 379520 60704
rect 296680 60664 296686 60676
rect 379514 60664 379520 60676
rect 379572 60664 379578 60716
rect 122834 60596 122840 60648
rect 122892 60636 122898 60648
rect 202874 60636 202880 60648
rect 122892 60608 202880 60636
rect 122892 60596 122898 60608
rect 202874 60596 202880 60608
rect 202932 60636 202938 60648
rect 204162 60636 204168 60648
rect 202932 60608 204168 60636
rect 202932 60596 202938 60608
rect 204162 60596 204168 60608
rect 204220 60596 204226 60648
rect 206002 60188 206008 60240
rect 206060 60228 206066 60240
rect 295334 60228 295340 60240
rect 206060 60200 295340 60228
rect 206060 60188 206066 60200
rect 295334 60188 295340 60200
rect 295392 60188 295398 60240
rect 204162 60120 204168 60172
rect 204220 60160 204226 60172
rect 232498 60160 232504 60172
rect 204220 60132 232504 60160
rect 204220 60120 204226 60132
rect 232498 60120 232504 60132
rect 232556 60120 232562 60172
rect 249058 60120 249064 60172
rect 249116 60160 249122 60172
rect 283558 60160 283564 60172
rect 249116 60132 283564 60160
rect 249116 60120 249122 60132
rect 283558 60120 283564 60132
rect 283616 60120 283622 60172
rect 283650 60120 283656 60172
rect 283708 60160 283714 60172
rect 386506 60160 386512 60172
rect 283708 60132 386512 60160
rect 283708 60120 283714 60132
rect 386506 60120 386512 60132
rect 386564 60120 386570 60172
rect 204070 60052 204076 60104
rect 204128 60092 204134 60104
rect 229186 60092 229192 60104
rect 204128 60064 229192 60092
rect 204128 60052 204134 60064
rect 229186 60052 229192 60064
rect 229244 60052 229250 60104
rect 229738 60052 229744 60104
rect 229796 60092 229802 60104
rect 364978 60092 364984 60104
rect 229796 60064 364984 60092
rect 229796 60052 229802 60064
rect 364978 60052 364984 60064
rect 365036 60052 365042 60104
rect 379882 60052 379888 60104
rect 379940 60092 379946 60104
rect 469214 60092 469220 60104
rect 379940 60064 469220 60092
rect 379940 60052 379946 60064
rect 469214 60052 469220 60064
rect 469272 60052 469278 60104
rect 191834 59984 191840 60036
rect 191892 60024 191898 60036
rect 204346 60024 204352 60036
rect 191892 59996 204352 60024
rect 191892 59984 191898 59996
rect 204346 59984 204352 59996
rect 204404 59984 204410 60036
rect 215938 59984 215944 60036
rect 215996 60024 216002 60036
rect 403618 60024 403624 60036
rect 215996 59996 403624 60024
rect 215996 59984 216002 59996
rect 403618 59984 403624 59996
rect 403676 59984 403682 60036
rect 180794 59304 180800 59356
rect 180852 59344 180858 59356
rect 200482 59344 200488 59356
rect 180852 59316 200488 59344
rect 180852 59304 180858 59316
rect 200482 59304 200488 59316
rect 200540 59344 200546 59356
rect 201402 59344 201408 59356
rect 200540 59316 201408 59344
rect 200540 59304 200546 59316
rect 201402 59304 201408 59316
rect 201460 59304 201466 59356
rect 323578 58964 323584 59016
rect 323636 59004 323642 59016
rect 336734 59004 336740 59016
rect 323636 58976 336740 59004
rect 323636 58964 323642 58976
rect 336734 58964 336740 58976
rect 336792 58964 336798 59016
rect 296530 58828 296536 58880
rect 296588 58868 296594 58880
rect 336826 58868 336832 58880
rect 296588 58840 336832 58868
rect 296588 58828 296594 58840
rect 336826 58828 336832 58840
rect 336884 58868 336890 58880
rect 336884 58840 345014 58868
rect 336884 58828 336890 58840
rect 201402 58760 201408 58812
rect 201460 58800 201466 58812
rect 308674 58800 308680 58812
rect 201460 58772 308680 58800
rect 201460 58760 201466 58772
rect 308674 58760 308680 58772
rect 308732 58760 308738 58812
rect 325234 58760 325240 58812
rect 325292 58800 325298 58812
rect 340966 58800 340972 58812
rect 325292 58772 340972 58800
rect 325292 58760 325298 58772
rect 340966 58760 340972 58772
rect 341024 58760 341030 58812
rect 184934 58692 184940 58744
rect 184992 58732 184998 58744
rect 310606 58732 310612 58744
rect 184992 58704 310612 58732
rect 184992 58692 184998 58704
rect 310606 58692 310612 58704
rect 310664 58692 310670 58744
rect 344986 58732 345014 58840
rect 368474 58732 368480 58744
rect 344986 58704 368480 58732
rect 368474 58692 368480 58704
rect 368532 58692 368538 58744
rect 195974 58624 195980 58676
rect 196032 58664 196038 58676
rect 381538 58664 381544 58676
rect 196032 58636 381544 58664
rect 196032 58624 196038 58636
rect 381538 58624 381544 58636
rect 381596 58624 381602 58676
rect 396442 58624 396448 58676
rect 396500 58664 396506 58676
rect 476114 58664 476120 58676
rect 396500 58636 476120 58664
rect 396500 58624 396506 58636
rect 476114 58624 476120 58636
rect 476172 58624 476178 58676
rect 153194 57876 153200 57928
rect 153252 57916 153258 57928
rect 200114 57916 200120 57928
rect 153252 57888 200120 57916
rect 153252 57876 153258 57888
rect 200114 57876 200120 57888
rect 200172 57916 200178 57928
rect 201402 57916 201408 57928
rect 200172 57888 201408 57916
rect 200172 57876 200178 57888
rect 201402 57876 201408 57888
rect 201460 57876 201466 57928
rect 258718 57876 258724 57928
rect 258776 57916 258782 57928
rect 262674 57916 262680 57928
rect 258776 57888 262680 57916
rect 258776 57876 258782 57888
rect 262674 57876 262680 57888
rect 262732 57876 262738 57928
rect 310514 57876 310520 57928
rect 310572 57916 310578 57928
rect 312354 57916 312360 57928
rect 310572 57888 312360 57916
rect 310572 57876 310578 57888
rect 312354 57876 312360 57888
rect 312412 57876 312418 57928
rect 161474 57808 161480 57860
rect 161532 57848 161538 57860
rect 201494 57848 201500 57860
rect 161532 57820 201500 57848
rect 161532 57808 161538 57820
rect 201494 57808 201500 57820
rect 201552 57848 201558 57860
rect 202782 57848 202788 57860
rect 201552 57820 202788 57848
rect 201552 57808 201558 57820
rect 202782 57808 202788 57820
rect 202840 57808 202846 57860
rect 274266 57604 274272 57656
rect 274324 57644 274330 57656
rect 311158 57644 311164 57656
rect 274324 57616 311164 57644
rect 274324 57604 274330 57616
rect 311158 57604 311164 57616
rect 311216 57604 311222 57656
rect 332594 57604 332600 57656
rect 332652 57644 332658 57656
rect 350442 57644 350448 57656
rect 332652 57616 350448 57644
rect 332652 57604 332658 57616
rect 350442 57604 350448 57616
rect 350500 57604 350506 57656
rect 277578 57536 277584 57588
rect 277636 57576 277642 57588
rect 341058 57576 341064 57588
rect 277636 57548 341064 57576
rect 277636 57536 277642 57548
rect 341058 57536 341064 57548
rect 341116 57536 341122 57588
rect 300118 57468 300124 57520
rect 300176 57508 300182 57520
rect 367002 57508 367008 57520
rect 300176 57480 367008 57508
rect 300176 57468 300182 57480
rect 367002 57468 367008 57480
rect 367060 57468 367066 57520
rect 300210 57400 300216 57452
rect 300268 57440 300274 57452
rect 383562 57440 383568 57452
rect 300268 57412 383568 57440
rect 300268 57400 300274 57412
rect 383562 57400 383568 57412
rect 383620 57400 383626 57452
rect 201402 57332 201408 57384
rect 201460 57372 201466 57384
rect 287514 57372 287520 57384
rect 201460 57344 287520 57372
rect 201460 57332 201466 57344
rect 287514 57332 287520 57344
rect 287572 57332 287578 57384
rect 298830 57332 298836 57384
rect 298888 57372 298894 57384
rect 385218 57372 385224 57384
rect 298888 57344 385224 57372
rect 298888 57332 298894 57344
rect 385218 57332 385224 57344
rect 385276 57332 385282 57384
rect 280890 57264 280896 57316
rect 280948 57304 280954 57316
rect 442258 57304 442264 57316
rect 280948 57276 442264 57304
rect 280948 57264 280954 57276
rect 442258 57264 442264 57276
rect 442316 57264 442322 57316
rect 202782 57196 202788 57248
rect 202840 57236 202846 57248
rect 290826 57236 290832 57248
rect 202840 57208 290832 57236
rect 202840 57196 202846 57208
rect 290826 57196 290832 57208
rect 290884 57196 290890 57248
rect 300762 57196 300768 57248
rect 300820 57236 300826 57248
rect 465718 57236 465724 57248
rect 300820 57208 465724 57236
rect 300820 57196 300826 57208
rect 465718 57196 465724 57208
rect 465776 57196 465782 57248
rect 315666 56584 315672 56636
rect 315724 56624 315730 56636
rect 317414 56624 317420 56636
rect 315724 56596 317420 56624
rect 315724 56584 315730 56596
rect 317414 56584 317420 56596
rect 317472 56584 317478 56636
rect 8938 56516 8944 56568
rect 8996 56556 9002 56568
rect 57514 56556 57520 56568
rect 8996 56528 57520 56556
rect 8996 56516 9002 56528
rect 57514 56516 57520 56528
rect 57572 56516 57578 56568
rect 102134 52640 102140 52692
rect 102192 52680 102198 52692
rect 104066 52680 104072 52692
rect 102192 52652 104072 52680
rect 102192 52640 102198 52652
rect 104066 52640 104072 52652
rect 104124 52640 104130 52692
rect 102134 52504 102140 52556
rect 102192 52544 102198 52556
rect 196158 52544 196164 52556
rect 102192 52516 196164 52544
rect 102192 52504 102198 52516
rect 196158 52504 196164 52516
rect 196216 52504 196222 52556
rect 17218 52368 17224 52420
rect 17276 52408 17282 52420
rect 57054 52408 57060 52420
rect 17276 52380 57060 52408
rect 17276 52368 17282 52380
rect 57054 52368 57060 52380
rect 57112 52368 57118 52420
rect 103054 52368 103060 52420
rect 103112 52408 103118 52420
rect 195974 52408 195980 52420
rect 103112 52380 195980 52408
rect 103112 52368 103118 52380
rect 195974 52368 195980 52380
rect 196032 52368 196038 52420
rect 102778 51008 102784 51060
rect 102836 51048 102842 51060
rect 195974 51048 195980 51060
rect 102836 51020 195980 51048
rect 102836 51008 102842 51020
rect 195974 51008 195980 51020
rect 196032 51008 196038 51060
rect 102594 49648 102600 49700
rect 102652 49688 102658 49700
rect 195974 49688 195980 49700
rect 102652 49660 195980 49688
rect 102652 49648 102658 49660
rect 195974 49648 195980 49660
rect 196032 49648 196038 49700
rect 102962 48220 102968 48272
rect 103020 48260 103026 48272
rect 195974 48260 195980 48272
rect 103020 48232 195980 48260
rect 103020 48220 103026 48232
rect 195974 48220 195980 48232
rect 196032 48220 196038 48272
rect 102226 48152 102232 48204
rect 102284 48192 102290 48204
rect 196066 48192 196072 48204
rect 102284 48164 196072 48192
rect 102284 48152 102290 48164
rect 196066 48152 196072 48164
rect 196124 48152 196130 48204
rect 3602 46860 3608 46912
rect 3660 46900 3666 46912
rect 57514 46900 57520 46912
rect 3660 46872 57520 46900
rect 3660 46860 3666 46872
rect 57514 46860 57520 46872
rect 57572 46860 57578 46912
rect 104066 46860 104072 46912
rect 104124 46900 104130 46912
rect 195974 46900 195980 46912
rect 104124 46872 195980 46900
rect 104124 46860 104130 46872
rect 195974 46860 195980 46872
rect 196032 46860 196038 46912
rect 103238 45500 103244 45552
rect 103296 45540 103302 45552
rect 195974 45540 195980 45552
rect 103296 45512 195980 45540
rect 103296 45500 103302 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 103054 44072 103060 44124
rect 103112 44112 103118 44124
rect 195974 44112 195980 44124
rect 103112 44084 195980 44112
rect 103112 44072 103118 44084
rect 195974 44072 195980 44084
rect 196032 44072 196038 44124
rect 103422 44004 103428 44056
rect 103480 44044 103486 44056
rect 196066 44044 196072 44056
rect 103480 44016 196072 44044
rect 103480 44004 103486 44016
rect 196066 44004 196072 44016
rect 196124 44004 196130 44056
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 57146 42752 57152 42764
rect 4948 42724 57152 42752
rect 4948 42712 4954 42724
rect 57146 42712 57152 42724
rect 57204 42712 57210 42764
rect 102686 42712 102692 42764
rect 102744 42752 102750 42764
rect 195974 42752 195980 42764
rect 102744 42724 195980 42752
rect 102744 42712 102750 42724
rect 195974 42712 195980 42724
rect 196032 42712 196038 42764
rect 102778 41352 102784 41404
rect 102836 41392 102842 41404
rect 195974 41392 195980 41404
rect 102836 41364 195980 41392
rect 102836 41352 102842 41364
rect 195974 41352 195980 41364
rect 196032 41352 196038 41404
rect 102502 39992 102508 40044
rect 102560 40032 102566 40044
rect 195974 40032 195980 40044
rect 102560 40004 195980 40032
rect 102560 39992 102566 40004
rect 195974 39992 195980 40004
rect 196032 39992 196038 40044
rect 102318 39924 102324 39976
rect 102376 39964 102382 39976
rect 196066 39964 196072 39976
rect 102376 39936 196072 39964
rect 102376 39924 102382 39936
rect 196066 39924 196072 39936
rect 196124 39924 196130 39976
rect 102134 38564 102140 38616
rect 102192 38604 102198 38616
rect 196066 38604 196072 38616
rect 102192 38576 196072 38604
rect 102192 38564 102198 38576
rect 196066 38564 196072 38576
rect 196124 38564 196130 38616
rect 102410 38496 102416 38548
rect 102468 38536 102474 38548
rect 195974 38536 195980 38548
rect 102468 38508 195980 38536
rect 102468 38496 102474 38508
rect 195974 38496 195980 38508
rect 196032 38496 196038 38548
rect 3694 37204 3700 37256
rect 3752 37244 3758 37256
rect 57054 37244 57060 37256
rect 3752 37216 57060 37244
rect 3752 37204 3758 37216
rect 57054 37204 57060 37216
rect 57112 37204 57118 37256
rect 102226 37204 102232 37256
rect 102284 37244 102290 37256
rect 195974 37244 195980 37256
rect 102284 37216 195980 37244
rect 102284 37204 102290 37216
rect 195974 37204 195980 37216
rect 196032 37204 196038 37256
rect 102870 35844 102876 35896
rect 102928 35884 102934 35896
rect 195974 35884 195980 35896
rect 102928 35856 195980 35884
rect 102928 35844 102934 35856
rect 195974 35844 195980 35856
rect 196032 35844 196038 35896
rect 102134 35776 102140 35828
rect 102192 35816 102198 35828
rect 196066 35816 196072 35828
rect 102192 35788 196072 35816
rect 102192 35776 102198 35788
rect 196066 35776 196072 35788
rect 196124 35776 196130 35828
rect 102594 34416 102600 34468
rect 102652 34456 102658 34468
rect 195974 34456 195980 34468
rect 102652 34428 195980 34456
rect 102652 34416 102658 34428
rect 195974 34416 195980 34428
rect 196032 34416 196038 34468
rect 102778 34348 102784 34400
rect 102836 34388 102842 34400
rect 196066 34388 196072 34400
rect 102836 34360 196072 34388
rect 102836 34348 102842 34360
rect 196066 34348 196072 34360
rect 196124 34348 196130 34400
rect 102134 33056 102140 33108
rect 102192 33096 102198 33108
rect 195974 33096 195980 33108
rect 102192 33068 195980 33096
rect 102192 33056 102198 33068
rect 195974 33056 195980 33068
rect 196032 33056 196038 33108
rect 3326 31764 3332 31816
rect 3384 31804 3390 31816
rect 59998 31804 60004 31816
rect 3384 31776 60004 31804
rect 3384 31764 3390 31776
rect 59998 31764 60004 31776
rect 60056 31764 60062 31816
rect 5074 31696 5080 31748
rect 5132 31736 5138 31748
rect 57606 31736 57612 31748
rect 5132 31708 57612 31736
rect 5132 31696 5138 31708
rect 57606 31696 57612 31708
rect 57664 31696 57670 31748
rect 102318 31696 102324 31748
rect 102376 31736 102382 31748
rect 195974 31736 195980 31748
rect 102376 31708 195980 31736
rect 102376 31696 102382 31708
rect 195974 31696 195980 31708
rect 196032 31696 196038 31748
rect 102134 31628 102140 31680
rect 102192 31668 102198 31680
rect 196066 31668 196072 31680
rect 102192 31640 196072 31668
rect 102192 31628 102198 31640
rect 196066 31628 196072 31640
rect 196124 31628 196130 31680
rect 102226 30268 102232 30320
rect 102284 30308 102290 30320
rect 195974 30308 195980 30320
rect 102284 30280 195980 30308
rect 102284 30268 102290 30280
rect 195974 30268 195980 30280
rect 196032 30268 196038 30320
rect 102134 30200 102140 30252
rect 102192 30240 102198 30252
rect 196066 30240 196072 30252
rect 102192 30212 196072 30240
rect 102192 30200 102198 30212
rect 196066 30200 196072 30212
rect 196124 30200 196130 30252
rect 102134 28908 102140 28960
rect 102192 28948 102198 28960
rect 195974 28948 195980 28960
rect 102192 28920 195980 28948
rect 102192 28908 102198 28920
rect 195974 28908 195980 28920
rect 196032 28908 196038 28960
rect 102134 28228 102140 28280
rect 102192 28268 102198 28280
rect 195974 28268 195980 28280
rect 102192 28240 195980 28268
rect 102192 28228 102198 28240
rect 195974 28228 195980 28240
rect 196032 28228 196038 28280
rect 21450 27548 21456 27600
rect 21508 27588 21514 27600
rect 57238 27588 57244 27600
rect 21508 27560 57244 27588
rect 21508 27548 21514 27560
rect 57238 27548 57244 27560
rect 57296 27548 57302 27600
rect 102134 27548 102140 27600
rect 102192 27588 102198 27600
rect 195974 27588 195980 27600
rect 102192 27560 195980 27588
rect 102192 27548 102198 27560
rect 195974 27548 195980 27560
rect 196032 27548 196038 27600
rect 102778 26188 102784 26240
rect 102836 26228 102842 26240
rect 195974 26228 195980 26240
rect 102836 26200 195980 26228
rect 102836 26188 102842 26200
rect 195974 26188 195980 26200
rect 196032 26188 196038 26240
rect 59998 24216 60004 24268
rect 60056 24256 60062 24268
rect 335538 24256 335544 24268
rect 60056 24228 335544 24256
rect 60056 24216 60062 24228
rect 335538 24216 335544 24228
rect 335596 24216 335602 24268
rect 3510 24148 3516 24200
rect 3568 24188 3574 24200
rect 364426 24188 364432 24200
rect 3568 24160 364432 24188
rect 3568 24148 3574 24160
rect 364426 24148 364432 24160
rect 364484 24148 364490 24200
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 367830 24120 367836 24132
rect 3476 24092 367836 24120
rect 3476 24080 3482 24092
rect 367830 24080 367836 24092
rect 367888 24080 367894 24132
rect 88978 23468 88984 23520
rect 89036 23508 89042 23520
rect 266354 23508 266360 23520
rect 89036 23480 266360 23508
rect 89036 23468 89042 23480
rect 266354 23468 266360 23480
rect 266412 23508 266418 23520
rect 267366 23508 267372 23520
rect 266412 23480 267372 23508
rect 266412 23468 266418 23480
rect 267366 23468 267372 23480
rect 267424 23468 267430 23520
rect 3602 22720 3608 22772
rect 3660 22760 3666 22772
rect 292574 22760 292580 22772
rect 3660 22732 292580 22760
rect 3660 22720 3666 22732
rect 292574 22720 292580 22732
rect 292632 22720 292638 22772
rect 3786 22108 3792 22160
rect 3844 22148 3850 22160
rect 350166 22148 350172 22160
rect 3844 22120 350172 22148
rect 3844 22108 3850 22120
rect 350166 22108 350172 22120
rect 350224 22108 350230 22160
rect 62298 22040 62304 22092
rect 62356 22080 62362 22092
rect 88978 22080 88984 22092
rect 62356 22052 88984 22080
rect 62356 22040 62362 22052
rect 88978 22040 88984 22052
rect 89036 22040 89042 22092
rect 200022 22040 200028 22092
rect 200080 22080 200086 22092
rect 378870 22080 378876 22092
rect 200080 22052 378876 22080
rect 200080 22040 200086 22052
rect 378870 22040 378876 22052
rect 378928 22040 378934 22092
rect 389634 22040 389640 22092
rect 389692 22080 389698 22092
rect 580258 22080 580264 22092
rect 389692 22052 580264 22080
rect 389692 22040 389698 22052
rect 580258 22040 580264 22052
rect 580316 22040 580322 22092
rect 21358 21972 21364 22024
rect 21416 22012 21422 22024
rect 360930 22012 360936 22024
rect 21416 21984 360936 22012
rect 21416 21972 21422 21984
rect 360930 21972 360936 21984
rect 360988 21972 360994 22024
rect 393222 21972 393228 22024
rect 393280 22012 393286 22024
rect 580350 22012 580356 22024
rect 393280 21984 580356 22012
rect 393280 21972 393286 21984
rect 580350 21972 580356 21984
rect 580408 21972 580414 22024
rect 21634 21904 21640 21956
rect 21692 21944 21698 21956
rect 346578 21944 346584 21956
rect 21692 21916 346584 21944
rect 21692 21904 21698 21916
rect 346578 21904 346584 21916
rect 346636 21904 346642 21956
rect 396810 21904 396816 21956
rect 396868 21944 396874 21956
rect 580442 21944 580448 21956
rect 396868 21916 580448 21944
rect 396868 21904 396874 21916
rect 580442 21904 580448 21916
rect 580500 21904 580506 21956
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 342990 21876 342996 21888
rect 21600 21848 342996 21876
rect 21600 21836 21606 21848
rect 342990 21836 342996 21848
rect 343048 21836 343054 21888
rect 386046 21836 386052 21888
rect 386104 21876 386110 21888
rect 527818 21876 527824 21888
rect 386104 21848 527824 21876
rect 386104 21836 386110 21848
rect 527818 21836 527824 21848
rect 527876 21836 527882 21888
rect 292574 21768 292580 21820
rect 292632 21808 292638 21820
rect 353754 21808 353760 21820
rect 292632 21780 353760 21808
rect 292632 21768 292638 21780
rect 353754 21768 353760 21780
rect 353812 21768 353818 21820
rect 382458 21768 382464 21820
rect 382516 21808 382522 21820
rect 485774 21808 485780 21820
rect 382516 21780 485780 21808
rect 382516 21768 382522 21780
rect 485774 21768 485780 21780
rect 485832 21768 485838 21820
rect 88794 21496 88800 21548
rect 88852 21536 88858 21548
rect 156598 21536 156604 21548
rect 88852 21508 156604 21536
rect 88852 21496 88858 21508
rect 156598 21496 156604 21508
rect 156656 21496 156662 21548
rect 149054 21428 149060 21480
rect 149112 21468 149118 21480
rect 292758 21468 292764 21480
rect 149112 21440 292764 21468
rect 149112 21428 149118 21440
rect 292758 21428 292764 21440
rect 292816 21428 292822 21480
rect 155954 21360 155960 21412
rect 156012 21400 156018 21412
rect 299934 21400 299940 21412
rect 156012 21372 299940 21400
rect 156012 21360 156018 21372
rect 299934 21360 299940 21372
rect 299992 21360 299998 21412
rect 178034 20068 178040 20120
rect 178092 20108 178098 20120
rect 256878 20108 256884 20120
rect 178092 20080 256884 20108
rect 178092 20068 178098 20080
rect 256878 20068 256884 20080
rect 256936 20068 256942 20120
rect 169754 20000 169760 20052
rect 169812 20040 169818 20052
rect 314286 20040 314292 20052
rect 169812 20012 314292 20040
rect 169812 20000 169818 20012
rect 314286 20000 314292 20012
rect 314344 20000 314350 20052
rect 138014 19932 138020 19984
rect 138072 19972 138078 19984
rect 281994 19972 282000 19984
rect 138072 19944 282000 19972
rect 138072 19932 138078 19944
rect 281994 19932 282000 19944
rect 282052 19932 282058 19984
rect 175274 18776 175280 18828
rect 175332 18816 175338 18828
rect 253290 18816 253296 18828
rect 175332 18788 253296 18816
rect 175332 18776 175338 18788
rect 253290 18776 253296 18788
rect 253348 18776 253354 18828
rect 150434 18708 150440 18760
rect 150492 18748 150498 18760
rect 228174 18748 228180 18760
rect 150492 18720 228180 18748
rect 150492 18708 150498 18720
rect 228174 18708 228180 18720
rect 228232 18708 228238 18760
rect 151814 18640 151820 18692
rect 151872 18680 151878 18692
rect 296346 18680 296352 18692
rect 151872 18652 296352 18680
rect 151872 18640 151878 18652
rect 296346 18640 296352 18652
rect 296404 18640 296410 18692
rect 184934 18572 184940 18624
rect 184992 18612 184998 18624
rect 328638 18612 328644 18624
rect 184992 18584 328644 18612
rect 184992 18572 184998 18584
rect 328638 18572 328644 18584
rect 328696 18572 328702 18624
rect 171134 17348 171140 17400
rect 171192 17388 171198 17400
rect 249702 17388 249708 17400
rect 171192 17360 249708 17388
rect 171192 17348 171198 17360
rect 249702 17348 249708 17360
rect 249760 17348 249766 17400
rect 131114 17280 131120 17332
rect 131172 17320 131178 17332
rect 274818 17320 274824 17332
rect 131172 17292 274824 17320
rect 131172 17280 131178 17292
rect 274818 17280 274824 17292
rect 274876 17280 274882 17332
rect 71130 17212 71136 17264
rect 71188 17252 71194 17264
rect 242894 17252 242900 17264
rect 71188 17224 242900 17252
rect 71188 17212 71194 17224
rect 242894 17212 242900 17224
rect 242952 17212 242958 17264
rect 168374 15988 168380 16040
rect 168432 16028 168438 16040
rect 245654 16028 245660 16040
rect 168432 16000 245660 16028
rect 168432 15988 168438 16000
rect 245654 15988 245660 16000
rect 245712 15988 245718 16040
rect 135254 15920 135260 15972
rect 135312 15960 135318 15972
rect 277394 15960 277400 15972
rect 135312 15932 277400 15960
rect 135312 15920 135318 15932
rect 277394 15920 277400 15932
rect 277452 15920 277458 15972
rect 74534 15852 74540 15904
rect 74592 15892 74598 15904
rect 245930 15892 245936 15904
rect 74592 15864 245936 15892
rect 74592 15852 74598 15864
rect 245930 15852 245936 15864
rect 245988 15852 245994 15904
rect 136450 14560 136456 14612
rect 136508 14600 136514 14612
rect 212534 14600 212540 14612
rect 136508 14572 212540 14600
rect 136508 14560 136514 14572
rect 212534 14560 212540 14572
rect 212592 14560 212598 14612
rect 164418 14492 164424 14544
rect 164476 14532 164482 14544
rect 241514 14532 241520 14544
rect 164476 14504 241520 14532
rect 164476 14492 164482 14504
rect 241514 14492 241520 14504
rect 241572 14492 241578 14544
rect 173894 14424 173900 14476
rect 173952 14464 173958 14476
rect 317414 14464 317420 14476
rect 173952 14436 317420 14464
rect 173952 14424 173958 14436
rect 317414 14424 317420 14436
rect 317472 14424 317478 14476
rect 139578 13200 139584 13252
rect 139636 13240 139642 13252
rect 216674 13240 216680 13252
rect 139636 13212 216680 13240
rect 139636 13200 139642 13212
rect 216674 13200 216680 13212
rect 216732 13200 216738 13252
rect 217318 13200 217324 13252
rect 217376 13240 217382 13252
rect 288434 13240 288440 13252
rect 217376 13212 288440 13240
rect 217376 13200 217382 13212
rect 288434 13200 288440 13212
rect 288492 13200 288498 13252
rect 160094 13132 160100 13184
rect 160152 13172 160158 13184
rect 238754 13172 238760 13184
rect 160152 13144 238760 13172
rect 160152 13132 160158 13144
rect 238754 13132 238760 13144
rect 238812 13132 238818 13184
rect 176654 13064 176660 13116
rect 176712 13104 176718 13116
rect 320174 13104 320180 13116
rect 176712 13076 320180 13104
rect 176712 13064 176718 13076
rect 320174 13064 320180 13076
rect 320232 13064 320238 13116
rect 153746 11908 153752 11960
rect 153804 11948 153810 11960
rect 230474 11948 230480 11960
rect 153804 11920 230480 11948
rect 153804 11908 153810 11920
rect 230474 11908 230480 11920
rect 230532 11908 230538 11960
rect 125594 11840 125600 11892
rect 125652 11880 125658 11892
rect 202874 11880 202880 11892
rect 125652 11852 202880 11880
rect 125652 11840 125658 11852
rect 202874 11840 202880 11852
rect 202932 11840 202938 11892
rect 186130 11772 186136 11824
rect 186188 11812 186194 11824
rect 263594 11812 263600 11824
rect 186188 11784 263600 11812
rect 186188 11772 186194 11784
rect 263594 11772 263600 11784
rect 263652 11772 263658 11824
rect 142154 11704 142160 11756
rect 142212 11744 142218 11756
rect 284294 11744 284300 11756
rect 142212 11716 284300 11744
rect 142212 11704 142218 11716
rect 284294 11704 284300 11716
rect 284352 11704 284358 11756
rect 147122 10412 147128 10464
rect 147180 10452 147186 10464
rect 223574 10452 223580 10464
rect 147180 10424 223580 10452
rect 147180 10412 147186 10424
rect 223574 10412 223580 10424
rect 223632 10412 223638 10464
rect 156598 10344 156604 10396
rect 156656 10384 156662 10396
rect 245194 10384 245200 10396
rect 156656 10356 245200 10384
rect 156656 10344 156662 10356
rect 245194 10344 245200 10356
rect 245252 10344 245258 10396
rect 3418 10276 3424 10328
rect 3476 10316 3482 10328
rect 338114 10316 338120 10328
rect 3476 10288 338120 10316
rect 3476 10276 3482 10288
rect 338114 10276 338120 10288
rect 338172 10276 338178 10328
rect 163682 9052 163688 9104
rect 163740 9092 163746 9104
rect 306374 9092 306380 9104
rect 163740 9064 306380 9092
rect 163740 9052 163746 9064
rect 306374 9052 306380 9064
rect 306432 9052 306438 9104
rect 167178 8984 167184 9036
rect 167236 9024 167242 9036
rect 310514 9024 310520 9036
rect 167236 8996 310520 9024
rect 167236 8984 167242 8996
rect 310514 8984 310520 8996
rect 310572 8984 310578 9036
rect 84194 8916 84200 8968
rect 84252 8956 84258 8968
rect 241698 8956 241704 8968
rect 84252 8928 241704 8956
rect 84252 8916 84258 8928
rect 241698 8916 241704 8928
rect 241756 8916 241762 8968
rect 157794 7760 157800 7812
rect 157852 7800 157858 7812
rect 234614 7800 234620 7812
rect 157852 7772 234620 7800
rect 157852 7760 157858 7772
rect 234614 7760 234620 7772
rect 234672 7760 234678 7812
rect 132954 7692 132960 7744
rect 133012 7732 133018 7744
rect 209774 7732 209780 7744
rect 133012 7704 209780 7732
rect 133012 7692 133018 7704
rect 209774 7692 209780 7704
rect 209832 7692 209838 7744
rect 188522 7624 188528 7676
rect 188580 7664 188586 7676
rect 331214 7664 331220 7676
rect 188580 7636 331220 7664
rect 188580 7624 188586 7636
rect 331214 7624 331220 7636
rect 331272 7624 331278 7676
rect 128170 7556 128176 7608
rect 128228 7596 128234 7608
rect 270494 7596 270500 7608
rect 128228 7568 270500 7596
rect 128228 7556 128234 7568
rect 270494 7556 270500 7568
rect 270552 7556 270558 7608
rect 143534 6264 143540 6316
rect 143592 6304 143598 6316
rect 220814 6304 220820 6316
rect 143592 6276 220820 6304
rect 143592 6264 143598 6276
rect 220814 6264 220820 6276
rect 220872 6264 220878 6316
rect 181438 6196 181444 6248
rect 181496 6236 181502 6248
rect 324314 6236 324320 6248
rect 181496 6208 324320 6236
rect 181496 6196 181502 6208
rect 324314 6196 324320 6208
rect 324372 6196 324378 6248
rect 78674 6128 78680 6180
rect 78732 6168 78738 6180
rect 249978 6168 249984 6180
rect 78732 6140 249984 6168
rect 78732 6128 78738 6140
rect 249978 6128 249984 6140
rect 250036 6128 250042 6180
rect 182542 4972 182548 5024
rect 182600 5012 182606 5024
rect 259454 5012 259460 5024
rect 182600 4984 259460 5012
rect 182600 4972 182606 4984
rect 259454 4972 259460 4984
rect 259512 4972 259518 5024
rect 129366 4904 129372 4956
rect 129424 4944 129430 4956
rect 205634 4944 205640 4956
rect 129424 4916 205640 4944
rect 129424 4904 129430 4916
rect 205634 4904 205640 4916
rect 205692 4904 205698 4956
rect 96614 4836 96620 4888
rect 96672 4876 96678 4888
rect 252370 4876 252376 4888
rect 96672 4848 252376 4876
rect 96672 4836 96678 4848
rect 252370 4836 252376 4848
rect 252428 4836 252434 4888
rect 92474 4768 92480 4820
rect 92532 4808 92538 4820
rect 248782 4808 248788 4820
rect 92532 4780 248788 4808
rect 92532 4768 92538 4780
rect 248782 4768 248788 4780
rect 248840 4768 248846 4820
rect 145926 3544 145932 3596
rect 145984 3584 145990 3596
rect 217318 3584 217324 3596
rect 145984 3556 217324 3584
rect 145984 3544 145990 3556
rect 217318 3544 217324 3556
rect 217376 3544 217382 3596
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153010 3516 153016 3528
rect 151872 3488 153016 3516
rect 151872 3476 151878 3488
rect 153010 3476 153016 3488
rect 153068 3476 153074 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 161382 3476 161388 3528
rect 161440 3516 161446 3528
rect 302234 3516 302240 3528
rect 161440 3488 302240 3516
rect 161440 3476 161446 3488
rect 302234 3476 302240 3488
rect 302292 3476 302298 3528
rect 66254 3408 66260 3460
rect 66312 3448 66318 3460
rect 239306 3448 239312 3460
rect 66312 3420 239312 3448
rect 66312 3408 66318 3420
rect 239306 3408 239312 3420
rect 239364 3408 239370 3460
rect 266354 3408 266360 3460
rect 266412 3448 266418 3460
rect 579798 3448 579804 3460
rect 266412 3420 579804 3448
rect 266412 3408 266418 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 177850 3380 177856 3392
rect 176712 3352 177856 3380
rect 176712 3340 176718 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 160094 2796 160100 2848
rect 160152 2836 160158 2848
rect 161382 2836 161388 2848
rect 160152 2808 161388 2836
rect 160152 2796 160158 2808
rect 161382 2796 161388 2808
rect 161440 2796 161446 2848
<< via1 >>
rect 8116 700952 8168 701004
rect 72976 700952 73028 701004
rect 397460 700952 397512 701004
rect 462320 700952 462372 701004
rect 463608 700952 463660 701004
rect 22008 700340 22060 700392
rect 89168 700340 89220 700392
rect 137836 700340 137888 700392
rect 198740 700340 198792 700392
rect 22192 700272 22244 700324
rect 154120 700272 154172 700324
rect 302240 700272 302292 700324
rect 413652 700272 413704 700324
rect 463608 700272 463660 700324
rect 485780 700272 485832 700324
rect 198740 699796 198792 699848
rect 200028 699796 200080 699848
rect 202788 699796 202840 699848
rect 22100 699660 22152 699712
rect 24308 699660 24360 699712
rect 527180 697552 527232 697604
rect 527824 697552 527876 697604
rect 580172 697552 580224 697604
rect 3424 671168 3476 671220
rect 8944 671168 8996 671220
rect 92940 586440 92992 586492
rect 96160 586440 96212 586492
rect 373264 586440 373316 586492
rect 376484 586440 376536 586492
rect 21824 586168 21876 586220
rect 34520 586168 34572 586220
rect 193128 586168 193180 586220
rect 200212 586168 200264 586220
rect 301780 586168 301832 586220
rect 310796 586168 310848 586220
rect 21640 586100 21692 586152
rect 42064 586100 42116 586152
rect 185676 586100 185728 586152
rect 200304 586100 200356 586152
rect 301872 586100 301924 586152
rect 314660 586100 314712 586152
rect 372620 586100 372672 586152
rect 373264 586100 373316 586152
rect 465356 586100 465408 586152
rect 479064 586100 479116 586152
rect 22928 586032 22980 586084
rect 45928 586032 45980 586084
rect 181812 586032 181864 586084
rect 198096 586032 198148 586084
rect 302700 586032 302752 586084
rect 318524 586032 318576 586084
rect 461492 586032 461544 586084
rect 478144 586032 478196 586084
rect 20536 585964 20588 586016
rect 49792 585964 49844 586016
rect 177948 585964 178000 586016
rect 198924 585964 198976 586016
rect 302148 585964 302200 586016
rect 322388 585964 322440 586016
rect 457628 585964 457680 586016
rect 478972 585964 479024 586016
rect 21732 585896 21784 585948
rect 53840 585896 53892 585948
rect 173808 585896 173860 585948
rect 198004 585896 198056 585948
rect 302884 585896 302936 585948
rect 326252 585896 326304 585948
rect 453764 585896 453816 585948
rect 477960 585896 478012 585948
rect 21916 585828 21968 585880
rect 30472 585828 30524 585880
rect 32404 585828 32456 585880
rect 65248 585828 65300 585880
rect 170220 585828 170272 585880
rect 198740 585828 198792 585880
rect 301964 585828 302016 585880
rect 330116 585828 330168 585880
rect 449900 585828 449952 585880
rect 479156 585828 479208 585880
rect 22836 585760 22888 585812
rect 38200 585760 38252 585812
rect 39304 585760 39356 585812
rect 88432 585760 88484 585812
rect 166356 585760 166408 585812
rect 197912 585760 197964 585812
rect 302792 585760 302844 585812
rect 333980 585760 334032 585812
rect 446036 585760 446088 585812
rect 477868 585760 477920 585812
rect 473084 585148 473136 585200
rect 478052 585148 478104 585200
rect 300676 583380 300728 583432
rect 341708 583380 341760 583432
rect 442172 583380 442224 583432
rect 481640 583380 481692 583432
rect 158628 583312 158680 583364
rect 201592 583312 201644 583364
rect 299296 583312 299348 583364
rect 353300 583312 353352 583364
rect 426716 583312 426768 583364
rect 481824 583312 481876 583364
rect 150900 583244 150952 583296
rect 198832 583244 198884 583296
rect 300768 583244 300820 583296
rect 357164 583244 357216 583296
rect 422852 583244 422904 583296
rect 480720 583244 480772 583296
rect 147036 583176 147088 583228
rect 201500 583176 201552 583228
rect 300584 583176 300636 583228
rect 361028 583176 361080 583228
rect 415124 583176 415176 583228
rect 478880 583176 478932 583228
rect 143172 583108 143224 583160
rect 200396 583108 200448 583160
rect 300492 583108 300544 583160
rect 364892 583108 364944 583160
rect 411260 583108 411312 583160
rect 484400 583108 484452 583160
rect 127716 583040 127768 583092
rect 200120 583040 200172 583092
rect 297824 583040 297876 583092
rect 368756 583040 368808 583092
rect 407396 583040 407448 583092
rect 483020 583040 483072 583092
rect 20628 582972 20680 583024
rect 73160 582972 73212 583024
rect 123852 582972 123904 583024
rect 199384 582972 199436 583024
rect 298008 582972 298060 583024
rect 380348 582972 380400 583024
rect 403532 582972 403584 583024
rect 480260 582972 480312 583024
rect 297916 580320 297968 580372
rect 384212 580320 384264 580372
rect 399668 580320 399720 580372
rect 483112 580320 483164 580372
rect 299388 580252 299440 580304
rect 388076 580252 388128 580304
rect 395804 580252 395856 580304
rect 483204 580252 483256 580304
rect 577504 577260 577556 577312
rect 579620 577260 579672 577312
rect 19156 572364 19208 572416
rect 32404 572364 32456 572416
rect 161480 572364 161532 572416
rect 201776 572364 201828 572416
rect 18880 572296 18932 572348
rect 39304 572296 39356 572348
rect 153200 572296 153252 572348
rect 201684 572296 201736 572348
rect 19064 572228 19116 572280
rect 75920 572228 75972 572280
rect 131120 572228 131172 572280
rect 202972 572228 203024 572280
rect 20352 572160 20404 572212
rect 80060 572160 80112 572212
rect 118700 572160 118752 572212
rect 202880 572160 202932 572212
rect 19984 572092 20036 572144
rect 99380 572092 99432 572144
rect 114560 572092 114612 572144
rect 203064 572092 203116 572144
rect 18972 572024 19024 572076
rect 103520 572024 103572 572076
rect 189080 572024 189132 572076
rect 298744 572024 298796 572076
rect 300400 572024 300452 572076
rect 345020 572024 345072 572076
rect 437480 572024 437532 572076
rect 480536 572024 480588 572076
rect 20444 571956 20496 572008
rect 107660 571956 107712 572008
rect 138020 571956 138072 572008
rect 245660 571956 245712 572008
rect 247040 571956 247092 572008
rect 418160 571956 418212 572008
rect 433340 571956 433392 572008
rect 481732 571956 481784 572008
rect 263600 570596 263652 570648
rect 373264 570596 373316 570648
rect 2780 565904 2832 565956
rect 4896 565904 4948 565956
rect 3424 514768 3476 514820
rect 7564 514768 7616 514820
rect 480904 470568 480956 470620
rect 580172 470568 580224 470620
rect 20260 465740 20312 465792
rect 20536 465740 20588 465792
rect 478788 462884 478840 462936
rect 480444 462884 480496 462936
rect 22100 462612 22152 462664
rect 23204 462612 23256 462664
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 199016 462340 199068 462392
rect 199384 462340 199436 462392
rect 204260 462340 204312 462392
rect 392216 462340 392268 462392
rect 478788 462340 478840 462392
rect 300308 462272 300360 462324
rect 300492 462272 300544 462324
rect 479156 462272 479208 462324
rect 479340 462272 479392 462324
rect 480628 462272 480680 462324
rect 481640 462272 481692 462324
rect 20168 461524 20220 461576
rect 20444 461524 20496 461576
rect 18604 461320 18656 461372
rect 18972 461320 19024 461372
rect 18880 461116 18932 461168
rect 88432 461116 88484 461168
rect 158628 461116 158680 461168
rect 201592 461116 201644 461168
rect 300308 461116 300360 461168
rect 364248 461116 364300 461168
rect 453948 461116 454000 461168
rect 477960 461116 478012 461168
rect 17776 461048 17828 461100
rect 19984 461048 20036 461100
rect 100346 461048 100398 461100
rect 146714 461048 146766 461100
rect 201500 461048 201552 461100
rect 300768 461048 300820 461100
rect 357164 461048 357216 461100
rect 449900 461048 449952 461100
rect 479340 461048 479392 461100
rect 18972 460980 19024 461032
rect 104210 460980 104262 461032
rect 142850 460980 142902 461032
rect 200396 460980 200448 461032
rect 300584 460980 300636 461032
rect 361028 460980 361080 461032
rect 446036 460980 446088 461032
rect 477868 460980 477920 461032
rect 20168 460912 20220 460964
rect 107752 460912 107804 460964
rect 123852 460912 123904 460964
rect 199016 460912 199068 460964
rect 297916 460912 297968 460964
rect 384212 460912 384264 460964
rect 442172 460912 442224 460964
rect 480628 460980 480680 461032
rect 177948 460844 178000 460896
rect 198924 460844 198976 460896
rect 473084 460844 473136 460896
rect 478052 460844 478104 460896
rect 22008 459484 22060 459536
rect 26608 459484 26660 459536
rect 92940 459484 92992 459536
rect 95884 459484 95936 459536
rect 115848 459484 115900 459536
rect 203248 459484 203300 459536
rect 372620 459484 372672 459536
rect 373264 459484 373316 459536
rect 376484 459484 376536 459536
rect 415124 459484 415176 459536
rect 418712 459484 418764 459536
rect 457628 459484 457680 459536
rect 461492 459484 461544 459536
rect 461584 459484 461636 459536
rect 463792 459484 463844 459536
rect 465356 459484 465408 459536
rect 469312 459484 469364 459536
rect 18972 459416 19024 459468
rect 76840 459416 76892 459468
rect 131580 459416 131632 459468
rect 202972 459416 203024 459468
rect 298008 459416 298060 459468
rect 380348 459416 380400 459468
rect 407396 459416 407448 459468
rect 483020 459416 483072 459468
rect 19248 459348 19300 459400
rect 61384 459348 61436 459400
rect 135168 459348 135220 459400
rect 197360 459348 197412 459400
rect 297824 459348 297876 459400
rect 368756 459348 368808 459400
rect 411260 459348 411312 459400
rect 484400 459348 484452 459400
rect 20352 459280 20404 459332
rect 80704 459280 80756 459332
rect 162492 459280 162544 459332
rect 201868 459280 201920 459332
rect 299296 459280 299348 459332
rect 353300 459280 353352 459332
rect 430580 459280 430632 459332
rect 479156 459280 479208 459332
rect 300492 459212 300544 459264
rect 345572 459212 345624 459264
rect 438308 459212 438360 459264
rect 480536 459212 480588 459264
rect 300676 459144 300728 459196
rect 341708 459144 341760 459196
rect 403532 459144 403584 459196
rect 480260 459144 480312 459196
rect 482100 459144 482152 459196
rect 299388 459076 299440 459128
rect 388076 459076 388128 459128
rect 19156 459008 19208 459060
rect 20444 459008 20496 459060
rect 42800 459008 42852 459060
rect 45928 459008 45980 459060
rect 20628 458940 20680 458992
rect 21456 458940 21508 458992
rect 22744 458940 22796 458992
rect 30472 458940 30524 458992
rect 154488 458940 154540 458992
rect 200396 458940 200448 458992
rect 201684 458940 201736 458992
rect 20444 458872 20496 458924
rect 65248 458872 65300 458924
rect 119988 458872 120040 458924
rect 197176 458872 197228 458924
rect 202880 458872 202932 458924
rect 469220 458872 469272 458924
rect 481640 458872 481692 458924
rect 21456 458804 21508 458856
rect 73160 458804 73212 458856
rect 139308 458804 139360 458856
rect 244280 458804 244332 458856
rect 283564 458804 283616 458856
rect 418988 458804 419040 458856
rect 434444 458804 434496 458856
rect 480352 458804 480404 458856
rect 481732 458804 481784 458856
rect 30380 458464 30432 458516
rect 34520 458464 34572 458516
rect 18788 458192 18840 458244
rect 19248 458192 19300 458244
rect 483020 458192 483072 458244
rect 484492 458192 484544 458244
rect 150900 458124 150952 458176
rect 198832 458124 198884 458176
rect 302792 458124 302844 458176
rect 333980 458124 334032 458176
rect 395804 458124 395856 458176
rect 483296 458124 483348 458176
rect 20260 458056 20312 458108
rect 49792 458056 49844 458108
rect 166356 458056 166408 458108
rect 197912 458056 197964 458108
rect 301964 458056 302016 458108
rect 330116 458056 330168 458108
rect 399668 458056 399720 458108
rect 483112 458056 483164 458108
rect 21916 457988 21968 458040
rect 22744 457988 22796 458040
rect 22928 457988 22980 458040
rect 42800 457988 42852 458040
rect 170220 457988 170272 458040
rect 198740 457988 198792 458040
rect 302884 457988 302936 458040
rect 326252 457988 326304 458040
rect 418712 457988 418764 458040
rect 478880 457988 478932 458040
rect 21732 457920 21784 457972
rect 53840 457920 53892 457972
rect 422852 457920 422904 457972
rect 480720 457920 480772 457972
rect 483204 457920 483256 457972
rect 426716 457852 426768 457904
rect 481824 457852 481876 457904
rect 21824 457444 21876 457496
rect 22836 457444 22888 457496
rect 30380 457444 30432 457496
rect 20536 456764 20588 456816
rect 22928 456764 22980 456816
rect 197912 456764 197964 456816
rect 198096 456764 198148 456816
rect 198832 456764 198884 456816
rect 199016 456764 199068 456816
rect 302608 456764 302660 456816
rect 302792 456764 302844 456816
rect 478788 456696 478840 456748
rect 480444 456696 480496 456748
rect 264980 445000 265032 445052
rect 373264 445000 373316 445052
rect 126980 444320 127032 444372
rect 200120 444320 200172 444372
rect 201776 444320 201828 444372
rect 21548 443912 21600 443964
rect 23480 443912 23532 443964
rect 197268 443708 197320 443760
rect 204352 443708 204404 443760
rect 95884 443640 95936 443692
rect 260840 443640 260892 443692
rect 2872 410184 2924 410236
rect 4988 410184 5040 410236
rect 479524 364352 479576 364404
rect 580172 364352 580224 364404
rect 3332 345040 3384 345092
rect 20904 345040 20956 345092
rect 200488 335248 200540 335300
rect 200580 335044 200632 335096
rect 21456 334636 21508 334688
rect 72976 334636 73028 334688
rect 18604 334568 18656 334620
rect 103888 334568 103940 334620
rect 17960 334092 18012 334144
rect 18604 334092 18656 334144
rect 19248 334024 19300 334076
rect 19156 333956 19208 334008
rect 21456 333956 21508 334008
rect 76840 333956 76892 334008
rect 442448 333956 442500 334008
rect 480628 333956 480680 334008
rect 478420 333276 478472 333328
rect 479156 333276 479208 333328
rect 438860 333208 438912 333260
rect 480536 333208 480588 333260
rect 482008 333208 482060 333260
rect 162492 332936 162544 332988
rect 201684 332936 201736 332988
rect 201868 332936 201920 332988
rect 158720 332868 158772 332920
rect 201592 332868 201644 332920
rect 201960 332868 202012 332920
rect 299296 332868 299348 332920
rect 300124 332868 300176 332920
rect 350540 332868 350592 332920
rect 8944 332800 8996 332852
rect 26608 332800 26660 332852
rect 154764 332800 154816 332852
rect 200304 332800 200356 332852
rect 302884 332800 302936 332852
rect 361580 332800 361632 332852
rect 20352 332732 20404 332784
rect 80704 332732 80756 332784
rect 137928 332732 137980 332784
rect 197360 332732 197412 332784
rect 297732 332732 297784 332784
rect 368756 332732 368808 332784
rect 433248 332732 433300 332784
rect 478420 332732 478472 332784
rect 16488 332664 16540 332716
rect 17776 332664 17828 332716
rect 100024 332664 100076 332716
rect 143172 332664 143224 332716
rect 200396 332664 200448 332716
rect 202052 332664 202104 332716
rect 297916 332664 297968 332716
rect 384212 332664 384264 332716
rect 395804 332664 395856 332716
rect 483204 332664 483256 332716
rect 20076 332596 20128 332648
rect 107752 332596 107804 332648
rect 123852 332596 123904 332648
rect 199936 332596 199988 332648
rect 3608 332528 3660 332580
rect 22928 332528 22980 332580
rect 92940 332528 92992 332580
rect 96436 332528 96488 332580
rect 135076 332528 135128 332580
rect 137928 332528 137980 332580
rect 166356 332528 166408 332580
rect 198096 332528 198148 332580
rect 306932 332596 306984 332648
rect 577504 332596 577556 332648
rect 204260 332528 204312 332580
rect 300492 332528 300544 332580
rect 345572 332528 345624 332580
rect 350540 332528 350592 332580
rect 353300 332528 353352 332580
rect 361580 332528 361632 332580
rect 364892 332528 364944 332580
rect 372620 332528 372672 332580
rect 376484 332528 376536 332580
rect 430580 332528 430632 332580
rect 433248 332528 433300 332580
rect 473084 332528 473136 332580
rect 478052 332528 478104 332580
rect 20168 332460 20220 332512
rect 49792 332460 49844 332512
rect 170220 332460 170272 332512
rect 198832 332460 198884 332512
rect 301964 332460 302016 332512
rect 330116 332460 330168 332512
rect 449900 332460 449952 332512
rect 479340 332460 479392 332512
rect 20536 332392 20588 332444
rect 45928 332392 45980 332444
rect 173716 332392 173768 332444
rect 198004 332392 198056 332444
rect 302792 332392 302844 332444
rect 326252 332392 326304 332444
rect 453764 332392 453816 332444
rect 477960 332392 478012 332444
rect 481916 332392 481968 332444
rect 22560 332324 22612 332376
rect 38200 332324 38252 332376
rect 177948 332324 178000 332376
rect 198924 332324 198976 332376
rect 301872 332324 301924 332376
rect 322388 332324 322440 332376
rect 457628 332324 457680 332376
rect 478972 332324 479024 332376
rect 22836 332256 22888 332308
rect 34520 332256 34572 332308
rect 181812 332256 181864 332308
rect 198188 332256 198240 332308
rect 302700 332256 302752 332308
rect 318524 332256 318576 332308
rect 461492 332256 461544 332308
rect 478144 332256 478196 332308
rect 22652 332188 22704 332240
rect 30472 332188 30524 332240
rect 185676 332188 185728 332240
rect 200212 332188 200264 332240
rect 200672 332188 200724 332240
rect 301504 332188 301556 332240
rect 314660 332188 314712 332240
rect 465356 332188 465408 332240
rect 479064 332188 479116 332240
rect 21916 332120 21968 332172
rect 53840 332120 53892 332172
rect 193036 332120 193088 332172
rect 200580 332120 200632 332172
rect 302056 332120 302108 332172
rect 310796 332120 310848 332172
rect 446036 332120 446088 332172
rect 477868 332120 477920 332172
rect 22192 331848 22244 331900
rect 42064 331848 42116 331900
rect 301688 331780 301740 331832
rect 302056 331780 302108 331832
rect 22008 331440 22060 331492
rect 22560 331440 22612 331492
rect 17776 331236 17828 331288
rect 21548 331236 21600 331288
rect 22652 331236 22704 331288
rect 22928 331236 22980 331288
rect 84568 331236 84620 331288
rect 197912 331236 197964 331288
rect 198096 331236 198148 331288
rect 301504 331236 301556 331288
rect 301780 331236 301832 331288
rect 399668 331236 399720 331288
rect 400864 331236 400916 331288
rect 403532 331236 403584 331288
rect 405004 331236 405056 331288
rect 415124 331236 415176 331288
rect 127716 331168 127768 331220
rect 477868 331236 477920 331288
rect 478328 331236 478380 331288
rect 478880 331236 478932 331288
rect 479064 331236 479116 331288
rect 418620 331168 418672 331220
rect 201868 331100 201920 331152
rect 18880 331032 18932 331084
rect 88432 331032 88484 331084
rect 21640 330964 21692 331016
rect 22192 330964 22244 331016
rect 147036 330556 147088 330608
rect 200396 330556 200448 330608
rect 201500 330556 201552 330608
rect 119988 330488 120040 330540
rect 203064 330488 203116 330540
rect 204352 330488 204404 330540
rect 18788 329740 18840 329792
rect 18972 329740 19024 329792
rect 20260 329740 20312 329792
rect 20444 329740 20496 329792
rect 65248 329740 65300 329792
rect 131028 329740 131080 329792
rect 202972 329740 203024 329792
rect 203156 329740 203208 329792
rect 407396 329740 407448 329792
rect 484492 329740 484544 329792
rect 61384 329672 61436 329724
rect 411260 329672 411312 329724
rect 484400 329672 484452 329724
rect 418620 329604 418672 329656
rect 477500 329604 477552 329656
rect 484400 329400 484452 329452
rect 484584 329400 484636 329452
rect 3608 318792 3660 318844
rect 21456 318792 21508 318844
rect 249800 318044 249852 318096
rect 418160 318044 418212 318096
rect 138020 316684 138072 316736
rect 241520 316684 241572 316736
rect 114560 315936 114612 315988
rect 203248 315936 203300 315988
rect 298008 315936 298060 315988
rect 379520 315936 379572 315988
rect 391940 315936 391992 315988
rect 480444 315936 480496 315988
rect 150348 315868 150400 315920
rect 199016 315868 199068 315920
rect 300584 315868 300636 315920
rect 360200 315868 360252 315920
rect 405004 315868 405056 315920
rect 482100 315868 482152 315920
rect 300768 315800 300820 315852
rect 356060 315800 356112 315852
rect 400864 315800 400916 315852
rect 476120 315800 476172 315852
rect 302148 315732 302200 315784
rect 349160 315732 349212 315784
rect 422300 315732 422352 315784
rect 483112 315732 483164 315784
rect 300676 315664 300728 315716
rect 340880 315664 340932 315716
rect 426440 315664 426492 315716
rect 481824 315664 481876 315716
rect 303528 315596 303580 315648
rect 336740 315596 336792 315648
rect 433340 315596 433392 315648
rect 480352 315596 480404 315648
rect 302608 315528 302660 315580
rect 333980 315528 334032 315580
rect 111800 315324 111852 315376
rect 200488 315324 200540 315376
rect 301596 315324 301648 315376
rect 302148 315324 302200 315376
rect 195980 315256 196032 315308
rect 298836 315256 298888 315308
rect 481732 315188 481784 315240
rect 482100 315188 482152 315240
rect 302608 314780 302660 314832
rect 302884 314780 302936 314832
rect 198740 314644 198792 314696
rect 199016 314644 199068 314696
rect 202972 314644 203024 314696
rect 203248 314644 203300 314696
rect 300584 314644 300636 314696
rect 300768 314644 300820 314696
rect 481824 314644 481876 314696
rect 483388 314644 483440 314696
rect 299388 314236 299440 314288
rect 300216 314236 300268 314288
rect 2780 292612 2832 292664
rect 5080 292612 5132 292664
rect 3332 240116 3384 240168
rect 17224 240116 17276 240168
rect 481180 207000 481232 207052
rect 483020 207000 483072 207052
rect 476120 206524 476172 206576
rect 480444 206524 480496 206576
rect 297916 206320 297968 206372
rect 313280 206320 313332 206372
rect 16396 206252 16448 206304
rect 17868 206252 17920 206304
rect 103888 206252 103940 206304
rect 300216 206252 300268 206304
rect 387800 206252 387852 206304
rect 162492 205844 162544 205896
rect 201500 205844 201552 205896
rect 158628 205776 158680 205828
rect 201776 205776 201828 205828
rect 201960 205776 202012 205828
rect 154580 205708 154632 205760
rect 200120 205708 200172 205760
rect 200304 205708 200356 205760
rect 438584 205708 438636 205760
rect 480720 205708 480772 205760
rect 482008 205708 482060 205760
rect 20352 205640 20404 205692
rect 28908 205640 28960 205692
rect 143172 205640 143224 205692
rect 201592 205640 201644 205692
rect 202052 205640 202104 205692
rect 392216 205640 392268 205692
rect 476120 205640 476172 205692
rect 299388 204892 299440 204944
rect 300124 204892 300176 204944
rect 349252 204892 349304 204944
rect 434720 204688 434772 204740
rect 480352 204688 480404 204740
rect 300676 204620 300728 204672
rect 341340 204620 341392 204672
rect 418712 204620 418764 204672
rect 479064 204620 479116 204672
rect 302884 204552 302936 204604
rect 333980 204552 334032 204604
rect 407028 204552 407080 204604
rect 481732 204552 481784 204604
rect 300584 204484 300636 204536
rect 357164 204484 357216 204536
rect 426716 204484 426768 204536
rect 483388 204484 483440 204536
rect 296628 204416 296680 204468
rect 298008 204416 298060 204468
rect 380348 204416 380400 204468
rect 422852 204416 422904 204468
rect 483112 204416 483164 204468
rect 306932 204348 306984 204400
rect 480904 204348 480956 204400
rect 7564 204212 7616 204264
rect 23020 204280 23072 204332
rect 147036 204280 147088 204332
rect 197360 204280 197412 204332
rect 22928 204212 22980 204264
rect 30472 204212 30524 204264
rect 92940 204212 92992 204264
rect 95884 204212 95936 204264
rect 96160 204212 96212 204264
rect 177948 204212 178000 204264
rect 179880 204212 179932 204264
rect 19064 204144 19116 204196
rect 19248 204144 19300 204196
rect 76840 204144 76892 204196
rect 123852 204144 123904 204196
rect 199936 204212 199988 204264
rect 202880 204280 202932 204332
rect 303068 204280 303120 204332
rect 580540 204280 580592 204332
rect 302700 204212 302752 204264
rect 318524 204212 318576 204264
rect 349252 204212 349304 204264
rect 353300 204212 353352 204264
rect 372620 204212 372672 204264
rect 376484 204212 376536 204264
rect 403532 204212 403584 204264
rect 407028 204212 407080 204264
rect 415124 204212 415176 204264
rect 418712 204212 418764 204264
rect 475476 204212 475528 204264
rect 477868 204212 477920 204264
rect 478144 204212 478196 204264
rect 197360 204144 197412 204196
rect 197820 204144 197872 204196
rect 200396 204144 200448 204196
rect 301964 204144 302016 204196
rect 330116 204144 330168 204196
rect 453764 204144 453816 204196
rect 478052 204144 478104 204196
rect 19156 204076 19208 204128
rect 73160 204076 73212 204128
rect 150900 204076 150952 204128
rect 18972 204008 19024 204060
rect 19248 204008 19300 204060
rect 30472 204008 30524 204060
rect 34520 204008 34572 204060
rect 34612 204008 34664 204060
rect 80704 204008 80756 204060
rect 173716 204008 173768 204060
rect 183468 204008 183520 204060
rect 193036 204076 193088 204128
rect 195888 204076 195940 204128
rect 198740 204076 198792 204128
rect 199016 204076 199068 204128
rect 302792 204076 302844 204128
rect 326252 204076 326304 204128
rect 411260 204076 411312 204128
rect 413928 204076 413980 204128
rect 457628 204076 457680 204128
rect 301872 204008 301924 204060
rect 322388 204008 322440 204060
rect 461492 204008 461544 204060
rect 475476 204008 475528 204060
rect 20444 203940 20496 203992
rect 65248 203940 65300 203992
rect 112260 203940 112312 203992
rect 200304 203940 200356 203992
rect 200488 203940 200540 203992
rect 301780 203940 301832 203992
rect 314660 203940 314712 203992
rect 465356 203940 465408 203992
rect 19248 203872 19300 203924
rect 61384 203872 61436 203924
rect 302056 203872 302108 203924
rect 310796 203872 310848 203924
rect 312544 203872 312596 203924
rect 313280 203872 313332 203924
rect 384212 203872 384264 203924
rect 449900 203872 449952 203924
rect 473084 203940 473136 203992
rect 476028 203940 476080 203992
rect 476948 204076 477000 204128
rect 480536 204076 480588 204128
rect 478972 203940 479024 203992
rect 17868 203804 17920 203856
rect 84568 203804 84620 203856
rect 181812 203804 181864 203856
rect 187884 203804 187936 203856
rect 478880 203872 478932 203924
rect 479156 203804 479208 203856
rect 28908 203736 28960 203788
rect 34612 203736 34664 203788
rect 34704 203736 34756 203788
rect 38200 203736 38252 203788
rect 127716 203668 127768 203720
rect 200764 203668 200816 203720
rect 201868 203668 201920 203720
rect 139308 203600 139360 203652
rect 240140 203600 240192 203652
rect 269120 203600 269172 203652
rect 372620 203600 372672 203652
rect 189540 203532 189592 203584
rect 300124 203532 300176 203584
rect 469220 203532 469272 203584
rect 481916 203532 481968 203584
rect 185676 203192 185728 203244
rect 188804 203192 188856 203244
rect 17776 202852 17828 202904
rect 22376 202852 22428 202904
rect 39028 202852 39080 202904
rect 42064 202852 42116 202904
rect 399668 202852 399720 202904
rect 22008 202784 22060 202836
rect 22744 202784 22796 202836
rect 21916 202716 21968 202768
rect 53840 202784 53892 202836
rect 166356 202784 166408 202836
rect 197912 202784 197964 202836
rect 407396 202852 407448 202904
rect 410800 202852 410852 202904
rect 477500 202784 477552 202836
rect 23756 202716 23808 202768
rect 49792 202716 49844 202768
rect 170220 202716 170272 202768
rect 198832 202716 198884 202768
rect 20536 202648 20588 202700
rect 45928 202648 45980 202700
rect 187884 202648 187936 202700
rect 197360 202648 197412 202700
rect 20628 202580 20680 202632
rect 22192 202580 22244 202632
rect 39028 202580 39080 202632
rect 20168 202512 20220 202564
rect 23756 202512 23808 202564
rect 198096 202240 198148 202292
rect 197360 202172 197412 202224
rect 200488 202172 200540 202224
rect 188804 202104 188856 202156
rect 198096 202104 198148 202156
rect 200212 202104 200264 202156
rect 22744 202036 22796 202088
rect 34704 202036 34756 202088
rect 135076 201492 135128 201544
rect 198648 201424 198700 201476
rect 297732 201424 297784 201476
rect 368756 201424 368808 201476
rect 395804 201424 395856 201476
rect 483204 201424 483256 201476
rect 410800 201356 410852 201408
rect 484400 201356 484452 201408
rect 413928 201288 413980 201340
rect 484584 201288 484636 201340
rect 484584 200744 484636 200796
rect 485872 200744 485924 200796
rect 483204 200608 483256 200660
rect 484492 200608 484544 200660
rect 296536 200132 296588 200184
rect 297732 200132 297784 200184
rect 20076 200064 20128 200116
rect 107660 200064 107712 200116
rect 16488 199384 16540 199436
rect 17684 199384 17736 199436
rect 99380 199384 99432 199436
rect 18880 198704 18932 198756
rect 20076 198704 20128 198756
rect 252560 189728 252612 189780
rect 418160 189728 418212 189780
rect 118700 188980 118752 189032
rect 203064 188980 203116 189032
rect 131120 188300 131172 188352
rect 202144 188300 202196 188352
rect 203156 188300 203208 188352
rect 2780 187960 2832 188012
rect 4896 187960 4948 188012
rect 299296 187620 299348 187672
rect 360200 187620 360252 187672
rect 302148 187552 302200 187604
rect 349160 187552 349212 187604
rect 195980 187008 196032 187060
rect 300216 187008 300268 187060
rect 95884 186940 95936 186992
rect 256700 186940 256752 186992
rect 298008 186940 298060 186992
rect 312544 186940 312596 186992
rect 3332 149336 3384 149388
rect 8944 149336 8996 149388
rect 2780 136688 2832 136740
rect 5172 136688 5224 136740
rect 3332 110440 3384 110492
rect 20904 110440 20956 110492
rect 3332 84192 3384 84244
rect 20904 84192 20956 84244
rect 20904 79296 20956 79348
rect 21640 79296 21692 79348
rect 301780 78344 301832 78396
rect 314752 78344 314804 78396
rect 302700 78276 302752 78328
rect 317420 78276 317472 78328
rect 318156 78276 318208 78328
rect 301872 78208 301924 78260
rect 316776 78208 316828 78260
rect 302792 78140 302844 78192
rect 318800 78140 318852 78192
rect 430672 78140 430724 78192
rect 478236 78140 478288 78192
rect 301964 78072 302016 78124
rect 329840 78072 329892 78124
rect 394700 78072 394752 78124
rect 480536 78072 480588 78124
rect 18788 78004 18840 78056
rect 88432 78004 88484 78056
rect 191840 78004 191892 78056
rect 192944 78004 192996 78056
rect 200396 78004 200448 78056
rect 307208 78004 307260 78056
rect 479524 78004 479576 78056
rect 16396 77936 16448 77988
rect 103980 77936 104032 77988
rect 185676 77936 185728 77988
rect 198096 77936 198148 77988
rect 302056 77936 302108 77988
rect 310520 77936 310572 77988
rect 311164 77936 311216 77988
rect 579620 77936 579672 77988
rect 372712 77256 372764 77308
rect 480260 77256 480312 77308
rect 99380 77052 99432 77104
rect 100346 77052 100398 77104
rect 283840 76508 283892 76560
rect 369860 76508 369912 76560
rect 17684 75964 17736 76016
rect 99380 75964 99432 76016
rect 18880 75896 18932 75948
rect 108304 75896 108356 75948
rect 422852 75896 422904 75948
rect 483296 75896 483348 75948
rect 19064 75828 19116 75880
rect 76840 75828 76892 75880
rect 92940 75828 92992 75880
rect 96436 75828 96488 75880
rect 150900 75828 150952 75880
rect 199016 75828 199068 75880
rect 300676 75828 300728 75880
rect 340972 75828 341024 75880
rect 372620 75828 372672 75880
rect 376484 75828 376536 75880
rect 19156 75760 19208 75812
rect 73344 75760 73396 75812
rect 158628 75760 158680 75812
rect 201776 75760 201828 75812
rect 202788 75760 202840 75812
rect 316776 75760 316828 75812
rect 316960 75760 317012 75812
rect 322388 75760 322440 75812
rect 17776 75692 17828 75744
rect 69572 75692 69624 75744
rect 177948 75692 178000 75744
rect 198924 75692 198976 75744
rect 318800 75692 318852 75744
rect 326252 75760 326304 75812
rect 433984 75760 434036 75812
rect 434444 75760 434496 75812
rect 480444 75760 480496 75812
rect 438308 75692 438360 75744
rect 480720 75692 480772 75744
rect 20444 75624 20496 75676
rect 65340 75624 65392 75676
rect 442264 75624 442316 75676
rect 483020 75624 483072 75676
rect 19248 75556 19300 75608
rect 61384 75556 61436 75608
rect 449900 75556 449952 75608
rect 479156 75556 479208 75608
rect 20352 75488 20404 75540
rect 50344 75488 50396 75540
rect 414664 75488 414716 75540
rect 415124 75488 415176 75540
rect 479064 75488 479116 75540
rect 4988 75420 5040 75472
rect 23020 75420 23072 75472
rect 189540 75352 189592 75404
rect 229744 75352 229796 75404
rect 322204 75352 322256 75404
rect 333980 75352 334032 75404
rect 375380 75352 375432 75404
rect 449900 75352 449952 75404
rect 96436 75284 96488 75336
rect 112444 75284 112496 75336
rect 199016 75284 199068 75336
rect 255964 75284 256016 75336
rect 327080 75284 327132 75336
rect 345572 75284 345624 75336
rect 376760 75284 376812 75336
rect 480352 75284 480404 75336
rect 112260 75216 112312 75268
rect 139216 75216 139268 75268
rect 147036 75216 147088 75268
rect 156604 75216 156656 75268
rect 202788 75216 202840 75268
rect 288440 75216 288492 75268
rect 300584 75216 300636 75268
rect 331220 75216 331272 75268
rect 357164 75216 357216 75268
rect 378140 75216 378192 75268
rect 481916 75216 481968 75268
rect 69572 75148 69624 75200
rect 122104 75148 122156 75200
rect 139308 75148 139360 75200
rect 238760 75148 238812 75200
rect 278780 75148 278832 75200
rect 438308 75148 438360 75200
rect 271880 74604 271932 74656
rect 422852 74604 422904 74656
rect 274640 74536 274692 74588
rect 430580 74536 430632 74588
rect 17868 74468 17920 74520
rect 84936 74468 84988 74520
rect 139216 74468 139268 74520
rect 200304 74468 200356 74520
rect 201408 74468 201460 74520
rect 427084 74468 427136 74520
rect 483388 74468 483440 74520
rect 21916 74400 21968 74452
rect 54484 74400 54536 74452
rect 446404 74400 446456 74452
rect 477960 74400 478012 74452
rect 20536 74332 20588 74384
rect 46204 74332 46256 74384
rect 453764 74332 453816 74384
rect 478052 74332 478104 74384
rect 20628 74264 20680 74316
rect 42064 74264 42116 74316
rect 457628 74264 457680 74316
rect 478972 74264 479024 74316
rect 22744 74196 22796 74248
rect 38108 74196 38160 74248
rect 461492 74196 461544 74248
rect 477868 74196 477920 74248
rect 22836 74128 22888 74180
rect 35164 74128 35216 74180
rect 465724 74128 465776 74180
rect 478880 74128 478932 74180
rect 22928 74060 22980 74112
rect 31024 74060 31076 74112
rect 473084 74060 473136 74112
rect 481824 74060 481876 74112
rect 198924 73992 198976 74044
rect 307024 73992 307076 74044
rect 311164 73992 311216 74044
rect 427084 73992 427136 74044
rect 201408 73924 201460 73976
rect 227720 73924 227772 73976
rect 298652 73924 298704 73976
rect 461492 73924 461544 73976
rect 212632 73856 212684 73908
rect 395804 73856 395856 73908
rect 73344 73788 73396 73840
rect 356704 73788 356756 73840
rect 119896 73108 119948 73160
rect 203064 73108 203116 73160
rect 403624 73108 403676 73160
rect 481732 73108 481784 73160
rect 173808 73040 173860 73092
rect 198004 73040 198056 73092
rect 407764 73040 407816 73092
rect 484400 73040 484452 73092
rect 411260 72972 411312 73024
rect 411904 72972 411956 73024
rect 485872 72972 485924 73024
rect 203064 72632 203116 72684
rect 230848 72632 230900 72684
rect 293960 72632 294012 72684
rect 375380 72632 375432 72684
rect 198004 72564 198056 72616
rect 305368 72564 305420 72616
rect 330300 72564 330352 72616
rect 353300 72564 353352 72616
rect 104440 72496 104492 72548
rect 224224 72496 224276 72548
rect 254032 72496 254084 72548
rect 418988 72496 419040 72548
rect 38108 72428 38160 72480
rect 340880 72428 340932 72480
rect 131488 71680 131540 71732
rect 202144 71680 202196 71732
rect 202788 71680 202840 71732
rect 299388 71680 299440 71732
rect 329840 71680 329892 71732
rect 330300 71680 330352 71732
rect 202788 71204 202840 71256
rect 236000 71204 236052 71256
rect 270592 71204 270644 71256
rect 372620 71204 372672 71256
rect 203064 71136 203116 71188
rect 473084 71136 473136 71188
rect 88984 71068 89036 71120
rect 363328 71068 363380 71120
rect 81256 71000 81308 71052
rect 360200 71000 360252 71052
rect 127624 70320 127676 70372
rect 200764 70320 200816 70372
rect 201408 70320 201460 70372
rect 170128 70252 170180 70304
rect 198832 70252 198884 70304
rect 199384 70252 199436 70304
rect 199384 69776 199436 69828
rect 303712 69776 303764 69828
rect 201408 69708 201460 69760
rect 234160 69708 234212 69760
rect 297088 69708 297140 69760
rect 457628 69708 457680 69760
rect 76840 69640 76892 69692
rect 358360 69640 358412 69692
rect 135168 68960 135220 69012
rect 198740 68960 198792 69012
rect 300768 68960 300820 69012
rect 327080 68960 327132 69012
rect 166264 68892 166316 68944
rect 197360 68892 197412 68944
rect 198740 68552 198792 68604
rect 237472 68552 237524 68604
rect 197360 68484 197412 68536
rect 197912 68484 197964 68536
rect 302240 68484 302292 68536
rect 233884 68416 233936 68468
rect 368572 68416 368624 68468
rect 108304 68348 108356 68400
rect 225880 68348 225932 68400
rect 295432 68348 295484 68400
rect 453764 68348 453816 68400
rect 84936 68280 84988 68332
rect 361672 68280 361724 68332
rect 302884 67532 302936 67584
rect 322204 67532 322256 67584
rect 112444 66988 112496 67040
rect 255688 66988 255740 67040
rect 255964 66988 256016 67040
rect 285680 66988 285732 67040
rect 302148 66988 302200 67040
rect 328552 66988 328604 67040
rect 349160 66988 349212 67040
rect 122104 66920 122156 66972
rect 355048 66920 355100 66972
rect 54484 66852 54536 66904
rect 348424 66852 348476 66904
rect 142160 66172 142212 66224
rect 201592 66172 201644 66224
rect 202788 66172 202840 66224
rect 202788 65696 202840 65748
rect 282184 65696 282236 65748
rect 292120 65696 292172 65748
rect 446404 65696 446456 65748
rect 220912 65628 220964 65680
rect 414664 65628 414716 65680
rect 46204 65560 46256 65612
rect 345112 65560 345164 65612
rect 31024 65492 31076 65544
rect 338488 65492 338540 65544
rect 300032 64812 300084 64864
rect 387800 64812 387852 64864
rect 299296 64336 299348 64388
rect 333520 64336 333572 64388
rect 360292 64336 360344 64388
rect 57244 64268 57296 64320
rect 332600 64268 332652 64320
rect 65524 64200 65576 64252
rect 353392 64200 353444 64252
rect 61384 64132 61436 64184
rect 351920 64132 351972 64184
rect 209320 63520 209372 63572
rect 300032 63520 300084 63572
rect 156604 63452 156656 63504
rect 197820 63452 197872 63504
rect 336832 63452 336884 63504
rect 364340 63452 364392 63504
rect 99380 62976 99432 63028
rect 222568 62976 222620 63028
rect 320272 62976 320324 63028
rect 329932 62976 329984 63028
rect 219440 62908 219492 62960
rect 411904 62908 411956 62960
rect 42064 62840 42116 62892
rect 343640 62840 343692 62892
rect 35164 62772 35216 62824
rect 340144 62772 340196 62824
rect 341064 62772 341116 62824
rect 433984 62772 434036 62824
rect 197820 62092 197872 62144
rect 283840 62092 283892 62144
rect 335360 62092 335412 62144
rect 336832 62092 336884 62144
rect 5172 62024 5224 62076
rect 57060 62024 57112 62076
rect 298008 62024 298060 62076
rect 383660 62024 383712 62076
rect 207664 61548 207716 61600
rect 298008 61548 298060 61600
rect 211160 61480 211212 61532
rect 392584 61480 392636 61532
rect 214288 61412 214340 61464
rect 399484 61412 399536 61464
rect 217600 61344 217652 61396
rect 407764 61344 407816 61396
rect 114560 60664 114612 60716
rect 202972 60664 203024 60716
rect 204076 60664 204128 60716
rect 295340 60664 295392 60716
rect 296628 60664 296680 60716
rect 379520 60664 379572 60716
rect 122840 60596 122892 60648
rect 202880 60596 202932 60648
rect 204168 60596 204220 60648
rect 206008 60188 206060 60240
rect 295340 60188 295392 60240
rect 204168 60120 204220 60172
rect 232504 60120 232556 60172
rect 249064 60120 249116 60172
rect 283564 60120 283616 60172
rect 283656 60120 283708 60172
rect 386512 60120 386564 60172
rect 204076 60052 204128 60104
rect 229192 60052 229244 60104
rect 229744 60052 229796 60104
rect 364984 60052 365036 60104
rect 379888 60052 379940 60104
rect 469220 60052 469272 60104
rect 191840 59984 191892 60036
rect 204352 59984 204404 60036
rect 215944 59984 215996 60036
rect 403624 59984 403676 60036
rect 180800 59304 180852 59356
rect 200488 59304 200540 59356
rect 201408 59304 201460 59356
rect 323584 58964 323636 59016
rect 336740 58964 336792 59016
rect 296536 58828 296588 58880
rect 336832 58828 336884 58880
rect 201408 58760 201460 58812
rect 308680 58760 308732 58812
rect 325240 58760 325292 58812
rect 340972 58760 341024 58812
rect 184940 58692 184992 58744
rect 310612 58692 310664 58744
rect 368480 58692 368532 58744
rect 195980 58624 196032 58676
rect 381544 58624 381596 58676
rect 396448 58624 396500 58676
rect 476120 58624 476172 58676
rect 153200 57876 153252 57928
rect 200120 57876 200172 57928
rect 201408 57876 201460 57928
rect 258724 57876 258776 57928
rect 262680 57876 262732 57928
rect 310520 57876 310572 57928
rect 312360 57876 312412 57928
rect 161480 57808 161532 57860
rect 201500 57808 201552 57860
rect 202788 57808 202840 57860
rect 274272 57604 274324 57656
rect 311164 57604 311216 57656
rect 332600 57604 332652 57656
rect 350448 57604 350500 57656
rect 277584 57536 277636 57588
rect 341064 57536 341116 57588
rect 300124 57468 300176 57520
rect 367008 57468 367060 57520
rect 300216 57400 300268 57452
rect 383568 57400 383620 57452
rect 201408 57332 201460 57384
rect 287520 57332 287572 57384
rect 298836 57332 298888 57384
rect 385224 57332 385276 57384
rect 280896 57264 280948 57316
rect 442264 57264 442316 57316
rect 202788 57196 202840 57248
rect 290832 57196 290884 57248
rect 300768 57196 300820 57248
rect 465724 57196 465776 57248
rect 315672 56584 315724 56636
rect 317420 56584 317472 56636
rect 8944 56516 8996 56568
rect 57520 56516 57572 56568
rect 102140 52640 102192 52692
rect 104072 52640 104124 52692
rect 102140 52504 102192 52556
rect 196164 52504 196216 52556
rect 17224 52368 17276 52420
rect 57060 52368 57112 52420
rect 103060 52368 103112 52420
rect 195980 52368 196032 52420
rect 102784 51008 102836 51060
rect 195980 51008 196032 51060
rect 102600 49648 102652 49700
rect 195980 49648 196032 49700
rect 102968 48220 103020 48272
rect 195980 48220 196032 48272
rect 102232 48152 102284 48204
rect 196072 48152 196124 48204
rect 3608 46860 3660 46912
rect 57520 46860 57572 46912
rect 104072 46860 104124 46912
rect 195980 46860 196032 46912
rect 103244 45500 103296 45552
rect 195980 45500 196032 45552
rect 103060 44072 103112 44124
rect 195980 44072 196032 44124
rect 103428 44004 103480 44056
rect 196072 44004 196124 44056
rect 4896 42712 4948 42764
rect 57152 42712 57204 42764
rect 102692 42712 102744 42764
rect 195980 42712 196032 42764
rect 102784 41352 102836 41404
rect 195980 41352 196032 41404
rect 102508 39992 102560 40044
rect 195980 39992 196032 40044
rect 102324 39924 102376 39976
rect 196072 39924 196124 39976
rect 102140 38564 102192 38616
rect 196072 38564 196124 38616
rect 102416 38496 102468 38548
rect 195980 38496 196032 38548
rect 3700 37204 3752 37256
rect 57060 37204 57112 37256
rect 102232 37204 102284 37256
rect 195980 37204 196032 37256
rect 102876 35844 102928 35896
rect 195980 35844 196032 35896
rect 102140 35776 102192 35828
rect 196072 35776 196124 35828
rect 102600 34416 102652 34468
rect 195980 34416 196032 34468
rect 102784 34348 102836 34400
rect 196072 34348 196124 34400
rect 102140 33056 102192 33108
rect 195980 33056 196032 33108
rect 3332 31764 3384 31816
rect 60004 31764 60056 31816
rect 5080 31696 5132 31748
rect 57612 31696 57664 31748
rect 102324 31696 102376 31748
rect 195980 31696 196032 31748
rect 102140 31628 102192 31680
rect 196072 31628 196124 31680
rect 102232 30268 102284 30320
rect 195980 30268 196032 30320
rect 102140 30200 102192 30252
rect 196072 30200 196124 30252
rect 102140 28908 102192 28960
rect 195980 28908 196032 28960
rect 102140 28228 102192 28280
rect 195980 28228 196032 28280
rect 21456 27548 21508 27600
rect 57244 27548 57296 27600
rect 102140 27548 102192 27600
rect 195980 27548 196032 27600
rect 102784 26188 102836 26240
rect 195980 26188 196032 26240
rect 60004 24216 60056 24268
rect 335544 24216 335596 24268
rect 3516 24148 3568 24200
rect 364432 24148 364484 24200
rect 3424 24080 3476 24132
rect 367836 24080 367888 24132
rect 88984 23468 89036 23520
rect 266360 23468 266412 23520
rect 267372 23468 267424 23520
rect 3608 22720 3660 22772
rect 292580 22720 292632 22772
rect 3792 22108 3844 22160
rect 350172 22108 350224 22160
rect 62304 22040 62356 22092
rect 88984 22040 89036 22092
rect 200028 22040 200080 22092
rect 378876 22040 378928 22092
rect 389640 22040 389692 22092
rect 580264 22040 580316 22092
rect 21364 21972 21416 22024
rect 360936 21972 360988 22024
rect 393228 21972 393280 22024
rect 580356 21972 580408 22024
rect 21640 21904 21692 21956
rect 346584 21904 346636 21956
rect 396816 21904 396868 21956
rect 580448 21904 580500 21956
rect 21548 21836 21600 21888
rect 342996 21836 343048 21888
rect 386052 21836 386104 21888
rect 527824 21836 527876 21888
rect 292580 21768 292632 21820
rect 353760 21768 353812 21820
rect 382464 21768 382516 21820
rect 485780 21768 485832 21820
rect 88800 21496 88852 21548
rect 156604 21496 156656 21548
rect 149060 21428 149112 21480
rect 292764 21428 292816 21480
rect 155960 21360 156012 21412
rect 299940 21360 299992 21412
rect 178040 20068 178092 20120
rect 256884 20068 256936 20120
rect 169760 20000 169812 20052
rect 314292 20000 314344 20052
rect 138020 19932 138072 19984
rect 282000 19932 282052 19984
rect 175280 18776 175332 18828
rect 253296 18776 253348 18828
rect 150440 18708 150492 18760
rect 228180 18708 228232 18760
rect 151820 18640 151872 18692
rect 296352 18640 296404 18692
rect 184940 18572 184992 18624
rect 328644 18572 328696 18624
rect 171140 17348 171192 17400
rect 249708 17348 249760 17400
rect 131120 17280 131172 17332
rect 274824 17280 274876 17332
rect 71136 17212 71188 17264
rect 242900 17212 242952 17264
rect 168380 15988 168432 16040
rect 245660 15988 245712 16040
rect 135260 15920 135312 15972
rect 277400 15920 277452 15972
rect 74540 15852 74592 15904
rect 245936 15852 245988 15904
rect 136456 14560 136508 14612
rect 212540 14560 212592 14612
rect 164424 14492 164476 14544
rect 241520 14492 241572 14544
rect 173900 14424 173952 14476
rect 317420 14424 317472 14476
rect 139584 13200 139636 13252
rect 216680 13200 216732 13252
rect 217324 13200 217376 13252
rect 288440 13200 288492 13252
rect 160100 13132 160152 13184
rect 238760 13132 238812 13184
rect 176660 13064 176712 13116
rect 320180 13064 320232 13116
rect 153752 11908 153804 11960
rect 230480 11908 230532 11960
rect 125600 11840 125652 11892
rect 202880 11840 202932 11892
rect 186136 11772 186188 11824
rect 263600 11772 263652 11824
rect 142160 11704 142212 11756
rect 284300 11704 284352 11756
rect 147128 10412 147180 10464
rect 223580 10412 223632 10464
rect 156604 10344 156656 10396
rect 245200 10344 245252 10396
rect 3424 10276 3476 10328
rect 338120 10276 338172 10328
rect 163688 9052 163740 9104
rect 306380 9052 306432 9104
rect 167184 8984 167236 9036
rect 310520 8984 310572 9036
rect 84200 8916 84252 8968
rect 241704 8916 241756 8968
rect 157800 7760 157852 7812
rect 234620 7760 234672 7812
rect 132960 7692 133012 7744
rect 209780 7692 209832 7744
rect 188528 7624 188580 7676
rect 331220 7624 331272 7676
rect 128176 7556 128228 7608
rect 270500 7556 270552 7608
rect 143540 6264 143592 6316
rect 220820 6264 220872 6316
rect 181444 6196 181496 6248
rect 324320 6196 324372 6248
rect 78680 6128 78732 6180
rect 249984 6128 250036 6180
rect 182548 4972 182600 5024
rect 259460 4972 259512 5024
rect 129372 4904 129424 4956
rect 205640 4904 205692 4956
rect 96620 4836 96672 4888
rect 252376 4836 252428 4888
rect 92480 4768 92532 4820
rect 248788 4768 248840 4820
rect 145932 3544 145984 3596
rect 217324 3544 217376 3596
rect 151820 3476 151872 3528
rect 153016 3476 153068 3528
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 161388 3476 161440 3528
rect 302240 3476 302292 3528
rect 66260 3408 66312 3460
rect 239312 3408 239364 3460
rect 266360 3408 266412 3460
rect 579804 3408 579856 3460
rect 176660 3340 176712 3392
rect 177856 3340 177908 3392
rect 160100 2796 160152 2848
rect 161388 2796 161440 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 701010 8156 703520
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 22008 700392 22060 700398
rect 22008 700334 22060 700340
rect 3422 671256 3478 671265
rect 3422 671191 3424 671200
rect 3476 671191 3478 671200
rect 8944 671220 8996 671226
rect 3424 671162 3476 671168
rect 8944 671162 8996 671168
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 607209 2820 658135
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 2778 607200 2834 607209
rect 2778 607135 2834 607144
rect 2778 566944 2834 566953
rect 2778 566879 2834 566888
rect 2792 565962 2820 566879
rect 2780 565956 2832 565962
rect 2780 565898 2832 565904
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 502353 2820 553823
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 2778 502344 2834 502353
rect 2778 502279 2834 502288
rect 3422 502344 3478 502353
rect 3422 502279 3478 502288
rect 2792 501809 2820 502279
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 398857 2820 449511
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 410242 2912 410479
rect 2872 410236 2924 410242
rect 2872 410178 2924 410184
rect 2778 398848 2834 398857
rect 2778 398783 2834 398792
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292670 2820 293111
rect 2780 292664 2832 292670
rect 2780 292606 2832 292612
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 240174 3372 241023
rect 3332 240168 3384 240174
rect 3332 240110 3384 240116
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 2792 188018 2820 188799
rect 2780 188012 2832 188018
rect 2780 187954 2832 187960
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 149394 3372 149767
rect 3332 149388 3384 149394
rect 3332 149330 3384 149336
rect 2778 136776 2834 136785
rect 2778 136711 2780 136720
rect 2832 136711 2834 136720
rect 2780 136682 2832 136688
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3344 110498 3372 110599
rect 3332 110492 3384 110498
rect 3332 110434 3384 110440
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3344 31822 3372 32399
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3436 24138 3464 502279
rect 3514 398848 3570 398857
rect 3514 398783 3570 398792
rect 3528 397497 3556 398783
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3528 24206 3556 397423
rect 3620 332586 3648 619103
rect 4896 565956 4948 565962
rect 4896 565898 4948 565904
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3608 332580 3660 332586
rect 3608 332522 3660 332528
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3620 318850 3648 319223
rect 3608 318844 3660 318850
rect 3608 318786 3660 318792
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3620 46918 3648 267135
rect 3698 214976 3754 214985
rect 3698 214911 3754 214920
rect 3608 46912 3660 46918
rect 3608 46854 3660 46860
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3620 22778 3648 45455
rect 3712 37262 3740 214911
rect 4816 75721 4844 462538
rect 4908 204105 4936 565898
rect 7564 514820 7616 514826
rect 7564 514762 7616 514768
rect 4988 410236 5040 410242
rect 4988 410178 5040 410184
rect 4894 204096 4950 204105
rect 4894 204031 4950 204040
rect 4896 188012 4948 188018
rect 4896 187954 4948 187960
rect 4802 75712 4858 75721
rect 4802 75647 4858 75656
rect 3790 71632 3846 71641
rect 3790 71567 3846 71576
rect 3700 37256 3752 37262
rect 3700 37198 3752 37204
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3804 22166 3832 71567
rect 4908 42770 4936 187954
rect 5000 75478 5028 410178
rect 5080 292664 5132 292670
rect 5080 292606 5132 292612
rect 4988 75472 5040 75478
rect 4988 75414 5040 75420
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 5092 31754 5120 292606
rect 7576 204270 7604 514762
rect 8956 332858 8984 671162
rect 21824 586220 21876 586226
rect 21824 586162 21876 586168
rect 21640 586152 21692 586158
rect 21640 586094 21692 586100
rect 20536 586016 20588 586022
rect 20536 585958 20588 585964
rect 19246 585712 19302 585721
rect 19246 585647 19302 585656
rect 19156 572416 19208 572422
rect 19156 572358 19208 572364
rect 18880 572348 18932 572354
rect 18880 572290 18932 572296
rect 18604 461372 18656 461378
rect 18604 461314 18656 461320
rect 17776 461100 17828 461106
rect 17776 461042 17828 461048
rect 8944 332852 8996 332858
rect 8944 332794 8996 332800
rect 17788 332722 17816 461042
rect 18616 334626 18644 461314
rect 18892 461174 18920 572290
rect 19064 572280 19116 572286
rect 19064 572222 19116 572228
rect 18972 572076 19024 572082
rect 18972 572018 19024 572024
rect 18984 461378 19012 572018
rect 18972 461372 19024 461378
rect 18972 461314 19024 461320
rect 18880 461168 18932 461174
rect 18880 461110 18932 461116
rect 18788 458244 18840 458250
rect 18788 458186 18840 458192
rect 18604 334620 18656 334626
rect 18604 334562 18656 334568
rect 18616 334150 18644 334562
rect 17960 334144 18012 334150
rect 17880 334092 17960 334098
rect 17880 334086 18012 334092
rect 18604 334144 18656 334150
rect 18604 334086 18656 334092
rect 17880 334070 18000 334086
rect 16488 332716 16540 332722
rect 16488 332658 16540 332664
rect 17776 332716 17828 332722
rect 17776 332658 17828 332664
rect 16396 206304 16448 206310
rect 16396 206246 16448 206252
rect 7564 204264 7616 204270
rect 7564 204206 7616 204212
rect 8944 149388 8996 149394
rect 8944 149330 8996 149336
rect 5172 136740 5224 136746
rect 5172 136682 5224 136688
rect 5184 62082 5212 136682
rect 5172 62076 5224 62082
rect 5172 62018 5224 62024
rect 8956 56574 8984 149330
rect 16408 77994 16436 206246
rect 16500 199442 16528 332658
rect 17776 331288 17828 331294
rect 17776 331230 17828 331236
rect 17224 240168 17276 240174
rect 17224 240110 17276 240116
rect 16488 199436 16540 199442
rect 16488 199378 16540 199384
rect 16396 77988 16448 77994
rect 16396 77930 16448 77936
rect 8944 56568 8996 56574
rect 8944 56510 8996 56516
rect 17236 52426 17264 240110
rect 17788 204626 17816 331230
rect 17880 206310 17908 334070
rect 18800 329798 18828 458186
rect 18892 331090 18920 461110
rect 18984 461038 19012 461314
rect 18972 461032 19024 461038
rect 18972 460974 19024 460980
rect 19076 460934 19104 572222
rect 18984 460906 19104 460934
rect 18984 459474 19012 460906
rect 18972 459468 19024 459474
rect 18972 459410 19024 459416
rect 18984 345014 19012 459410
rect 19168 459066 19196 572358
rect 19260 459406 19288 585647
rect 20352 572212 20404 572218
rect 20352 572154 20404 572160
rect 19984 572144 20036 572150
rect 19984 572086 20036 572092
rect 19996 461106 20024 572086
rect 20260 465792 20312 465798
rect 20260 465734 20312 465740
rect 20168 461576 20220 461582
rect 20168 461518 20220 461524
rect 19984 461100 20036 461106
rect 19984 461042 20036 461048
rect 20180 460970 20208 461518
rect 20168 460964 20220 460970
rect 20168 460906 20220 460912
rect 19248 459400 19300 459406
rect 19248 459342 19300 459348
rect 19156 459060 19208 459066
rect 19156 459002 19208 459008
rect 19260 458250 19288 459342
rect 19248 458244 19300 458250
rect 19248 458186 19300 458192
rect 20180 345014 20208 460906
rect 20272 458114 20300 465734
rect 20364 459338 20392 572154
rect 20444 572008 20496 572014
rect 20444 571950 20496 571956
rect 20456 461582 20484 571950
rect 20548 465798 20576 585958
rect 20628 583024 20680 583030
rect 20628 582966 20680 582972
rect 20536 465792 20588 465798
rect 20536 465734 20588 465740
rect 20444 461576 20496 461582
rect 20444 461518 20496 461524
rect 20352 459332 20404 459338
rect 20352 459274 20404 459280
rect 20260 458108 20312 458114
rect 20260 458050 20312 458056
rect 18984 344986 19288 345014
rect 19260 334082 19288 344986
rect 20088 344986 20208 345014
rect 19248 334076 19300 334082
rect 19248 334018 19300 334024
rect 19156 334008 19208 334014
rect 19156 333950 19208 333956
rect 18880 331084 18932 331090
rect 18880 331026 18932 331032
rect 18788 329792 18840 329798
rect 18788 329734 18840 329740
rect 17868 206304 17920 206310
rect 17868 206246 17920 206252
rect 17788 204598 17908 204626
rect 17880 203862 17908 204598
rect 18892 204241 18920 331026
rect 18972 329792 19024 329798
rect 18972 329734 19024 329740
rect 18878 204232 18934 204241
rect 18878 204167 18934 204176
rect 17868 203856 17920 203862
rect 17868 203798 17920 203804
rect 17776 202904 17828 202910
rect 17776 202846 17828 202852
rect 17684 199436 17736 199442
rect 17684 199378 17736 199384
rect 17696 76022 17724 199378
rect 17684 76016 17736 76022
rect 17684 75958 17736 75964
rect 17788 75750 17816 202846
rect 17776 75744 17828 75750
rect 17776 75686 17828 75692
rect 17880 74526 17908 203798
rect 18892 200114 18920 204167
rect 18984 204066 19012 329734
rect 19064 204196 19116 204202
rect 19064 204138 19116 204144
rect 18972 204060 19024 204066
rect 18972 204002 19024 204008
rect 18800 200086 18920 200114
rect 18800 78062 18828 200086
rect 18880 198756 18932 198762
rect 18880 198698 18932 198704
rect 18788 78056 18840 78062
rect 18788 77998 18840 78004
rect 18892 75954 18920 198698
rect 18880 75948 18932 75954
rect 18880 75890 18932 75896
rect 19076 75886 19104 204138
rect 19168 204134 19196 333950
rect 19260 204202 19288 334018
rect 20088 332654 20116 344986
rect 20272 335354 20300 458050
rect 20180 335326 20300 335354
rect 20076 332648 20128 332654
rect 20076 332590 20128 332596
rect 19248 204196 19300 204202
rect 19248 204138 19300 204144
rect 19156 204128 19208 204134
rect 19156 204070 19208 204076
rect 19064 75880 19116 75886
rect 19064 75822 19116 75828
rect 19168 75818 19196 204070
rect 19248 204060 19300 204066
rect 19248 204002 19300 204008
rect 19260 203930 19288 204002
rect 19248 203924 19300 203930
rect 19248 203866 19300 203872
rect 19156 75812 19208 75818
rect 19156 75754 19208 75760
rect 19260 75614 19288 203866
rect 20088 200122 20116 332590
rect 20180 332518 20208 335326
rect 20364 332790 20392 459274
rect 20444 459060 20496 459066
rect 20444 459002 20496 459008
rect 20456 458930 20484 459002
rect 20640 458998 20668 582966
rect 21652 460873 21680 586094
rect 21732 585948 21784 585954
rect 21732 585890 21784 585896
rect 21638 460864 21694 460873
rect 21638 460799 21694 460808
rect 20628 458992 20680 458998
rect 20628 458934 20680 458940
rect 21456 458992 21508 458998
rect 21456 458934 21508 458940
rect 20444 458924 20496 458930
rect 20444 458866 20496 458872
rect 20352 332784 20404 332790
rect 20352 332726 20404 332732
rect 20168 332512 20220 332518
rect 20168 332454 20220 332460
rect 20180 202570 20208 332454
rect 20260 329792 20312 329798
rect 20260 329734 20312 329740
rect 20272 204626 20300 329734
rect 20364 205737 20392 332726
rect 20456 329798 20484 458866
rect 21468 458862 21496 458934
rect 21456 458856 21508 458862
rect 21456 458798 21508 458804
rect 20536 456816 20588 456822
rect 20536 456758 20588 456764
rect 20548 332450 20576 456758
rect 20904 345092 20956 345098
rect 20904 345034 20956 345040
rect 20916 335354 20944 345034
rect 20916 335326 21404 335354
rect 20536 332444 20588 332450
rect 20536 332386 20588 332392
rect 20444 329792 20496 329798
rect 20444 329734 20496 329740
rect 20350 205728 20406 205737
rect 20350 205663 20352 205672
rect 20404 205663 20406 205672
rect 20352 205634 20404 205640
rect 20364 205603 20392 205634
rect 20272 204598 20484 204626
rect 20456 203998 20484 204598
rect 20444 203992 20496 203998
rect 20444 203934 20496 203940
rect 20168 202564 20220 202570
rect 20168 202506 20220 202512
rect 20076 200116 20128 200122
rect 20180 200114 20208 202506
rect 20180 200086 20392 200114
rect 20076 200058 20128 200064
rect 20088 198762 20116 200058
rect 20076 198756 20128 198762
rect 20076 198698 20128 198704
rect 19248 75608 19300 75614
rect 19248 75550 19300 75556
rect 20364 75546 20392 200086
rect 20456 75682 20484 203934
rect 20548 202706 20576 332386
rect 20536 202700 20588 202706
rect 20536 202642 20588 202648
rect 20444 75676 20496 75682
rect 20444 75618 20496 75624
rect 20352 75540 20404 75546
rect 20352 75482 20404 75488
rect 17868 74520 17920 74526
rect 17868 74462 17920 74468
rect 20548 74390 20576 202642
rect 20628 202632 20680 202638
rect 20628 202574 20680 202580
rect 20536 74384 20588 74390
rect 20536 74326 20588 74332
rect 20640 74322 20668 202574
rect 20904 110492 20956 110498
rect 20904 110434 20956 110440
rect 20916 110401 20944 110434
rect 20902 110392 20958 110401
rect 20902 110327 20958 110336
rect 20904 84244 20956 84250
rect 20904 84186 20956 84192
rect 20916 79354 20944 84186
rect 20904 79348 20956 79354
rect 20904 79290 20956 79296
rect 20628 74316 20680 74322
rect 20628 74258 20680 74264
rect 17224 52420 17276 52426
rect 17224 52362 17276 52368
rect 5080 31748 5132 31754
rect 5080 31690 5132 31696
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 21376 22030 21404 335326
rect 21468 334694 21496 458798
rect 21548 443964 21600 443970
rect 21548 443906 21600 443912
rect 21456 334688 21508 334694
rect 21456 334630 21508 334636
rect 21468 334014 21496 334630
rect 21456 334008 21508 334014
rect 21456 333950 21508 333956
rect 21560 331294 21588 443906
rect 21548 331288 21600 331294
rect 21548 331230 21600 331236
rect 21652 331022 21680 460799
rect 21744 457978 21772 585890
rect 21732 457972 21784 457978
rect 21732 457914 21784 457920
rect 21744 451274 21772 457914
rect 21836 457502 21864 586162
rect 21916 585880 21968 585886
rect 21916 585822 21968 585828
rect 21928 458046 21956 585822
rect 22020 459542 22048 700334
rect 22192 700324 22244 700330
rect 22192 700266 22244 700272
rect 22100 699712 22152 699718
rect 22100 699654 22152 699660
rect 22112 462670 22140 699654
rect 22204 596174 22232 700266
rect 24320 699718 24348 703520
rect 72988 701010 73016 703520
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 72988 700369 73016 700946
rect 89180 700398 89208 703520
rect 137848 700398 137876 703520
rect 89168 700392 89220 700398
rect 72974 700360 73030 700369
rect 89168 700334 89220 700340
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 154132 700330 154160 703520
rect 198740 700392 198792 700398
rect 198740 700334 198792 700340
rect 72974 700295 73030 700304
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 198752 699854 198780 700334
rect 202800 699854 202828 703520
rect 198740 699848 198792 699854
rect 198740 699790 198792 699796
rect 200028 699848 200080 699854
rect 200028 699790 200080 699796
rect 202788 699848 202840 699854
rect 202788 699790 202840 699796
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 22204 596146 22692 596174
rect 22664 588690 22692 596146
rect 22664 588662 23092 588690
rect 26956 587302 27292 587330
rect 27264 586401 27292 587302
rect 30484 587302 30820 587330
rect 34532 587302 34684 587330
rect 38212 587302 38548 587330
rect 42076 587302 42412 587330
rect 45940 587302 46276 587330
rect 49804 587302 50140 587330
rect 53852 587302 54004 587330
rect 57532 587302 57868 587330
rect 61396 587302 61732 587330
rect 65260 587302 65596 587330
rect 69032 587302 69460 587330
rect 73172 587302 73324 587330
rect 75932 587302 77188 587330
rect 80072 587302 81052 587330
rect 84580 587302 84916 587330
rect 88444 587302 88780 587330
rect 92644 587302 92980 587330
rect 27250 586392 27306 586401
rect 27250 586327 27306 586336
rect 22928 586084 22980 586090
rect 22928 586026 22980 586032
rect 22836 585812 22888 585818
rect 22836 585754 22888 585760
rect 22100 462664 22152 462670
rect 22100 462606 22152 462612
rect 22848 460934 22876 585754
rect 22664 460906 22876 460934
rect 22008 459536 22060 459542
rect 22664 459513 22692 460906
rect 22008 459478 22060 459484
rect 22650 459504 22706 459513
rect 22650 459439 22706 459448
rect 21916 458040 21968 458046
rect 21916 457982 21968 457988
rect 21824 457496 21876 457502
rect 21824 457438 21876 457444
rect 21744 451246 22048 451274
rect 22020 335354 22048 451246
rect 22664 335354 22692 459439
rect 22744 458992 22796 458998
rect 22744 458934 22796 458940
rect 22756 458046 22784 458934
rect 22940 458046 22968 586026
rect 30484 585886 30512 587302
rect 34532 586226 34560 587302
rect 34520 586220 34572 586226
rect 34520 586162 34572 586168
rect 30472 585880 30524 585886
rect 30472 585822 30524 585828
rect 32404 585880 32456 585886
rect 32404 585822 32456 585828
rect 32416 572422 32444 585822
rect 38212 585818 38240 587302
rect 42076 586158 42104 587302
rect 42064 586152 42116 586158
rect 42064 586094 42116 586100
rect 45940 586090 45968 587302
rect 45928 586084 45980 586090
rect 45928 586026 45980 586032
rect 49804 586022 49832 587302
rect 49792 586016 49844 586022
rect 49792 585958 49844 585964
rect 53852 585954 53880 587302
rect 53840 585948 53892 585954
rect 53840 585890 53892 585896
rect 57532 585857 57560 587302
rect 57518 585848 57574 585857
rect 38200 585812 38252 585818
rect 38200 585754 38252 585760
rect 39304 585812 39356 585818
rect 57518 585783 57574 585792
rect 39304 585754 39356 585760
rect 32404 572416 32456 572422
rect 32404 572358 32456 572364
rect 39316 572354 39344 585754
rect 61396 585721 61424 587302
rect 65260 585886 65288 587302
rect 65248 585880 65300 585886
rect 65248 585822 65300 585828
rect 61382 585712 61438 585721
rect 61382 585647 61438 585656
rect 39304 572348 39356 572354
rect 39304 572290 39356 572296
rect 69032 571985 69060 587302
rect 73172 583030 73200 587302
rect 73160 583024 73212 583030
rect 73160 582966 73212 582972
rect 75932 572286 75960 587302
rect 75920 572280 75972 572286
rect 75920 572222 75972 572228
rect 80072 572218 80100 587302
rect 84580 583001 84608 587302
rect 88444 585818 88472 587302
rect 92952 586498 92980 587302
rect 96172 587302 96508 587330
rect 99392 587302 100372 587330
rect 103532 587302 104236 587330
rect 107672 587302 108100 587330
rect 111964 587302 112300 587330
rect 96172 586498 96200 587302
rect 92940 586492 92992 586498
rect 92940 586434 92992 586440
rect 96160 586492 96212 586498
rect 96160 586434 96212 586440
rect 88432 585812 88484 585818
rect 88432 585754 88484 585760
rect 96172 585721 96200 586434
rect 96158 585712 96214 585721
rect 96158 585647 96214 585656
rect 84566 582992 84622 583001
rect 84566 582927 84622 582936
rect 80060 572212 80112 572218
rect 80060 572154 80112 572160
rect 99392 572150 99420 587302
rect 99380 572144 99432 572150
rect 99380 572086 99432 572092
rect 103532 572082 103560 587302
rect 103520 572076 103572 572082
rect 103520 572018 103572 572024
rect 107672 572014 107700 587302
rect 112272 583001 112300 587302
rect 114572 587302 115828 587330
rect 118712 587302 119692 587330
rect 123556 587302 123892 587330
rect 127420 587302 127756 587330
rect 112258 582992 112314 583001
rect 112258 582927 112314 582936
rect 114572 572150 114600 587302
rect 118712 572218 118740 587302
rect 123864 583030 123892 587302
rect 127728 583098 127756 587302
rect 131132 587302 131284 587330
rect 133892 587302 135148 587330
rect 138032 587302 139012 587330
rect 142876 587302 143212 587330
rect 146740 587302 147076 587330
rect 150604 587302 150940 587330
rect 127716 583092 127768 583098
rect 127716 583034 127768 583040
rect 123852 583024 123904 583030
rect 123852 582966 123904 582972
rect 131132 572286 131160 587302
rect 131120 572280 131172 572286
rect 131120 572222 131172 572228
rect 118700 572212 118752 572218
rect 118700 572154 118752 572160
rect 114560 572144 114612 572150
rect 133892 572121 133920 587302
rect 114560 572086 114612 572092
rect 133878 572112 133934 572121
rect 133878 572047 133934 572056
rect 138032 572014 138060 587302
rect 143184 583166 143212 587302
rect 147048 583234 147076 587302
rect 150912 583302 150940 587302
rect 153212 587302 154468 587330
rect 158332 587302 158668 587330
rect 150900 583296 150952 583302
rect 150900 583238 150952 583244
rect 147036 583228 147088 583234
rect 147036 583170 147088 583176
rect 143172 583160 143224 583166
rect 143172 583102 143224 583108
rect 153212 572354 153240 587302
rect 158640 583370 158668 587302
rect 161492 587302 162196 587330
rect 166060 587302 166396 587330
rect 169924 587302 170260 587330
rect 158628 583364 158680 583370
rect 158628 583306 158680 583312
rect 161492 572422 161520 587302
rect 166368 585818 166396 587302
rect 170232 585886 170260 587302
rect 173774 587058 173802 587316
rect 177652 587302 177988 587330
rect 181516 587302 181852 587330
rect 185380 587302 185716 587330
rect 173774 587030 173848 587058
rect 173820 585954 173848 587030
rect 177960 586022 177988 587302
rect 181824 586090 181852 587302
rect 185688 586158 185716 587302
rect 189092 587302 189244 587330
rect 185676 586152 185728 586158
rect 185676 586094 185728 586100
rect 181812 586084 181864 586090
rect 181812 586026 181864 586032
rect 177948 586016 178000 586022
rect 177948 585958 178000 585964
rect 173808 585948 173860 585954
rect 173808 585890 173860 585896
rect 170220 585880 170272 585886
rect 170220 585822 170272 585828
rect 166356 585812 166408 585818
rect 166356 585754 166408 585760
rect 161480 572416 161532 572422
rect 161480 572358 161532 572364
rect 153200 572348 153252 572354
rect 153200 572290 153252 572296
rect 189092 572082 189120 587302
rect 193094 587058 193122 587316
rect 195992 587302 196972 587330
rect 193094 587030 193168 587058
rect 193140 586226 193168 587030
rect 193128 586220 193180 586226
rect 193128 586162 193180 586168
rect 189080 572076 189132 572082
rect 189080 572018 189132 572024
rect 107660 572008 107712 572014
rect 69018 571976 69074 571985
rect 107660 571950 107712 571956
rect 138020 572008 138072 572014
rect 195992 571985 196020 587302
rect 198096 586084 198148 586090
rect 198096 586026 198148 586032
rect 198004 585948 198056 585954
rect 198004 585890 198056 585896
rect 197912 585812 197964 585818
rect 197912 585754 197964 585760
rect 138020 571950 138072 571956
rect 195978 571976 196034 571985
rect 69018 571911 69074 571920
rect 195978 571911 196034 571920
rect 23204 462664 23256 462670
rect 23092 462612 23204 462618
rect 23092 462606 23256 462612
rect 23092 462590 23244 462606
rect 26620 461230 26956 461258
rect 30484 461230 30820 461258
rect 34532 461230 34684 461258
rect 38212 461230 38548 461258
rect 42076 461230 42412 461258
rect 45940 461230 46276 461258
rect 49804 461230 50140 461258
rect 53852 461230 54004 461258
rect 57532 461230 57868 461258
rect 61396 461230 61732 461258
rect 65260 461230 65596 461258
rect 69124 461230 69460 461258
rect 73172 461230 73324 461258
rect 76852 461230 77188 461258
rect 80716 461230 81052 461258
rect 84580 461230 84916 461258
rect 88444 461230 88780 461258
rect 92644 461230 92980 461258
rect 26620 459542 26648 461230
rect 26608 459536 26660 459542
rect 26608 459478 26660 459484
rect 30484 458998 30512 461230
rect 30472 458992 30524 458998
rect 30472 458934 30524 458940
rect 23478 458824 23534 458833
rect 23478 458759 23534 458768
rect 22744 458040 22796 458046
rect 22744 457982 22796 457988
rect 22928 458040 22980 458046
rect 22928 457982 22980 457988
rect 21928 335326 22048 335354
rect 22572 335326 22692 335354
rect 21928 332178 21956 335326
rect 22572 332382 22600 335326
rect 22756 333418 22784 457982
rect 22836 457496 22888 457502
rect 22836 457438 22888 457444
rect 22664 333390 22784 333418
rect 22560 332376 22612 332382
rect 22560 332318 22612 332324
rect 21916 332172 21968 332178
rect 21916 332114 21968 332120
rect 21640 331016 21692 331022
rect 21640 330958 21692 330964
rect 21456 318844 21508 318850
rect 21456 318786 21508 318792
rect 21468 27606 21496 318786
rect 21928 202774 21956 332114
rect 22192 331900 22244 331906
rect 22192 331842 22244 331848
rect 22008 331492 22060 331498
rect 22008 331434 22060 331440
rect 22020 202842 22048 331434
rect 22204 331022 22232 331842
rect 22572 331498 22600 332318
rect 22664 332246 22692 333390
rect 22848 332314 22876 457438
rect 22940 456822 22968 457982
rect 22928 456816 22980 456822
rect 22928 456758 22980 456764
rect 23492 443970 23520 458759
rect 34532 458522 34560 461230
rect 38212 459513 38240 461230
rect 42076 460873 42104 461230
rect 42062 460864 42118 460873
rect 42062 460799 42118 460808
rect 38198 459504 38254 459513
rect 38198 459439 38254 459448
rect 45940 459066 45968 461230
rect 42800 459060 42852 459066
rect 42800 459002 42852 459008
rect 45928 459060 45980 459066
rect 45928 459002 45980 459008
rect 30380 458516 30432 458522
rect 30380 458458 30432 458464
rect 34520 458516 34572 458522
rect 34520 458458 34572 458464
rect 30392 457502 30420 458458
rect 42812 458046 42840 459002
rect 49804 458114 49832 461230
rect 49792 458108 49844 458114
rect 49792 458050 49844 458056
rect 42800 458040 42852 458046
rect 42800 457982 42852 457988
rect 53852 457978 53880 461230
rect 57532 458153 57560 461230
rect 61396 459406 61424 461230
rect 61384 459400 61436 459406
rect 61384 459342 61436 459348
rect 65260 458930 65288 461230
rect 69124 458969 69152 461230
rect 69110 458960 69166 458969
rect 65248 458924 65300 458930
rect 69110 458895 69166 458904
rect 65248 458866 65300 458872
rect 73172 458862 73200 461230
rect 76852 459474 76880 461230
rect 76840 459468 76892 459474
rect 76840 459410 76892 459416
rect 80716 459338 80744 461230
rect 80704 459332 80756 459338
rect 80704 459274 80756 459280
rect 73160 458856 73212 458862
rect 84580 458833 84608 461230
rect 88444 461174 88472 461230
rect 88432 461168 88484 461174
rect 88432 461110 88484 461116
rect 92952 459542 92980 461230
rect 96172 461230 96508 461258
rect 96172 460934 96200 461230
rect 100358 461106 100386 461244
rect 100346 461100 100398 461106
rect 100346 461042 100398 461048
rect 104222 461038 104250 461244
rect 107764 461230 108100 461258
rect 111964 461230 112300 461258
rect 104210 461032 104262 461038
rect 104210 460974 104262 460980
rect 107764 460970 107792 461230
rect 95896 460906 96200 460934
rect 107752 460964 107804 460970
rect 107752 460906 107804 460912
rect 95896 459542 95924 460906
rect 92940 459536 92992 459542
rect 92940 459478 92992 459484
rect 95884 459536 95936 459542
rect 95884 459478 95936 459484
rect 73160 458798 73212 458804
rect 84566 458824 84622 458833
rect 84566 458759 84622 458768
rect 57518 458144 57574 458153
rect 57518 458079 57574 458088
rect 53840 457972 53892 457978
rect 53840 457914 53892 457920
rect 30380 457496 30432 457502
rect 30380 457438 30432 457444
rect 23480 443964 23532 443970
rect 23480 443906 23532 443912
rect 95896 443698 95924 459478
rect 112272 458153 112300 461230
rect 115814 461122 115842 461244
rect 119692 461230 120028 461258
rect 123556 461230 123892 461258
rect 115814 461094 115888 461122
rect 115860 459542 115888 461094
rect 115848 459536 115900 459542
rect 115848 459478 115900 459484
rect 120000 458930 120028 461230
rect 123864 460970 123892 461230
rect 126992 461230 127420 461258
rect 131284 461230 131620 461258
rect 123852 460964 123904 460970
rect 123852 460906 123904 460912
rect 119988 458924 120040 458930
rect 119988 458866 120040 458872
rect 112258 458144 112314 458153
rect 112258 458079 112314 458088
rect 126992 444378 127020 461230
rect 131592 459474 131620 461230
rect 135134 461122 135162 461244
rect 139012 461230 139348 461258
rect 135134 461094 135208 461122
rect 131580 459468 131632 459474
rect 131580 459410 131632 459416
rect 135180 459406 135208 461094
rect 135168 459400 135220 459406
rect 135168 459342 135220 459348
rect 139320 458862 139348 461230
rect 142862 461038 142890 461244
rect 146726 461106 146754 461244
rect 150604 461230 150940 461258
rect 146714 461100 146766 461106
rect 146714 461042 146766 461048
rect 142850 461032 142902 461038
rect 142850 460974 142902 460980
rect 139308 458856 139360 458862
rect 139308 458798 139360 458804
rect 150912 458182 150940 461230
rect 154454 461122 154482 461244
rect 158332 461230 158668 461258
rect 162196 461230 162532 461258
rect 166060 461230 166396 461258
rect 169924 461230 170260 461258
rect 158640 461174 158668 461230
rect 158628 461168 158680 461174
rect 154454 461094 154528 461122
rect 158628 461110 158680 461116
rect 154500 458998 154528 461094
rect 162504 459338 162532 461230
rect 162492 459332 162544 459338
rect 162492 459274 162544 459280
rect 154488 458992 154540 458998
rect 154488 458934 154540 458940
rect 150900 458176 150952 458182
rect 150900 458118 150952 458124
rect 166368 458114 166396 461230
rect 166356 458108 166408 458114
rect 166356 458050 166408 458056
rect 170232 458046 170260 461230
rect 173774 461122 173802 461244
rect 177652 461230 177988 461258
rect 181516 461230 181852 461258
rect 185380 461230 185716 461258
rect 189244 461230 189580 461258
rect 173774 461094 173848 461122
rect 170220 458040 170272 458046
rect 173820 458017 173848 461094
rect 177960 460902 177988 461230
rect 177948 460896 178000 460902
rect 181824 460873 181852 461230
rect 177948 460838 178000 460844
rect 181810 460864 181866 460873
rect 181810 460799 181866 460808
rect 185688 460737 185716 461230
rect 185674 460728 185730 460737
rect 185674 460663 185730 460672
rect 189552 458833 189580 461230
rect 193094 461122 193122 461244
rect 196972 461230 197308 461258
rect 193094 461094 193168 461122
rect 193140 459513 193168 461094
rect 193126 459504 193182 459513
rect 193126 459439 193182 459448
rect 197280 458969 197308 461230
rect 197360 459400 197412 459406
rect 197358 459368 197360 459377
rect 197412 459368 197414 459377
rect 197358 459303 197414 459312
rect 197266 458960 197322 458969
rect 197176 458924 197228 458930
rect 197266 458895 197322 458904
rect 197176 458866 197228 458872
rect 189538 458824 189594 458833
rect 189538 458759 189594 458768
rect 170220 457982 170272 457988
rect 173806 458008 173862 458017
rect 173806 457943 173862 457952
rect 197188 451274 197216 458866
rect 197924 458114 197952 585754
rect 197912 458108 197964 458114
rect 197912 458050 197964 458056
rect 197924 456822 197952 458050
rect 198016 458017 198044 585890
rect 198108 480254 198136 586026
rect 198924 586016 198976 586022
rect 198924 585958 198976 585964
rect 198740 585880 198792 585886
rect 198740 585822 198792 585828
rect 198108 480226 198228 480254
rect 198200 460873 198228 480226
rect 198186 460864 198242 460873
rect 198186 460799 198242 460808
rect 198002 458008 198058 458017
rect 198002 457943 198058 457952
rect 197912 456816 197964 456822
rect 197912 456758 197964 456764
rect 197188 451246 197308 451274
rect 126980 444372 127032 444378
rect 126980 444314 127032 444320
rect 197280 443766 197308 451246
rect 197268 443760 197320 443766
rect 197268 443702 197320 443708
rect 95884 443692 95936 443698
rect 95884 443634 95936 443640
rect 72976 334688 73028 334694
rect 73028 334636 73324 334642
rect 72976 334630 73324 334636
rect 72988 334614 73324 334630
rect 103900 334626 104236 334642
rect 103888 334620 104236 334626
rect 103940 334614 104236 334620
rect 103888 334562 103940 334568
rect 76840 334008 76892 334014
rect 76892 333956 77188 333962
rect 76840 333950 77188 333956
rect 76852 333934 77188 333950
rect 96448 333390 96508 333418
rect 22940 333254 23092 333282
rect 26620 333254 26956 333282
rect 30484 333254 30820 333282
rect 34532 333254 34684 333282
rect 38212 333254 38548 333282
rect 42076 333254 42412 333282
rect 45940 333254 46276 333282
rect 49804 333254 50140 333282
rect 53852 333254 54004 333282
rect 57532 333254 57868 333282
rect 61396 333254 61732 333282
rect 65260 333254 65596 333282
rect 69124 333254 69460 333282
rect 80716 333254 81052 333282
rect 84580 333254 84916 333282
rect 88444 333254 88780 333282
rect 92644 333254 92980 333282
rect 22940 332586 22968 333254
rect 26620 332858 26648 333254
rect 26608 332852 26660 332858
rect 26608 332794 26660 332800
rect 22928 332580 22980 332586
rect 22928 332522 22980 332528
rect 22836 332308 22888 332314
rect 22836 332250 22888 332256
rect 22652 332240 22704 332246
rect 22652 332182 22704 332188
rect 22560 331492 22612 331498
rect 22560 331434 22612 331440
rect 22664 331294 22692 332182
rect 22652 331288 22704 331294
rect 22652 331230 22704 331236
rect 22192 331016 22244 331022
rect 22192 330958 22244 330964
rect 22008 202836 22060 202842
rect 22008 202778 22060 202784
rect 21916 202768 21968 202774
rect 21916 202710 21968 202716
rect 21546 110392 21602 110401
rect 21546 110327 21602 110336
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21560 21894 21588 110327
rect 21640 79348 21692 79354
rect 21640 79290 21692 79296
rect 21652 21962 21680 79290
rect 21928 74458 21956 202710
rect 22204 202638 22232 330958
rect 22848 203561 22876 332250
rect 30484 332246 30512 333254
rect 34532 332314 34560 333254
rect 38212 332382 38240 333254
rect 38200 332376 38252 332382
rect 38200 332318 38252 332324
rect 34520 332308 34572 332314
rect 34520 332250 34572 332256
rect 30472 332240 30524 332246
rect 30472 332182 30524 332188
rect 42076 331906 42104 333254
rect 45940 332450 45968 333254
rect 49804 332518 49832 333254
rect 49792 332512 49844 332518
rect 49792 332454 49844 332460
rect 45928 332444 45980 332450
rect 45928 332386 45980 332392
rect 53852 332178 53880 333254
rect 57532 332353 57560 333254
rect 57518 332344 57574 332353
rect 57518 332279 57574 332288
rect 53840 332172 53892 332178
rect 53840 332114 53892 332120
rect 42064 331900 42116 331906
rect 42064 331842 42116 331848
rect 22928 331288 22980 331294
rect 22928 331230 22980 331236
rect 22940 204270 22968 331230
rect 61396 329730 61424 333254
rect 65260 329798 65288 333254
rect 69124 332489 69152 333254
rect 80716 332790 80744 333254
rect 80704 332784 80756 332790
rect 80704 332726 80756 332732
rect 69110 332480 69166 332489
rect 69110 332415 69166 332424
rect 84580 331294 84608 333254
rect 84568 331288 84620 331294
rect 84568 331230 84620 331236
rect 88444 331090 88472 333254
rect 92952 332586 92980 333254
rect 96448 332586 96476 333390
rect 100036 333254 100372 333282
rect 107764 333254 108100 333282
rect 111812 333254 111964 333282
rect 114572 333254 115828 333282
rect 119692 333254 120028 333282
rect 123556 333254 123892 333282
rect 127420 333254 127756 333282
rect 100036 332722 100064 333254
rect 100024 332716 100076 332722
rect 100024 332658 100076 332664
rect 107764 332654 107792 333254
rect 107752 332648 107804 332654
rect 107752 332590 107804 332596
rect 92940 332580 92992 332586
rect 92940 332522 92992 332528
rect 96436 332580 96488 332586
rect 96436 332522 96488 332528
rect 96448 331809 96476 332522
rect 96434 331800 96490 331809
rect 96434 331735 96490 331744
rect 88432 331084 88484 331090
rect 88432 331026 88484 331032
rect 65248 329792 65300 329798
rect 65248 329734 65300 329740
rect 61384 329724 61436 329730
rect 61384 329666 61436 329672
rect 111812 315382 111840 333254
rect 114572 315994 114600 333254
rect 120000 330546 120028 333254
rect 123864 332654 123892 333254
rect 123852 332648 123904 332654
rect 123852 332590 123904 332596
rect 127728 331226 127756 333254
rect 131132 333254 131284 333282
rect 135088 333254 135148 333282
rect 138032 333254 139012 333282
rect 142876 333254 143212 333282
rect 146740 333254 147076 333282
rect 131132 331242 131160 333254
rect 135088 332586 135116 333254
rect 137928 332784 137980 332790
rect 137928 332726 137980 332732
rect 137940 332586 137968 332726
rect 135076 332580 135128 332586
rect 135076 332522 135128 332528
rect 137928 332580 137980 332586
rect 137928 332522 137980 332528
rect 127716 331220 127768 331226
rect 127716 331162 127768 331168
rect 131040 331214 131160 331242
rect 119988 330540 120040 330546
rect 119988 330482 120040 330488
rect 131040 329798 131068 331214
rect 131028 329792 131080 329798
rect 131028 329734 131080 329740
rect 138032 316742 138060 333254
rect 143184 332722 143212 333254
rect 143172 332716 143224 332722
rect 143172 332658 143224 332664
rect 147048 330614 147076 333254
rect 150452 333254 150604 333282
rect 154468 333254 154804 333282
rect 158332 333254 158760 333282
rect 162196 333254 162532 333282
rect 166060 333254 166396 333282
rect 169924 333254 170260 333282
rect 150452 331242 150480 333254
rect 154776 332858 154804 333254
rect 158732 332926 158760 333254
rect 162504 332994 162532 333254
rect 162492 332988 162544 332994
rect 162492 332930 162544 332936
rect 158720 332920 158772 332926
rect 158720 332862 158772 332868
rect 154764 332852 154816 332858
rect 154764 332794 154816 332800
rect 166368 332586 166396 333254
rect 166356 332580 166408 332586
rect 166356 332522 166408 332528
rect 170232 332518 170260 333254
rect 173728 333254 173788 333282
rect 177652 333254 177988 333282
rect 181516 333254 181852 333282
rect 185380 333254 185716 333282
rect 189244 333254 189580 333282
rect 170220 332512 170272 332518
rect 170220 332454 170272 332460
rect 173728 332450 173756 333254
rect 173716 332444 173768 332450
rect 173716 332386 173768 332392
rect 177960 332382 177988 333254
rect 177948 332376 178000 332382
rect 177948 332318 178000 332324
rect 181824 332314 181852 333254
rect 181812 332308 181864 332314
rect 181812 332250 181864 332256
rect 185688 332246 185716 333254
rect 185676 332240 185728 332246
rect 185676 332182 185728 332188
rect 189552 331945 189580 333254
rect 193048 333254 193108 333282
rect 195992 333254 196972 333282
rect 193048 332178 193076 333254
rect 193036 332172 193088 332178
rect 193036 332114 193088 332120
rect 189538 331936 189594 331945
rect 189538 331871 189594 331880
rect 150360 331214 150480 331242
rect 147036 330608 147088 330614
rect 147036 330550 147088 330556
rect 138020 316736 138072 316742
rect 138020 316678 138072 316684
rect 114560 315988 114612 315994
rect 114560 315930 114612 315936
rect 150360 315926 150388 331214
rect 150348 315920 150400 315926
rect 150348 315862 150400 315868
rect 111800 315376 111852 315382
rect 111800 315318 111852 315324
rect 195992 315314 196020 333254
rect 197360 332784 197412 332790
rect 197358 332752 197360 332761
rect 197412 332752 197414 332761
rect 197358 332687 197414 332696
rect 198016 332450 198044 457943
rect 198096 456816 198148 456822
rect 198096 456758 198148 456764
rect 198108 332586 198136 456758
rect 198096 332580 198148 332586
rect 198096 332522 198148 332528
rect 198004 332444 198056 332450
rect 198004 332386 198056 332392
rect 197912 331288 197964 331294
rect 197912 331230 197964 331236
rect 195980 315308 196032 315314
rect 195980 315250 196032 315256
rect 103888 206304 103940 206310
rect 103940 206252 104236 206258
rect 103888 206246 104236 206252
rect 103900 206230 104236 206246
rect 162492 205896 162544 205902
rect 158332 205834 158668 205850
rect 162196 205844 162492 205850
rect 162196 205838 162544 205844
rect 158332 205828 158680 205834
rect 158332 205822 158628 205828
rect 162196 205822 162532 205838
rect 158628 205770 158680 205776
rect 154580 205760 154632 205766
rect 142876 205698 143212 205714
rect 154468 205708 154580 205714
rect 154468 205702 154632 205708
rect 28908 205692 28960 205698
rect 142876 205692 143224 205698
rect 142876 205686 143172 205692
rect 28908 205634 28960 205640
rect 154468 205686 154620 205702
rect 143172 205634 143224 205640
rect 23032 205278 23092 205306
rect 26620 205278 26956 205306
rect 23032 204338 23060 205278
rect 23020 204332 23072 204338
rect 23020 204274 23072 204280
rect 22928 204264 22980 204270
rect 22928 204206 22980 204212
rect 22834 203552 22890 203561
rect 22834 203487 22890 203496
rect 22376 202904 22428 202910
rect 22374 202872 22376 202881
rect 22428 202872 22430 202881
rect 22374 202807 22430 202816
rect 22744 202836 22796 202842
rect 22744 202778 22796 202784
rect 22192 202632 22244 202638
rect 22192 202574 22244 202580
rect 22756 202094 22784 202778
rect 22744 202088 22796 202094
rect 22744 202030 22796 202036
rect 21916 74452 21968 74458
rect 21916 74394 21968 74400
rect 22756 74254 22784 202030
rect 22744 74248 22796 74254
rect 22744 74190 22796 74196
rect 22848 74186 22876 203487
rect 22836 74180 22888 74186
rect 22836 74122 22888 74128
rect 22940 74118 22968 204206
rect 26620 204105 26648 205278
rect 26606 204096 26662 204105
rect 26606 204031 26662 204040
rect 28920 203794 28948 205634
rect 30484 205278 30820 205306
rect 34532 205278 34684 205306
rect 38212 205278 38548 205306
rect 42076 205278 42412 205306
rect 45940 205278 46276 205306
rect 49804 205278 50140 205306
rect 53852 205278 54004 205306
rect 57532 205278 57868 205306
rect 61396 205278 61732 205306
rect 65260 205278 65596 205306
rect 69124 205278 69460 205306
rect 73172 205278 73324 205306
rect 76852 205278 77188 205306
rect 80716 205278 81052 205306
rect 84580 205278 84916 205306
rect 88444 205278 88780 205306
rect 92644 205278 92980 205306
rect 30484 204270 30512 205278
rect 30472 204264 30524 204270
rect 30472 204206 30524 204212
rect 34532 204066 34560 205278
rect 30472 204060 30524 204066
rect 30472 204002 30524 204008
rect 34520 204060 34572 204066
rect 34520 204002 34572 204008
rect 34612 204060 34664 204066
rect 34612 204002 34664 204008
rect 28908 203788 28960 203794
rect 28908 203730 28960 203736
rect 30484 203561 30512 204002
rect 34624 203794 34652 204002
rect 38212 203794 38240 205278
rect 34612 203788 34664 203794
rect 34612 203730 34664 203736
rect 34704 203788 34756 203794
rect 34704 203730 34756 203736
rect 38200 203788 38252 203794
rect 38200 203730 38252 203736
rect 30470 203552 30526 203561
rect 30470 203487 30526 203496
rect 23756 202768 23808 202774
rect 23756 202710 23808 202716
rect 23768 202570 23796 202710
rect 23756 202564 23808 202570
rect 23756 202506 23808 202512
rect 34716 202094 34744 203730
rect 42076 202910 42104 205278
rect 39028 202904 39080 202910
rect 39028 202846 39080 202852
rect 42064 202904 42116 202910
rect 42064 202846 42116 202852
rect 39040 202638 39068 202846
rect 45940 202706 45968 205278
rect 49804 202774 49832 205278
rect 53852 202842 53880 205278
rect 53840 202836 53892 202842
rect 53840 202778 53892 202784
rect 49792 202768 49844 202774
rect 57532 202745 57560 205278
rect 61396 203930 61424 205278
rect 65260 203998 65288 205278
rect 65248 203992 65300 203998
rect 65248 203934 65300 203940
rect 61384 203924 61436 203930
rect 61384 203866 61436 203872
rect 69124 202881 69152 205278
rect 73172 204134 73200 205278
rect 76852 204202 76880 205278
rect 76840 204196 76892 204202
rect 76840 204138 76892 204144
rect 73160 204128 73212 204134
rect 73160 204070 73212 204076
rect 80716 204066 80744 205278
rect 80704 204060 80756 204066
rect 80704 204002 80756 204008
rect 84580 203862 84608 205278
rect 88444 204241 88472 205278
rect 92952 204270 92980 205278
rect 96172 205278 96508 205306
rect 99392 205278 100372 205306
rect 107672 205278 108100 205306
rect 111964 205278 112300 205306
rect 96172 204270 96200 205278
rect 92940 204264 92992 204270
rect 88430 204232 88486 204241
rect 92940 204206 92992 204212
rect 95884 204264 95936 204270
rect 95884 204206 95936 204212
rect 96160 204264 96212 204270
rect 96160 204206 96212 204212
rect 88430 204167 88486 204176
rect 84568 203856 84620 203862
rect 84568 203798 84620 203804
rect 69110 202872 69166 202881
rect 69110 202807 69166 202816
rect 49792 202710 49844 202716
rect 57518 202736 57574 202745
rect 45928 202700 45980 202706
rect 57518 202671 57574 202680
rect 45928 202642 45980 202648
rect 39028 202632 39080 202638
rect 39028 202574 39080 202580
rect 34704 202088 34756 202094
rect 34704 202030 34756 202036
rect 95896 186998 95924 204206
rect 99392 199442 99420 205278
rect 107672 200122 107700 205278
rect 112272 203998 112300 205278
rect 115768 205278 115828 205306
rect 118712 205278 119692 205306
rect 123556 205278 123892 205306
rect 127420 205278 127756 205306
rect 115768 204241 115796 205278
rect 115754 204232 115810 204241
rect 115754 204167 115810 204176
rect 112260 203992 112312 203998
rect 112260 203934 112312 203940
rect 107660 200116 107712 200122
rect 107660 200058 107712 200064
rect 99380 199436 99432 199442
rect 99380 199378 99432 199384
rect 118712 189038 118740 205278
rect 123864 204202 123892 205278
rect 123852 204196 123904 204202
rect 123852 204138 123904 204144
rect 127728 203726 127756 205278
rect 131132 205278 131284 205306
rect 135088 205278 135148 205306
rect 139012 205278 139348 205306
rect 146740 205278 147076 205306
rect 150604 205278 150940 205306
rect 166060 205278 166396 205306
rect 169924 205278 170260 205306
rect 127716 203720 127768 203726
rect 127716 203662 127768 203668
rect 118700 189032 118752 189038
rect 118700 188974 118752 188980
rect 131132 188358 131160 205278
rect 135088 201550 135116 205278
rect 139320 203658 139348 205278
rect 147048 204338 147076 205278
rect 147036 204332 147088 204338
rect 147036 204274 147088 204280
rect 150912 204134 150940 205278
rect 150900 204128 150952 204134
rect 150900 204070 150952 204076
rect 139308 203652 139360 203658
rect 139308 203594 139360 203600
rect 166368 202842 166396 205278
rect 166356 202836 166408 202842
rect 166356 202778 166408 202784
rect 170232 202774 170260 205278
rect 173728 205278 173788 205306
rect 177652 205278 177988 205306
rect 181516 205278 181852 205306
rect 185380 205278 185716 205306
rect 189244 205278 189580 205306
rect 173728 204066 173756 205278
rect 177960 204270 177988 205278
rect 177948 204264 178000 204270
rect 177948 204206 178000 204212
rect 179880 204264 179932 204270
rect 179880 204206 179932 204212
rect 173716 204060 173768 204066
rect 173716 204002 173768 204008
rect 179892 203561 179920 204206
rect 181824 203862 181852 205278
rect 183466 204368 183522 204377
rect 183466 204303 183522 204312
rect 183480 204066 183508 204303
rect 183468 204060 183520 204066
rect 183468 204002 183520 204008
rect 181812 203856 181864 203862
rect 181812 203798 181864 203804
rect 179878 203552 179934 203561
rect 179878 203487 179934 203496
rect 185688 203250 185716 205278
rect 187884 203856 187936 203862
rect 187884 203798 187936 203804
rect 185676 203244 185728 203250
rect 185676 203186 185728 203192
rect 170220 202768 170272 202774
rect 170220 202710 170272 202716
rect 187896 202706 187924 203798
rect 189552 203590 189580 205278
rect 193048 205278 193108 205306
rect 195992 205278 196972 205306
rect 193048 204134 193076 205278
rect 193036 204128 193088 204134
rect 193036 204070 193088 204076
rect 195888 204128 195940 204134
rect 195888 204070 195940 204076
rect 195900 203969 195928 204070
rect 195886 203960 195942 203969
rect 195886 203895 195942 203904
rect 189540 203584 189592 203590
rect 189540 203526 189592 203532
rect 188804 203244 188856 203250
rect 188804 203186 188856 203192
rect 187884 202700 187936 202706
rect 187884 202642 187936 202648
rect 188816 202162 188844 203186
rect 188804 202156 188856 202162
rect 188804 202098 188856 202104
rect 135076 201544 135128 201550
rect 135076 201486 135128 201492
rect 131120 188352 131172 188358
rect 131120 188294 131172 188300
rect 195992 187066 196020 205278
rect 197360 204332 197412 204338
rect 197360 204274 197412 204280
rect 197372 204202 197400 204274
rect 197360 204196 197412 204202
rect 197360 204138 197412 204144
rect 197820 204196 197872 204202
rect 197820 204138 197872 204144
rect 197832 203017 197860 204138
rect 197818 203008 197874 203017
rect 197818 202943 197874 202952
rect 197924 202842 197952 331230
rect 198016 204377 198044 332386
rect 198108 331294 198136 332522
rect 198200 332314 198228 460799
rect 198752 458046 198780 585822
rect 198832 583296 198884 583302
rect 198832 583238 198884 583244
rect 198844 458182 198872 583238
rect 198936 460902 198964 585958
rect 199384 583024 199436 583030
rect 199384 582966 199436 582972
rect 199396 462398 199424 582966
rect 199016 462392 199068 462398
rect 199016 462334 199068 462340
rect 199384 462392 199436 462398
rect 199384 462334 199436 462340
rect 199028 460970 199056 462334
rect 199016 460964 199068 460970
rect 199016 460906 199068 460912
rect 198924 460896 198976 460902
rect 198924 460838 198976 460844
rect 198832 458176 198884 458182
rect 198832 458118 198884 458124
rect 198740 458040 198792 458046
rect 198740 457982 198792 457988
rect 198752 451274 198780 457982
rect 198844 456822 198872 458118
rect 198832 456816 198884 456822
rect 198832 456758 198884 456764
rect 198752 451246 198872 451274
rect 198844 332518 198872 451246
rect 198832 332512 198884 332518
rect 198832 332454 198884 332460
rect 198188 332308 198240 332314
rect 198188 332250 198240 332256
rect 198096 331288 198148 331294
rect 198096 331230 198148 331236
rect 198200 316034 198228 332250
rect 198108 316006 198228 316034
rect 198002 204368 198058 204377
rect 198002 204303 198058 204312
rect 197912 202836 197964 202842
rect 197912 202778 197964 202784
rect 197360 202700 197412 202706
rect 197360 202642 197412 202648
rect 197372 202230 197400 202642
rect 197360 202224 197412 202230
rect 197360 202166 197412 202172
rect 195980 187060 196032 187066
rect 195980 187002 196032 187008
rect 95884 186992 95936 186998
rect 95884 186934 95936 186940
rect 88432 78056 88484 78062
rect 191840 78056 191892 78062
rect 88484 78004 89024 78010
rect 88432 77998 89024 78004
rect 88444 77982 89024 77998
rect 184952 77994 185716 78010
rect 191840 77998 191892 78004
rect 192944 78056 192996 78062
rect 192996 78004 193108 78010
rect 192944 77998 193108 78004
rect 23032 77302 23092 77330
rect 26620 77302 26956 77330
rect 30820 77302 31064 77330
rect 34684 77302 35204 77330
rect 23032 75478 23060 77302
rect 26620 75721 26648 77302
rect 26606 75712 26662 75721
rect 26606 75647 26662 75656
rect 23020 75472 23072 75478
rect 23020 75414 23072 75420
rect 31036 74118 31064 77302
rect 35176 74186 35204 77302
rect 38120 77302 38548 77330
rect 42076 77302 42412 77330
rect 46216 77302 46276 77330
rect 50140 77302 50384 77330
rect 54004 77302 54524 77330
rect 38120 74254 38148 77302
rect 42076 74322 42104 77302
rect 46216 74390 46244 77302
rect 50356 75546 50384 77302
rect 50344 75540 50396 75546
rect 50344 75482 50396 75488
rect 50356 75177 50384 75482
rect 50342 75168 50398 75177
rect 50342 75103 50398 75112
rect 54496 74458 54524 77302
rect 57256 77302 57868 77330
rect 61396 77302 61732 77330
rect 65352 77302 65596 77330
rect 69460 77302 69612 77330
rect 57256 74497 57284 77302
rect 61396 75614 61424 77302
rect 65352 75682 65380 77302
rect 69584 75750 69612 77302
rect 73310 77058 73338 77316
rect 76852 77302 77188 77330
rect 81052 77302 81296 77330
rect 73310 77030 73384 77058
rect 73356 75818 73384 77030
rect 76852 75886 76880 77302
rect 76840 75880 76892 75886
rect 81268 75857 81296 77302
rect 84902 77058 84930 77316
rect 84902 77030 84976 77058
rect 76840 75822 76892 75828
rect 81254 75848 81310 75857
rect 73344 75812 73396 75818
rect 73344 75754 73396 75760
rect 69572 75744 69624 75750
rect 69572 75686 69624 75692
rect 65340 75676 65392 75682
rect 65340 75618 65392 75624
rect 61384 75608 61436 75614
rect 61384 75550 61436 75556
rect 57242 74488 57298 74497
rect 54484 74452 54536 74458
rect 57242 74423 57298 74432
rect 54484 74394 54536 74400
rect 46204 74384 46256 74390
rect 46204 74326 46256 74332
rect 42064 74316 42116 74322
rect 42064 74258 42116 74264
rect 38108 74248 38160 74254
rect 38108 74190 38160 74196
rect 35164 74180 35216 74186
rect 35164 74122 35216 74128
rect 22928 74112 22980 74118
rect 22928 74054 22980 74060
rect 31024 74112 31076 74118
rect 31024 74054 31076 74060
rect 31036 65550 31064 74054
rect 31024 65544 31076 65550
rect 31024 65486 31076 65492
rect 35176 62830 35204 74122
rect 38120 72486 38148 74190
rect 38108 72480 38160 72486
rect 38108 72422 38160 72428
rect 42076 62898 42104 74258
rect 46216 65618 46244 74326
rect 54496 66910 54524 74394
rect 54484 66904 54536 66910
rect 54484 66846 54536 66852
rect 46204 65612 46256 65618
rect 46204 65554 46256 65560
rect 57256 64326 57284 74423
rect 57244 64320 57296 64326
rect 57244 64262 57296 64268
rect 61396 64190 61424 75550
rect 65352 74534 65380 75618
rect 69584 75206 69612 75686
rect 69572 75200 69624 75206
rect 69572 75142 69624 75148
rect 65352 74506 65564 74534
rect 65536 64258 65564 74506
rect 73356 73846 73384 75754
rect 73344 73840 73396 73846
rect 73344 73782 73396 73788
rect 76852 69698 76880 75822
rect 81254 75783 81310 75792
rect 81268 71058 81296 75783
rect 84948 74526 84976 77030
rect 84936 74520 84988 74526
rect 84936 74462 84988 74468
rect 81256 71052 81308 71058
rect 81256 70994 81308 71000
rect 76840 69692 76892 69698
rect 76840 69634 76892 69640
rect 84948 68338 84976 74462
rect 88996 71126 89024 77982
rect 103980 77988 104032 77994
rect 103980 77930 104032 77936
rect 184952 77988 185728 77994
rect 184952 77982 185676 77988
rect 96448 77438 96508 77466
rect 92644 77302 92980 77330
rect 92952 75886 92980 77302
rect 96448 75886 96476 77438
rect 103992 77330 104020 77930
rect 100358 77110 100386 77316
rect 103992 77302 104480 77330
rect 108100 77302 108344 77330
rect 111964 77302 112300 77330
rect 99380 77104 99432 77110
rect 99380 77046 99432 77052
rect 100346 77104 100398 77110
rect 100346 77046 100398 77052
rect 99392 76022 99420 77046
rect 99380 76016 99432 76022
rect 99380 75958 99432 75964
rect 92940 75880 92992 75886
rect 92940 75822 92992 75828
rect 96436 75880 96488 75886
rect 96436 75822 96488 75828
rect 96448 75342 96476 75822
rect 96436 75336 96488 75342
rect 96436 75278 96488 75284
rect 88984 71120 89036 71126
rect 88984 71062 89036 71068
rect 84936 68332 84988 68338
rect 84936 68274 84988 68280
rect 65524 64252 65576 64258
rect 65524 64194 65576 64200
rect 61384 64184 61436 64190
rect 61384 64126 61436 64132
rect 99392 63034 99420 75958
rect 104452 72554 104480 77302
rect 108316 75954 108344 77302
rect 108304 75948 108356 75954
rect 108304 75890 108356 75896
rect 104440 72548 104492 72554
rect 104440 72490 104492 72496
rect 108316 68406 108344 75890
rect 112272 75274 112300 77302
rect 114572 77302 115828 77330
rect 119692 77302 119936 77330
rect 112444 75336 112496 75342
rect 112444 75278 112496 75284
rect 112260 75268 112312 75274
rect 112260 75210 112312 75216
rect 108304 68400 108356 68406
rect 108304 68342 108356 68348
rect 112456 67046 112484 75278
rect 112444 67040 112496 67046
rect 112444 66982 112496 66988
rect 99380 63028 99432 63034
rect 99380 62970 99432 62976
rect 42064 62892 42116 62898
rect 42064 62834 42116 62840
rect 35164 62824 35216 62830
rect 35164 62766 35216 62772
rect 57060 62076 57112 62082
rect 57060 62018 57112 62024
rect 57072 61577 57100 62018
rect 57058 61568 57114 61577
rect 57058 61503 57114 61512
rect 114572 60722 114600 77302
rect 119908 73166 119936 77302
rect 122852 77302 123556 77330
rect 127420 77302 127664 77330
rect 131284 77302 131528 77330
rect 122104 75200 122156 75206
rect 122104 75142 122156 75148
rect 119896 73160 119948 73166
rect 119896 73102 119948 73108
rect 122116 66978 122144 75142
rect 122104 66972 122156 66978
rect 122104 66914 122156 66920
rect 114560 60716 114612 60722
rect 114560 60658 114612 60664
rect 122852 60654 122880 77302
rect 127636 70378 127664 77302
rect 131500 71738 131528 77302
rect 135134 77058 135162 77316
rect 139012 77302 139348 77330
rect 135134 77030 135208 77058
rect 131488 71732 131540 71738
rect 131488 71674 131540 71680
rect 127624 70372 127676 70378
rect 127624 70314 127676 70320
rect 135180 69018 135208 77030
rect 139216 75268 139268 75274
rect 139216 75210 139268 75216
rect 139228 74526 139256 75210
rect 139320 75206 139348 77302
rect 142172 77302 142876 77330
rect 146740 77302 147076 77330
rect 150604 77302 150940 77330
rect 139308 75200 139360 75206
rect 139308 75142 139360 75148
rect 139216 74520 139268 74526
rect 139216 74462 139268 74468
rect 135168 69012 135220 69018
rect 135168 68954 135220 68960
rect 142172 66230 142200 77302
rect 147048 75274 147076 77302
rect 150912 75886 150940 77302
rect 153212 77302 154468 77330
rect 158332 77302 158668 77330
rect 150900 75880 150952 75886
rect 150900 75822 150952 75828
rect 147036 75268 147088 75274
rect 147036 75210 147088 75216
rect 142160 66224 142212 66230
rect 142160 66166 142212 66172
rect 122840 60648 122892 60654
rect 122840 60590 122892 60596
rect 103058 59664 103114 59673
rect 103058 59599 103114 59608
rect 102782 58576 102838 58585
rect 102782 58511 102838 58520
rect 102598 56672 102654 56681
rect 102598 56607 102654 56616
rect 57520 56568 57572 56574
rect 57520 56510 57572 56516
rect 57532 56409 57560 56510
rect 57518 56400 57574 56409
rect 57518 56335 57574 56344
rect 102230 54224 102286 54233
rect 102230 54159 102286 54168
rect 102138 53544 102194 53553
rect 102138 53479 102194 53488
rect 102152 52698 102180 53479
rect 102140 52692 102192 52698
rect 102140 52634 102192 52640
rect 102138 52592 102194 52601
rect 102138 52527 102140 52536
rect 102192 52527 102194 52536
rect 102140 52498 102192 52504
rect 57060 52420 57112 52426
rect 57060 52362 57112 52368
rect 57072 51785 57100 52362
rect 57058 51776 57114 51785
rect 57058 51711 57114 51720
rect 102244 48210 102272 54159
rect 102612 49706 102640 56607
rect 102796 51066 102824 58511
rect 102966 55584 103022 55593
rect 102966 55519 103022 55528
rect 102784 51060 102836 51066
rect 102784 51002 102836 51008
rect 102600 49700 102652 49706
rect 102600 49642 102652 49648
rect 102980 48278 103008 55519
rect 103072 52426 103100 59599
rect 153212 57934 153240 77302
rect 158640 75818 158668 77302
rect 161492 77302 162196 77330
rect 166060 77302 166304 77330
rect 169924 77302 170168 77330
rect 158628 75812 158680 75818
rect 158628 75754 158680 75760
rect 156604 75268 156656 75274
rect 156604 75210 156656 75216
rect 156616 63510 156644 75210
rect 156604 63504 156656 63510
rect 156604 63446 156656 63452
rect 153200 57928 153252 57934
rect 153200 57870 153252 57876
rect 161492 57866 161520 77302
rect 166276 68950 166304 77302
rect 170140 70310 170168 77302
rect 173774 77058 173802 77316
rect 177652 77302 177988 77330
rect 173774 77030 173848 77058
rect 173820 73098 173848 77030
rect 177960 75750 177988 77302
rect 180812 77302 181516 77330
rect 177948 75744 178000 75750
rect 177948 75686 178000 75692
rect 173808 73092 173860 73098
rect 173808 73034 173860 73040
rect 170128 70304 170180 70310
rect 170128 70246 170180 70252
rect 166264 68944 166316 68950
rect 166264 68886 166316 68892
rect 180812 59362 180840 77302
rect 180800 59356 180852 59362
rect 180800 59298 180852 59304
rect 184952 58750 184980 77982
rect 185676 77930 185728 77936
rect 189244 77302 189580 77330
rect 189552 75410 189580 77302
rect 189540 75404 189592 75410
rect 189540 75346 189592 75352
rect 191852 60042 191880 77998
rect 192956 77982 193108 77998
rect 196544 77302 196972 77330
rect 196544 64874 196572 77302
rect 197360 68944 197412 68950
rect 197360 68886 197412 68892
rect 197372 68542 197400 68886
rect 197924 68542 197952 202778
rect 198016 73098 198044 204303
rect 198108 202298 198136 316006
rect 198740 314696 198792 314702
rect 198740 314638 198792 314644
rect 198752 204134 198780 314638
rect 198740 204128 198792 204134
rect 198740 204070 198792 204076
rect 198844 202774 198872 332454
rect 198936 332382 198964 460838
rect 199016 456816 199068 456822
rect 199016 456758 199068 456764
rect 198924 332376 198976 332382
rect 198924 332318 198976 332324
rect 198936 203561 198964 332318
rect 199028 315926 199056 456758
rect 199936 332648 199988 332654
rect 199936 332590 199988 332596
rect 199016 315920 199068 315926
rect 199016 315862 199068 315868
rect 199028 314702 199056 315862
rect 199016 314696 199068 314702
rect 199016 314638 199068 314644
rect 199948 204270 199976 332590
rect 199936 204264 199988 204270
rect 199936 204206 199988 204212
rect 199016 204128 199068 204134
rect 199016 204070 199068 204076
rect 198922 203552 198978 203561
rect 198922 203487 198978 203496
rect 198832 202768 198884 202774
rect 198832 202710 198884 202716
rect 198096 202292 198148 202298
rect 198096 202234 198148 202240
rect 198096 202156 198148 202162
rect 198096 202098 198148 202104
rect 198108 77994 198136 202098
rect 198648 201476 198700 201482
rect 198648 201418 198700 201424
rect 198660 201362 198688 201418
rect 198738 201376 198794 201385
rect 198660 201334 198738 201362
rect 198738 201311 198794 201320
rect 198096 77988 198148 77994
rect 198096 77930 198148 77936
rect 198004 73092 198056 73098
rect 198004 73034 198056 73040
rect 198016 72622 198044 73034
rect 198004 72616 198056 72622
rect 198004 72558 198056 72564
rect 198752 69018 198780 201311
rect 198844 70310 198872 202710
rect 198936 75750 198964 203487
rect 199028 75886 199056 204070
rect 199016 75880 199068 75886
rect 199016 75822 199068 75828
rect 198924 75744 198976 75750
rect 198924 75686 198976 75692
rect 198936 74050 198964 75686
rect 199028 75342 199056 75822
rect 199016 75336 199068 75342
rect 199016 75278 199068 75284
rect 198924 74044 198976 74050
rect 198924 73986 198976 73992
rect 198832 70304 198884 70310
rect 198832 70246 198884 70252
rect 199384 70304 199436 70310
rect 199384 70246 199436 70252
rect 199396 69834 199424 70246
rect 199384 69828 199436 69834
rect 199384 69770 199436 69776
rect 198740 69012 198792 69018
rect 198740 68954 198792 68960
rect 198752 68610 198780 68954
rect 198740 68604 198792 68610
rect 198740 68546 198792 68552
rect 197360 68536 197412 68542
rect 197360 68478 197412 68484
rect 197912 68536 197964 68542
rect 197912 68478 197964 68484
rect 195992 64846 196572 64874
rect 191840 60036 191892 60042
rect 191840 59978 191892 59984
rect 184940 58744 184992 58750
rect 184940 58686 184992 58692
rect 195992 58682 196020 64846
rect 197820 63504 197872 63510
rect 197818 63472 197820 63481
rect 197872 63472 197874 63481
rect 197818 63407 197874 63416
rect 197832 62150 197860 63407
rect 197820 62144 197872 62150
rect 197820 62086 197872 62092
rect 195980 58676 196032 58682
rect 195980 58618 196032 58624
rect 161480 57860 161532 57866
rect 161480 57802 161532 57808
rect 104072 52692 104124 52698
rect 104072 52634 104124 52640
rect 103060 52420 103112 52426
rect 103060 52362 103112 52368
rect 103242 51096 103298 51105
rect 103242 51031 103298 51040
rect 103058 49872 103114 49881
rect 103058 49807 103114 49816
rect 102968 48272 103020 48278
rect 102968 48214 103020 48220
rect 102232 48204 102284 48210
rect 102232 48146 102284 48152
rect 102690 47016 102746 47025
rect 102690 46951 102746 46960
rect 57520 46912 57572 46918
rect 57518 46880 57520 46889
rect 57572 46880 57574 46889
rect 57518 46815 57574 46824
rect 102506 44432 102562 44441
rect 102506 44367 102562 44376
rect 102322 43344 102378 43353
rect 102322 43279 102378 43288
rect 57152 42764 57204 42770
rect 57152 42706 57204 42712
rect 57164 42129 57192 42706
rect 57150 42120 57206 42129
rect 57150 42055 57206 42064
rect 102138 41440 102194 41449
rect 102138 41375 102194 41384
rect 102152 38622 102180 41375
rect 102230 40080 102286 40089
rect 102230 40015 102286 40024
rect 102140 38616 102192 38622
rect 102140 38558 102192 38564
rect 102138 37904 102194 37913
rect 102138 37839 102194 37848
rect 57060 37256 57112 37262
rect 57060 37198 57112 37204
rect 57072 36961 57100 37198
rect 57058 36952 57114 36961
rect 57058 36887 57114 36896
rect 102152 35834 102180 37839
rect 102244 37262 102272 40015
rect 102336 39982 102364 43279
rect 102414 42936 102470 42945
rect 102414 42871 102470 42880
rect 102324 39976 102376 39982
rect 102324 39918 102376 39924
rect 102428 38554 102456 42871
rect 102520 40050 102548 44367
rect 102704 42770 102732 46951
rect 102782 45792 102838 45801
rect 102782 45727 102838 45736
rect 102692 42764 102744 42770
rect 102692 42706 102744 42712
rect 102796 41410 102824 45727
rect 103072 44130 103100 49807
rect 103256 45558 103284 51031
rect 103426 48784 103482 48793
rect 103426 48719 103482 48728
rect 103244 45552 103296 45558
rect 103244 45494 103296 45500
rect 103060 44124 103112 44130
rect 103060 44066 103112 44072
rect 103440 44062 103468 48719
rect 104084 46918 104112 52634
rect 196164 52556 196216 52562
rect 196164 52498 196216 52504
rect 195980 52420 196032 52426
rect 195980 52362 196032 52368
rect 195992 51377 196020 52362
rect 195978 51368 196034 51377
rect 195978 51303 196034 51312
rect 195980 51060 196032 51066
rect 195980 51002 196032 51008
rect 195992 50969 196020 51002
rect 195978 50960 196034 50969
rect 195978 50895 196034 50904
rect 195980 49700 196032 49706
rect 195980 49642 196032 49648
rect 195992 49473 196020 49642
rect 195978 49464 196034 49473
rect 195978 49399 196034 49408
rect 195980 48272 196032 48278
rect 195978 48240 195980 48249
rect 196032 48240 196034 48249
rect 195978 48175 196034 48184
rect 196072 48204 196124 48210
rect 196072 48146 196124 48152
rect 196084 47705 196112 48146
rect 196070 47696 196126 47705
rect 196070 47631 196126 47640
rect 104072 46912 104124 46918
rect 195980 46912 196032 46918
rect 104072 46854 104124 46860
rect 195978 46880 195980 46889
rect 196032 46880 196034 46889
rect 195978 46815 196034 46824
rect 196176 46209 196204 52498
rect 196162 46200 196218 46209
rect 196162 46135 196218 46144
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 195992 45257 196020 45494
rect 195978 45248 196034 45257
rect 195978 45183 196034 45192
rect 195980 44124 196032 44130
rect 195980 44066 196032 44072
rect 103428 44056 103480 44062
rect 195992 44033 196020 44066
rect 196072 44056 196124 44062
rect 103428 43998 103480 44004
rect 195978 44024 196034 44033
rect 196072 43998 196124 44004
rect 195978 43959 196034 43968
rect 196084 43625 196112 43998
rect 196070 43616 196126 43625
rect 196070 43551 196126 43560
rect 195980 42764 196032 42770
rect 195980 42706 196032 42712
rect 195992 41585 196020 42706
rect 195978 41576 196034 41585
rect 195978 41511 196034 41520
rect 102784 41404 102836 41410
rect 102784 41346 102836 41352
rect 195980 41404 196032 41410
rect 195980 41346 196032 41352
rect 195992 41177 196020 41346
rect 195978 41168 196034 41177
rect 195978 41103 196034 41112
rect 102508 40044 102560 40050
rect 102508 39986 102560 39992
rect 195980 40044 196032 40050
rect 195980 39986 196032 39992
rect 195992 39953 196020 39986
rect 196072 39976 196124 39982
rect 195978 39944 196034 39953
rect 196072 39918 196124 39924
rect 195978 39879 196034 39888
rect 196084 39545 196112 39918
rect 196070 39536 196126 39545
rect 196070 39471 196126 39480
rect 102874 38992 102930 39001
rect 102874 38927 102930 38936
rect 102416 38548 102468 38554
rect 102416 38490 102468 38496
rect 102598 37360 102654 37369
rect 102598 37295 102654 37304
rect 102232 37256 102284 37262
rect 102232 37198 102284 37204
rect 102140 35828 102192 35834
rect 102140 35770 102192 35776
rect 102138 34640 102194 34649
rect 102138 34575 102194 34584
rect 102152 33114 102180 34575
rect 102612 34474 102640 37295
rect 102782 36136 102838 36145
rect 102782 36071 102838 36080
rect 102600 34468 102652 34474
rect 102600 34410 102652 34416
rect 102796 34406 102824 36071
rect 102888 35902 102916 38927
rect 196072 38616 196124 38622
rect 196072 38558 196124 38564
rect 195980 38548 196032 38554
rect 195980 38490 196032 38496
rect 195992 38457 196020 38490
rect 195978 38448 196034 38457
rect 195978 38383 196034 38392
rect 196084 38049 196112 38558
rect 196070 38040 196126 38049
rect 196070 37975 196126 37984
rect 195980 37256 196032 37262
rect 195980 37198 196032 37204
rect 195992 37097 196020 37198
rect 195978 37088 196034 37097
rect 195978 37023 196034 37032
rect 102876 35896 102928 35902
rect 195980 35896 196032 35902
rect 102876 35838 102928 35844
rect 195978 35864 195980 35873
rect 196032 35864 196034 35873
rect 195978 35799 196034 35808
rect 196072 35828 196124 35834
rect 196072 35770 196124 35776
rect 196084 35465 196112 35770
rect 196070 35456 196126 35465
rect 196070 35391 196126 35400
rect 195980 34468 196032 34474
rect 195980 34410 196032 34416
rect 102784 34400 102836 34406
rect 195992 34377 196020 34410
rect 196072 34400 196124 34406
rect 102784 34342 102836 34348
rect 195978 34368 196034 34377
rect 196072 34342 196124 34348
rect 195978 34303 196034 34312
rect 196084 33833 196112 34342
rect 196070 33824 196126 33833
rect 196070 33759 196126 33768
rect 102322 33552 102378 33561
rect 102322 33487 102378 33496
rect 102140 33108 102192 33114
rect 102140 33050 102192 33056
rect 102138 32464 102194 32473
rect 102138 32399 102194 32408
rect 60004 31816 60056 31822
rect 60004 31758 60056 31764
rect 57612 31748 57664 31754
rect 57612 31690 57664 31696
rect 57624 31657 57652 31690
rect 57610 31648 57666 31657
rect 57610 31583 57666 31592
rect 57244 27600 57296 27606
rect 57244 27542 57296 27548
rect 57256 27169 57284 27542
rect 57242 27160 57298 27169
rect 57242 27095 57298 27104
rect 60016 24274 60044 31758
rect 102152 31686 102180 32399
rect 102230 31784 102286 31793
rect 102336 31754 102364 33487
rect 195980 33108 196032 33114
rect 195980 33050 196032 33056
rect 195992 33017 196020 33050
rect 195978 33008 196034 33017
rect 195978 32943 196034 32952
rect 102230 31719 102286 31728
rect 102324 31748 102376 31754
rect 102140 31680 102192 31686
rect 102140 31622 102192 31628
rect 102138 30560 102194 30569
rect 102138 30495 102194 30504
rect 102152 30258 102180 30495
rect 102244 30326 102272 31719
rect 102324 31690 102376 31696
rect 195980 31748 196032 31754
rect 195980 31690 196032 31696
rect 195992 31657 196020 31690
rect 196072 31680 196124 31686
rect 195978 31648 196034 31657
rect 196072 31622 196124 31628
rect 195978 31583 196034 31592
rect 196084 31249 196112 31622
rect 196070 31240 196126 31249
rect 196070 31175 196126 31184
rect 102232 30320 102284 30326
rect 195980 30320 196032 30326
rect 102232 30262 102284 30268
rect 195978 30288 195980 30297
rect 196032 30288 196034 30297
rect 102140 30252 102192 30258
rect 195978 30223 196034 30232
rect 196072 30252 196124 30258
rect 102140 30194 102192 30200
rect 196072 30194 196124 30200
rect 196084 29753 196112 30194
rect 196070 29744 196126 29753
rect 196070 29679 196126 29688
rect 102138 29336 102194 29345
rect 102138 29271 102194 29280
rect 102152 28966 102180 29271
rect 102140 28960 102192 28966
rect 195980 28960 196032 28966
rect 102140 28902 102192 28908
rect 195978 28928 195980 28937
rect 196032 28928 196034 28937
rect 195978 28863 196034 28872
rect 102138 28520 102194 28529
rect 102138 28455 102194 28464
rect 102152 28286 102180 28455
rect 102140 28280 102192 28286
rect 102140 28222 102192 28228
rect 195980 28280 196032 28286
rect 195980 28222 196032 28228
rect 195992 28121 196020 28222
rect 195978 28112 196034 28121
rect 195978 28047 196034 28056
rect 102138 27704 102194 27713
rect 102138 27639 102194 27648
rect 102152 27606 102180 27639
rect 102140 27600 102192 27606
rect 102140 27542 102192 27548
rect 195980 27600 196032 27606
rect 195980 27542 196032 27548
rect 195992 27305 196020 27542
rect 195978 27296 196034 27305
rect 195978 27231 196034 27240
rect 102782 26344 102838 26353
rect 102782 26279 102838 26288
rect 102796 26246 102824 26279
rect 102784 26240 102836 26246
rect 195980 26240 196032 26246
rect 102784 26182 102836 26188
rect 195978 26208 195980 26217
rect 196032 26208 196034 26217
rect 195978 26143 196034 26152
rect 60004 24268 60056 24274
rect 60004 24210 60056 24216
rect 62316 22098 62344 24140
rect 66272 24126 66746 24154
rect 62304 22092 62356 22098
rect 62304 22034 62356 22040
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 3424 10328 3476 10334
rect 3424 10270 3476 10276
rect 3436 6497 3464 10270
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 66272 3466 66300 24126
rect 71148 17270 71176 24140
rect 74552 24126 75578 24154
rect 78692 24126 79994 24154
rect 84212 24126 84410 24154
rect 71136 17264 71188 17270
rect 71136 17206 71188 17212
rect 74552 15910 74580 24126
rect 74540 15904 74592 15910
rect 74540 15846 74592 15852
rect 78692 6186 78720 24126
rect 84212 8974 84240 24126
rect 88812 21554 88840 24140
rect 92492 24126 93242 24154
rect 96632 24126 97658 24154
rect 88984 23520 89036 23526
rect 88984 23462 89036 23468
rect 88996 22098 89024 23462
rect 88984 22092 89036 22098
rect 88984 22034 89036 22040
rect 88800 21548 88852 21554
rect 88800 21490 88852 21496
rect 84200 8968 84252 8974
rect 84200 8910 84252 8916
rect 78680 6180 78732 6186
rect 78680 6122 78732 6128
rect 92492 4826 92520 24126
rect 96632 4894 96660 24126
rect 200040 22098 200068 699790
rect 218072 586401 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700330 413692 703520
rect 462332 701010 462360 703520
rect 478524 702434 478552 703520
rect 477880 702406 478552 702434
rect 462320 701004 462372 701010
rect 462320 700946 462372 700952
rect 463608 701004 463660 701010
rect 463608 700946 463660 700952
rect 463620 700330 463648 700946
rect 302240 700324 302292 700330
rect 302240 700266 302292 700272
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 463608 700324 463660 700330
rect 463608 700266 463660 700272
rect 302252 596174 302280 700266
rect 302252 596146 302648 596174
rect 302620 588690 302648 596146
rect 302620 588662 303094 588690
rect 306944 586401 306972 587316
rect 218058 586392 218114 586401
rect 218058 586327 218114 586336
rect 306930 586392 306986 586401
rect 306930 586327 306986 586336
rect 310808 586226 310836 587316
rect 200212 586220 200264 586226
rect 200212 586162 200264 586168
rect 301780 586220 301832 586226
rect 301780 586162 301832 586168
rect 310796 586220 310848 586226
rect 310796 586162 310848 586168
rect 200120 583092 200172 583098
rect 200120 583034 200172 583040
rect 200132 444378 200160 583034
rect 200224 459513 200252 586162
rect 200304 586152 200356 586158
rect 200304 586094 200356 586100
rect 200316 460737 200344 586094
rect 258722 585712 258778 585721
rect 258722 585647 258778 585656
rect 201592 583364 201644 583370
rect 201592 583306 201644 583312
rect 201500 583228 201552 583234
rect 201500 583170 201552 583176
rect 200396 583160 200448 583166
rect 200396 583102 200448 583108
rect 200408 461038 200436 583102
rect 201512 461106 201540 583170
rect 201604 461174 201632 583306
rect 201776 572416 201828 572422
rect 201776 572358 201828 572364
rect 201684 572348 201736 572354
rect 201684 572290 201736 572296
rect 201592 461168 201644 461174
rect 201592 461110 201644 461116
rect 201500 461100 201552 461106
rect 201500 461042 201552 461048
rect 200396 461032 200448 461038
rect 200396 460974 200448 460980
rect 200408 460934 200436 460974
rect 200408 460906 200620 460934
rect 200302 460728 200358 460737
rect 200302 460663 200358 460672
rect 200316 459649 200344 460663
rect 200302 459640 200358 459649
rect 200302 459575 200358 459584
rect 200210 459504 200266 459513
rect 200210 459439 200266 459448
rect 200486 459504 200542 459513
rect 200486 459439 200542 459448
rect 200396 458992 200448 458998
rect 200396 458934 200448 458940
rect 200120 444372 200172 444378
rect 200120 444314 200172 444320
rect 200408 335354 200436 458934
rect 200316 335326 200436 335354
rect 200316 332858 200344 335326
rect 200500 335306 200528 459439
rect 200488 335300 200540 335306
rect 200488 335242 200540 335248
rect 200592 335186 200620 460906
rect 200670 459640 200726 459649
rect 200670 459575 200726 459584
rect 200408 335158 200620 335186
rect 200304 332852 200356 332858
rect 200304 332794 200356 332800
rect 200212 332240 200264 332246
rect 200212 332182 200264 332188
rect 200120 205760 200172 205766
rect 200120 205702 200172 205708
rect 200132 57934 200160 205702
rect 200224 202162 200252 332182
rect 200316 205766 200344 332794
rect 200408 332722 200436 335158
rect 200580 335096 200632 335102
rect 200580 335038 200632 335044
rect 200396 332716 200448 332722
rect 200396 332658 200448 332664
rect 200592 332178 200620 335038
rect 200684 332246 200712 459575
rect 200672 332240 200724 332246
rect 200672 332182 200724 332188
rect 200580 332172 200632 332178
rect 200580 332114 200632 332120
rect 200396 330608 200448 330614
rect 200396 330550 200448 330556
rect 200304 205760 200356 205766
rect 200304 205702 200356 205708
rect 200408 204202 200436 330550
rect 200486 316024 200542 316033
rect 200486 315959 200542 315968
rect 200500 315382 200528 315959
rect 200488 315376 200540 315382
rect 200488 315318 200540 315324
rect 200396 204196 200448 204202
rect 200396 204138 200448 204144
rect 200500 203998 200528 315318
rect 200304 203992 200356 203998
rect 200488 203992 200540 203998
rect 200304 203934 200356 203940
rect 200394 203960 200450 203969
rect 200212 202156 200264 202162
rect 200212 202098 200264 202104
rect 200316 74526 200344 203934
rect 200592 203969 200620 332114
rect 201512 330614 201540 461042
rect 201604 332926 201632 461110
rect 201696 458998 201724 572290
rect 201788 480254 201816 572358
rect 202972 572280 203024 572286
rect 202972 572222 203024 572228
rect 202880 572212 202932 572218
rect 202880 572154 202932 572160
rect 201788 480226 201908 480254
rect 201880 459338 201908 480226
rect 201868 459332 201920 459338
rect 201868 459274 201920 459280
rect 201684 458992 201736 458998
rect 201684 458934 201736 458940
rect 201776 444372 201828 444378
rect 201776 444314 201828 444320
rect 201684 332988 201736 332994
rect 201684 332930 201736 332936
rect 201592 332920 201644 332926
rect 201592 332862 201644 332868
rect 201500 330608 201552 330614
rect 201500 330550 201552 330556
rect 201696 209774 201724 332930
rect 201788 331242 201816 444314
rect 201880 332994 201908 459274
rect 202892 458930 202920 572154
rect 202984 459474 203012 572222
rect 203064 572144 203116 572150
rect 203064 572086 203116 572092
rect 203076 460934 203104 572086
rect 245660 572008 245712 572014
rect 245660 571950 245712 571956
rect 247040 572008 247092 572014
rect 247040 571950 247092 571956
rect 204260 462392 204312 462398
rect 204260 462334 204312 462340
rect 203076 460906 203288 460934
rect 203260 459542 203288 460906
rect 203248 459536 203300 459542
rect 203248 459478 203300 459484
rect 202972 459468 203024 459474
rect 202972 459410 203024 459416
rect 202880 458924 202932 458930
rect 202880 458866 202932 458872
rect 201868 332988 201920 332994
rect 201868 332930 201920 332936
rect 201960 332920 202012 332926
rect 201960 332862 202012 332868
rect 201788 331214 201908 331242
rect 201880 331158 201908 331214
rect 201868 331152 201920 331158
rect 201868 331094 201920 331100
rect 201512 209746 201724 209774
rect 201512 205902 201540 209746
rect 201500 205896 201552 205902
rect 201500 205838 201552 205844
rect 200488 203934 200540 203940
rect 200578 203960 200634 203969
rect 200394 203895 200450 203904
rect 200578 203895 200634 203904
rect 200408 78062 200436 203895
rect 200764 203720 200816 203726
rect 200764 203662 200816 203668
rect 200488 202224 200540 202230
rect 200488 202166 200540 202172
rect 200396 78056 200448 78062
rect 200396 77998 200448 78004
rect 200304 74520 200356 74526
rect 200304 74462 200356 74468
rect 200500 59362 200528 202166
rect 200776 70378 200804 203662
rect 201408 74520 201460 74526
rect 201408 74462 201460 74468
rect 201420 73982 201448 74462
rect 201408 73976 201460 73982
rect 201408 73918 201460 73924
rect 200764 70372 200816 70378
rect 200764 70314 200816 70320
rect 201408 70372 201460 70378
rect 201408 70314 201460 70320
rect 201420 69766 201448 70314
rect 201408 69760 201460 69766
rect 201408 69702 201460 69708
rect 200488 59356 200540 59362
rect 200488 59298 200540 59304
rect 201408 59356 201460 59362
rect 201408 59298 201460 59304
rect 201420 58818 201448 59298
rect 201408 58812 201460 58818
rect 201408 58754 201460 58760
rect 200120 57928 200172 57934
rect 200120 57870 200172 57876
rect 201408 57928 201460 57934
rect 201408 57870 201460 57876
rect 201420 57390 201448 57870
rect 201512 57866 201540 205838
rect 201776 205828 201828 205834
rect 201776 205770 201828 205776
rect 201592 205692 201644 205698
rect 201592 205634 201644 205640
rect 201604 66230 201632 205634
rect 201788 75818 201816 205770
rect 201880 203726 201908 331094
rect 201972 205834 202000 332862
rect 202052 332716 202104 332722
rect 202052 332658 202104 332664
rect 201960 205828 202012 205834
rect 201960 205770 202012 205776
rect 202064 205698 202092 332658
rect 202984 329798 203012 459410
rect 203064 330540 203116 330546
rect 203064 330482 203116 330488
rect 202972 329792 203024 329798
rect 202972 329734 203024 329740
rect 202972 314696 203024 314702
rect 202972 314638 203024 314644
rect 202052 205692 202104 205698
rect 202052 205634 202104 205640
rect 202880 204332 202932 204338
rect 202880 204274 202932 204280
rect 201868 203720 201920 203726
rect 201868 203662 201920 203668
rect 202144 188352 202196 188358
rect 202144 188294 202196 188300
rect 201776 75812 201828 75818
rect 201776 75754 201828 75760
rect 202156 71738 202184 188294
rect 202788 75812 202840 75818
rect 202788 75754 202840 75760
rect 202800 75274 202828 75754
rect 202788 75268 202840 75274
rect 202788 75210 202840 75216
rect 202144 71732 202196 71738
rect 202144 71674 202196 71680
rect 202788 71732 202840 71738
rect 202788 71674 202840 71680
rect 202800 71262 202828 71674
rect 202788 71256 202840 71262
rect 202788 71198 202840 71204
rect 201592 66224 201644 66230
rect 201592 66166 201644 66172
rect 202788 66224 202840 66230
rect 202788 66166 202840 66172
rect 202800 65754 202828 66166
rect 202788 65748 202840 65754
rect 202788 65690 202840 65696
rect 202892 60654 202920 204274
rect 202984 204241 203012 314638
rect 202970 204232 203026 204241
rect 202970 204167 203026 204176
rect 202984 60722 203012 204167
rect 203076 189038 203104 330482
rect 203156 329792 203208 329798
rect 203156 329734 203208 329740
rect 203064 189032 203116 189038
rect 203064 188974 203116 188980
rect 203076 73166 203104 188974
rect 203168 188358 203196 329734
rect 203260 315994 203288 459478
rect 204272 332586 204300 462334
rect 244280 458856 244332 458862
rect 244280 458798 244332 458804
rect 204352 443760 204404 443766
rect 204352 443702 204404 443708
rect 204260 332580 204312 332586
rect 204260 332522 204312 332528
rect 204364 330546 204392 443702
rect 233882 331936 233938 331945
rect 233882 331871 233938 331880
rect 204352 330540 204404 330546
rect 204352 330482 204404 330488
rect 203248 315988 203300 315994
rect 203248 315930 203300 315936
rect 203260 314702 203288 315930
rect 203248 314696 203300 314702
rect 203248 314638 203300 314644
rect 203156 188352 203208 188358
rect 203156 188294 203208 188300
rect 229744 75404 229796 75410
rect 229744 75346 229796 75352
rect 227720 73976 227772 73982
rect 227720 73918 227772 73924
rect 212632 73908 212684 73914
rect 212632 73850 212684 73856
rect 203064 73160 203116 73166
rect 203064 73102 203116 73108
rect 203076 72690 203104 73102
rect 203064 72684 203116 72690
rect 203064 72626 203116 72632
rect 203064 71188 203116 71194
rect 203064 71130 203116 71136
rect 202972 60716 203024 60722
rect 202972 60658 203024 60664
rect 202880 60648 202932 60654
rect 202880 60590 202932 60596
rect 201500 57860 201552 57866
rect 201500 57802 201552 57808
rect 202788 57860 202840 57866
rect 202788 57802 202840 57808
rect 201408 57384 201460 57390
rect 201408 57326 201460 57332
rect 202800 57254 202828 57802
rect 202788 57248 202840 57254
rect 202788 57190 202840 57196
rect 203076 54740 203104 71130
rect 209320 63572 209372 63578
rect 209320 63514 209372 63520
rect 207664 61600 207716 61606
rect 207664 61542 207716 61548
rect 204076 60716 204128 60722
rect 204076 60658 204128 60664
rect 204088 60110 204116 60658
rect 204168 60648 204220 60654
rect 204168 60590 204220 60596
rect 204180 60178 204208 60590
rect 206008 60240 206060 60246
rect 206008 60182 206060 60188
rect 204168 60172 204220 60178
rect 204168 60114 204220 60120
rect 204076 60104 204128 60110
rect 204076 60046 204128 60052
rect 204352 60036 204404 60042
rect 204352 59978 204404 59984
rect 204364 54754 204392 59978
rect 206020 54754 206048 60182
rect 207676 54754 207704 61542
rect 209332 54754 209360 63514
rect 211160 61532 211212 61538
rect 211160 61474 211212 61480
rect 211172 54754 211200 61474
rect 212644 54754 212672 73850
rect 224224 72548 224276 72554
rect 224224 72490 224276 72496
rect 220912 65680 220964 65686
rect 220912 65622 220964 65628
rect 219440 62960 219492 62966
rect 219440 62902 219492 62908
rect 214288 61464 214340 61470
rect 214288 61406 214340 61412
rect 214300 54754 214328 61406
rect 217600 61396 217652 61402
rect 217600 61338 217652 61344
rect 215944 60036 215996 60042
rect 215944 59978 215996 59984
rect 215956 54754 215984 59978
rect 217612 54754 217640 61338
rect 219452 54754 219480 62902
rect 220924 54754 220952 65622
rect 222568 63028 222620 63034
rect 222568 62970 222620 62976
rect 222580 54754 222608 62970
rect 224236 54754 224264 72490
rect 225880 68400 225932 68406
rect 225880 68342 225932 68348
rect 225892 54754 225920 68342
rect 227732 54754 227760 73918
rect 229756 60110 229784 75346
rect 230848 72684 230900 72690
rect 230848 72626 230900 72632
rect 229192 60104 229244 60110
rect 229192 60046 229244 60052
rect 229744 60104 229796 60110
rect 229744 60046 229796 60052
rect 229204 54754 229232 60046
rect 230860 54754 230888 72626
rect 233896 68474 233924 331871
rect 241520 316736 241572 316742
rect 241520 316678 241572 316684
rect 240140 203652 240192 203658
rect 240140 203594 240192 203600
rect 238760 75200 238812 75206
rect 238760 75142 238812 75148
rect 238772 74534 238800 75142
rect 240152 74534 240180 203594
rect 241532 74534 241560 316678
rect 238772 74506 239168 74534
rect 240152 74506 240824 74534
rect 241532 74506 242480 74534
rect 236000 71256 236052 71262
rect 236000 71198 236052 71204
rect 234160 69760 234212 69766
rect 234160 69702 234212 69708
rect 233884 68468 233936 68474
rect 233884 68410 233936 68416
rect 232504 60172 232556 60178
rect 232504 60114 232556 60120
rect 232516 54754 232544 60114
rect 234172 54754 234200 69702
rect 236012 54754 236040 71198
rect 237472 68604 237524 68610
rect 237472 68546 237524 68552
rect 237484 54754 237512 68546
rect 239140 54754 239168 74506
rect 240796 54754 240824 74506
rect 242452 54754 242480 74506
rect 244292 54754 244320 458798
rect 245672 74534 245700 571950
rect 247052 74534 247080 571950
rect 258078 331800 258134 331809
rect 258078 331735 258134 331744
rect 249800 318096 249852 318102
rect 249800 318038 249852 318044
rect 249812 74534 249840 318038
rect 252560 189780 252612 189786
rect 252560 189722 252612 189728
rect 245672 74506 245792 74534
rect 247052 74506 247448 74534
rect 249812 74506 250760 74534
rect 245764 54754 245792 74506
rect 247420 54754 247448 74506
rect 249064 60172 249116 60178
rect 249064 60114 249116 60120
rect 249076 54754 249104 60114
rect 250732 54754 250760 74506
rect 252572 54754 252600 189722
rect 256700 186992 256752 186998
rect 256700 186934 256752 186940
rect 255964 75336 256016 75342
rect 255964 75278 256016 75284
rect 254032 72548 254084 72554
rect 254032 72490 254084 72496
rect 254044 54754 254072 72490
rect 255976 67046 256004 75278
rect 256712 74534 256740 186934
rect 258092 74534 258120 331735
rect 256712 74506 257384 74534
rect 258092 74506 258672 74534
rect 255688 67040 255740 67046
rect 255688 66982 255740 66988
rect 255964 67040 256016 67046
rect 255964 66982 256016 66988
rect 255700 54754 255728 66982
rect 257356 54754 257384 74506
rect 258644 55214 258672 74506
rect 258736 57934 258764 585647
rect 300676 583432 300728 583438
rect 300676 583374 300728 583380
rect 299296 583364 299348 583370
rect 299296 583306 299348 583312
rect 297824 583092 297876 583098
rect 297824 583034 297876 583040
rect 263600 570648 263652 570654
rect 263600 570590 263652 570596
rect 260840 443692 260892 443698
rect 260840 443634 260892 443640
rect 258724 57928 258776 57934
rect 258724 57870 258776 57876
rect 258644 55186 259040 55214
rect 259012 54754 259040 55186
rect 260852 54754 260880 443634
rect 263612 74534 263640 570590
rect 297836 459406 297864 583034
rect 298008 583024 298060 583030
rect 298008 582966 298060 582972
rect 297916 580372 297968 580378
rect 297916 580314 297968 580320
rect 297928 460970 297956 580314
rect 297916 460964 297968 460970
rect 297916 460906 297968 460912
rect 297824 459400 297876 459406
rect 297824 459342 297876 459348
rect 283654 458960 283710 458969
rect 283654 458895 283710 458904
rect 283564 458856 283616 458862
rect 283564 458798 283616 458804
rect 264980 445052 265032 445058
rect 264980 444994 265032 445000
rect 264992 74534 265020 444994
rect 266358 331800 266414 331809
rect 266358 331735 266414 331744
rect 266372 74534 266400 331735
rect 269120 203652 269172 203658
rect 269120 203594 269172 203600
rect 263612 74506 264008 74534
rect 264992 74506 265664 74534
rect 266372 74506 267320 74534
rect 262680 57928 262732 57934
rect 262680 57870 262732 57876
rect 204364 54726 204746 54754
rect 206020 54726 206402 54754
rect 207676 54726 208058 54754
rect 209332 54726 209714 54754
rect 211172 54726 211370 54754
rect 212644 54726 213026 54754
rect 214300 54726 214682 54754
rect 215956 54726 216338 54754
rect 217612 54726 217994 54754
rect 219452 54726 219650 54754
rect 220924 54726 221306 54754
rect 222580 54726 222962 54754
rect 224236 54726 224618 54754
rect 225892 54726 226274 54754
rect 227732 54726 227930 54754
rect 229204 54726 229586 54754
rect 230860 54726 231242 54754
rect 232516 54726 232898 54754
rect 234172 54726 234554 54754
rect 236012 54726 236210 54754
rect 237484 54726 237866 54754
rect 239140 54726 239522 54754
rect 240796 54726 241178 54754
rect 242452 54726 242834 54754
rect 244292 54726 244490 54754
rect 245764 54726 246146 54754
rect 247420 54726 247802 54754
rect 249076 54726 249458 54754
rect 250732 54726 251114 54754
rect 252572 54726 252770 54754
rect 254044 54726 254426 54754
rect 255700 54726 256082 54754
rect 257356 54726 257738 54754
rect 259012 54726 259394 54754
rect 260852 54726 261050 54754
rect 262692 54740 262720 57870
rect 263980 54754 264008 74506
rect 265636 54754 265664 74506
rect 267292 54754 267320 74506
rect 269132 54754 269160 203594
rect 278780 75200 278832 75206
rect 278780 75142 278832 75148
rect 271880 74656 271932 74662
rect 271880 74598 271932 74604
rect 271892 74534 271920 74598
rect 274640 74588 274692 74594
rect 274640 74534 274692 74536
rect 278792 74534 278820 75142
rect 271892 74506 272288 74534
rect 274640 74530 275600 74534
rect 274652 74506 275600 74530
rect 278792 74506 278912 74534
rect 270592 71256 270644 71262
rect 270592 71198 270644 71204
rect 270604 54754 270632 71198
rect 272260 54754 272288 74506
rect 274272 57656 274324 57662
rect 274272 57598 274324 57604
rect 263980 54726 264362 54754
rect 265636 54726 266018 54754
rect 267292 54726 267674 54754
rect 269132 54726 269330 54754
rect 270604 54726 270986 54754
rect 272260 54726 272642 54754
rect 274284 54740 274312 57598
rect 275572 54754 275600 74506
rect 277584 57588 277636 57594
rect 277584 57530 277636 57536
rect 275572 54726 275954 54754
rect 277596 54740 277624 57530
rect 278884 54754 278912 74506
rect 282184 65748 282236 65754
rect 282184 65690 282236 65696
rect 280896 57316 280948 57322
rect 280896 57258 280948 57264
rect 278884 54726 279266 54754
rect 280908 54740 280936 57258
rect 282196 54754 282224 65690
rect 283576 60178 283604 458798
rect 283668 60178 283696 458895
rect 283838 458824 283894 458833
rect 283838 458759 283894 458768
rect 283852 76566 283880 458759
rect 297836 335354 297864 459342
rect 297744 335326 297864 335354
rect 297744 332790 297772 335326
rect 297732 332784 297784 332790
rect 297732 332726 297784 332732
rect 296628 204468 296680 204474
rect 296628 204410 296680 204416
rect 296536 200184 296588 200190
rect 296536 200126 296588 200132
rect 283840 76560 283892 76566
rect 283840 76502 283892 76508
rect 288440 75268 288492 75274
rect 288440 75210 288492 75216
rect 288452 74534 288480 75210
rect 288452 74506 288848 74534
rect 285680 67040 285732 67046
rect 285680 66982 285732 66988
rect 283840 62144 283892 62150
rect 283840 62086 283892 62092
rect 283564 60172 283616 60178
rect 283564 60114 283616 60120
rect 283656 60172 283708 60178
rect 283656 60114 283708 60120
rect 283852 54754 283880 62086
rect 285692 54754 285720 66982
rect 287520 57384 287572 57390
rect 287520 57326 287572 57332
rect 282196 54726 282578 54754
rect 283852 54726 284234 54754
rect 285692 54726 285890 54754
rect 287532 54740 287560 57326
rect 288820 54754 288848 74506
rect 293960 72684 294012 72690
rect 293960 72626 294012 72632
rect 292120 65748 292172 65754
rect 292120 65690 292172 65696
rect 290832 57248 290884 57254
rect 290832 57190 290884 57196
rect 288820 54726 289202 54754
rect 290844 54740 290872 57190
rect 292132 54754 292160 65690
rect 293972 54754 294000 72626
rect 295432 68400 295484 68406
rect 295432 68342 295484 68348
rect 295340 60716 295392 60722
rect 295340 60658 295392 60664
rect 295352 60246 295380 60658
rect 295340 60240 295392 60246
rect 295340 60182 295392 60188
rect 295444 54754 295472 68342
rect 296548 58886 296576 200126
rect 296640 60722 296668 204410
rect 297744 201482 297772 332726
rect 297928 332722 297956 460906
rect 298020 459474 298048 582966
rect 298744 572076 298796 572082
rect 298744 572018 298796 572024
rect 298008 459468 298060 459474
rect 298008 459410 298060 459416
rect 297916 332716 297968 332722
rect 297916 332658 297968 332664
rect 297928 206378 297956 332658
rect 298020 315994 298048 459410
rect 298008 315988 298060 315994
rect 298008 315930 298060 315936
rect 297916 206372 297968 206378
rect 297916 206314 297968 206320
rect 298020 204474 298048 315930
rect 298008 204468 298060 204474
rect 298008 204410 298060 204416
rect 297732 201476 297784 201482
rect 297732 201418 297784 201424
rect 297744 200190 297772 201418
rect 297732 200184 297784 200190
rect 297732 200126 297784 200132
rect 298008 186992 298060 186998
rect 298008 186934 298060 186940
rect 297088 69760 297140 69766
rect 297088 69702 297140 69708
rect 296628 60716 296680 60722
rect 296628 60658 296680 60664
rect 296536 58880 296588 58886
rect 296536 58822 296588 58828
rect 297100 54754 297128 69702
rect 298020 62082 298048 186934
rect 298652 73976 298704 73982
rect 298652 73918 298704 73924
rect 298008 62076 298060 62082
rect 298008 62018 298060 62024
rect 298020 61606 298048 62018
rect 298008 61600 298060 61606
rect 298008 61542 298060 61548
rect 298664 55214 298692 73918
rect 298756 57361 298784 572018
rect 299308 459338 299336 583306
rect 300584 583228 300636 583234
rect 300584 583170 300636 583176
rect 300492 583160 300544 583166
rect 300492 583102 300544 583108
rect 299388 580304 299440 580310
rect 299388 580246 299440 580252
rect 299296 459332 299348 459338
rect 299296 459274 299348 459280
rect 299308 332926 299336 459274
rect 299400 459134 299428 580246
rect 300400 572076 300452 572082
rect 300400 572018 300452 572024
rect 300308 462324 300360 462330
rect 300308 462266 300360 462272
rect 300320 461174 300348 462266
rect 300308 461168 300360 461174
rect 300308 461110 300360 461116
rect 299388 459128 299440 459134
rect 299388 459070 299440 459076
rect 299296 332920 299348 332926
rect 299296 332862 299348 332868
rect 299400 315330 299428 459070
rect 300124 332920 300176 332926
rect 300124 332862 300176 332868
rect 299478 315344 299534 315353
rect 298836 315308 298888 315314
rect 298836 315250 298888 315256
rect 299400 315302 299478 315330
rect 298848 57390 298876 315250
rect 299294 314800 299350 314809
rect 299294 314735 299350 314744
rect 299308 187678 299336 314735
rect 299400 314294 299428 315302
rect 299478 315279 299534 315288
rect 299388 314288 299440 314294
rect 299388 314230 299440 314236
rect 300136 204950 300164 332862
rect 300320 332489 300348 461110
rect 300412 460934 300440 572018
rect 300504 462330 300532 583102
rect 300492 462324 300544 462330
rect 300492 462266 300544 462272
rect 300596 462233 300624 583170
rect 300582 462224 300638 462233
rect 300582 462159 300638 462168
rect 300596 461038 300624 462159
rect 300584 461032 300636 461038
rect 300584 460974 300636 460980
rect 300412 460906 300532 460934
rect 300504 459270 300532 460906
rect 300492 459264 300544 459270
rect 300492 459206 300544 459212
rect 300504 332586 300532 459206
rect 300688 459202 300716 583374
rect 300768 583296 300820 583302
rect 300768 583238 300820 583244
rect 300780 461106 300808 583238
rect 300768 461100 300820 461106
rect 300768 461042 300820 461048
rect 300676 459196 300728 459202
rect 300676 459138 300728 459144
rect 300492 332580 300544 332586
rect 300492 332522 300544 332528
rect 300306 332480 300362 332489
rect 300306 332415 300362 332424
rect 300216 314288 300268 314294
rect 300216 314230 300268 314236
rect 300228 206310 300256 314230
rect 300216 206304 300268 206310
rect 300216 206246 300268 206252
rect 300228 205737 300256 206246
rect 300214 205728 300270 205737
rect 300214 205663 300270 205672
rect 299388 204944 299440 204950
rect 299388 204886 299440 204892
rect 300124 204944 300176 204950
rect 300124 204886 300176 204892
rect 299296 187672 299348 187678
rect 299296 187614 299348 187620
rect 299308 64394 299336 187614
rect 299400 71738 299428 204886
rect 300504 204241 300532 332522
rect 300584 315920 300636 315926
rect 300582 315888 300584 315897
rect 300636 315888 300638 315897
rect 300582 315823 300638 315832
rect 300688 315722 300716 459138
rect 300780 315858 300808 461042
rect 301792 460934 301820 586162
rect 314672 586158 314700 587316
rect 301872 586152 301924 586158
rect 301872 586094 301924 586100
rect 314660 586152 314712 586158
rect 314660 586094 314712 586100
rect 301700 460906 301820 460934
rect 301700 459241 301728 460906
rect 301884 459377 301912 586094
rect 318536 586090 318564 587316
rect 302700 586084 302752 586090
rect 302700 586026 302752 586032
rect 318524 586084 318576 586090
rect 318524 586026 318576 586032
rect 302148 586016 302200 586022
rect 302148 585958 302200 585964
rect 301964 585880 302016 585886
rect 301964 585822 302016 585828
rect 301870 459368 301926 459377
rect 301870 459303 301926 459312
rect 301686 459232 301742 459241
rect 301686 459167 301742 459176
rect 301502 458280 301558 458289
rect 301502 458215 301558 458224
rect 301516 332246 301544 458215
rect 301594 457056 301650 457065
rect 301594 456991 301650 457000
rect 301504 332240 301556 332246
rect 301504 332182 301556 332188
rect 301516 331294 301544 332182
rect 301504 331288 301556 331294
rect 301504 331230 301556 331236
rect 300768 315852 300820 315858
rect 300768 315794 300820 315800
rect 300676 315716 300728 315722
rect 300676 315658 300728 315664
rect 300584 314696 300636 314702
rect 300584 314638 300636 314644
rect 300596 204542 300624 314638
rect 300688 204678 300716 315658
rect 300780 314702 300808 315794
rect 301608 315382 301636 456991
rect 301700 331838 301728 459167
rect 301884 458289 301912 459303
rect 301870 458280 301926 458289
rect 301870 458215 301926 458224
rect 301976 458114 302004 585822
rect 302054 585712 302110 585721
rect 302054 585647 302110 585656
rect 302068 458153 302096 585647
rect 302054 458144 302110 458153
rect 301964 458108 302016 458114
rect 302054 458079 302110 458088
rect 301964 458050 302016 458056
rect 301870 456920 301926 456929
rect 301870 456855 301926 456864
rect 301884 332382 301912 456855
rect 301976 332518 302004 458050
rect 302068 457065 302096 458079
rect 302160 457881 302188 585958
rect 302712 459513 302740 586026
rect 322400 586022 322428 587316
rect 322388 586016 322440 586022
rect 322388 585958 322440 585964
rect 326264 585954 326292 587316
rect 302884 585948 302936 585954
rect 302884 585890 302936 585896
rect 326252 585948 326304 585954
rect 326252 585890 326304 585896
rect 302792 585812 302844 585818
rect 302792 585754 302844 585760
rect 302698 459504 302754 459513
rect 302698 459439 302754 459448
rect 302146 457872 302202 457881
rect 302146 457807 302202 457816
rect 302054 457056 302110 457065
rect 302054 456991 302110 457000
rect 302160 456929 302188 457807
rect 302146 456920 302202 456929
rect 302146 456855 302202 456864
rect 302608 456816 302660 456822
rect 302608 456758 302660 456764
rect 301964 332512 302016 332518
rect 301964 332454 302016 332460
rect 301872 332376 301924 332382
rect 301872 332318 301924 332324
rect 301688 331832 301740 331838
rect 301688 331774 301740 331780
rect 301780 331288 301832 331294
rect 301780 331230 301832 331236
rect 301596 315376 301648 315382
rect 301596 315318 301648 315324
rect 300768 314696 300820 314702
rect 300768 314638 300820 314644
rect 300676 204672 300728 204678
rect 300676 204614 300728 204620
rect 300584 204536 300636 204542
rect 300584 204478 300636 204484
rect 300490 204232 300546 204241
rect 300490 204167 300546 204176
rect 300124 203584 300176 203590
rect 300124 203526 300176 203532
rect 299388 71732 299440 71738
rect 299388 71674 299440 71680
rect 300032 64864 300084 64870
rect 300030 64832 300032 64841
rect 300084 64832 300086 64841
rect 300030 64767 300086 64776
rect 299296 64388 299348 64394
rect 299296 64330 299348 64336
rect 300044 63578 300072 64767
rect 300032 63572 300084 63578
rect 300032 63514 300084 63520
rect 300136 57526 300164 203526
rect 300216 187060 300268 187066
rect 300216 187002 300268 187008
rect 300124 57520 300176 57526
rect 300124 57462 300176 57468
rect 300228 57458 300256 187002
rect 300596 75274 300624 204478
rect 300688 75886 300716 204614
rect 300766 204232 300822 204241
rect 300766 204167 300822 204176
rect 300676 75880 300728 75886
rect 300676 75822 300728 75828
rect 300584 75268 300636 75274
rect 300584 75210 300636 75216
rect 300780 69018 300808 204167
rect 301792 203998 301820 331230
rect 301884 204066 301912 332318
rect 301976 204202 302004 332454
rect 302056 332172 302108 332178
rect 302056 332114 302108 332120
rect 302068 331838 302096 332114
rect 302056 331832 302108 331838
rect 302056 331774 302108 331780
rect 301964 204196 302016 204202
rect 301964 204138 302016 204144
rect 301872 204060 301924 204066
rect 301872 204002 301924 204008
rect 301780 203992 301832 203998
rect 301780 203934 301832 203940
rect 301792 78402 301820 203934
rect 301780 78396 301832 78402
rect 301780 78338 301832 78344
rect 301884 78266 301912 204002
rect 301872 78260 301924 78266
rect 301872 78202 301924 78208
rect 301976 78130 302004 204138
rect 302068 203930 302096 331774
rect 302148 315784 302200 315790
rect 302148 315726 302200 315732
rect 302160 315382 302188 315726
rect 302620 315586 302648 456758
rect 302712 332314 302740 459439
rect 302804 458182 302832 585754
rect 302792 458176 302844 458182
rect 302792 458118 302844 458124
rect 302804 456822 302832 458118
rect 302896 458046 302924 585890
rect 330128 585886 330156 587316
rect 330116 585880 330168 585886
rect 330116 585822 330168 585828
rect 333992 585818 334020 587316
rect 333980 585812 334032 585818
rect 333980 585754 334032 585760
rect 337856 583001 337884 587316
rect 341720 583438 341748 587316
rect 345032 587302 345598 587330
rect 341708 583432 341760 583438
rect 341708 583374 341760 583380
rect 337842 582992 337898 583001
rect 337842 582927 337898 582936
rect 345032 572082 345060 587302
rect 349448 585721 349476 587316
rect 349434 585712 349490 585721
rect 349434 585647 349490 585656
rect 353312 583370 353340 587316
rect 353300 583364 353352 583370
rect 353300 583306 353352 583312
rect 357176 583302 357204 587316
rect 357164 583296 357216 583302
rect 357164 583238 357216 583244
rect 361040 583234 361068 587316
rect 361028 583228 361080 583234
rect 361028 583170 361080 583176
rect 364904 583166 364932 587316
rect 364892 583160 364944 583166
rect 364892 583102 364944 583108
rect 368768 583098 368796 587316
rect 372632 586158 372660 587316
rect 376496 586498 376524 587316
rect 373264 586492 373316 586498
rect 373264 586434 373316 586440
rect 376484 586492 376536 586498
rect 376484 586434 376536 586440
rect 373276 586158 373304 586434
rect 372620 586152 372672 586158
rect 372620 586094 372672 586100
rect 373264 586152 373316 586158
rect 373264 586094 373316 586100
rect 368756 583092 368808 583098
rect 368756 583034 368808 583040
rect 345020 572076 345072 572082
rect 345020 572018 345072 572024
rect 373276 570654 373304 586094
rect 380360 583030 380388 587316
rect 380348 583024 380400 583030
rect 380348 582966 380400 582972
rect 384224 580378 384252 587316
rect 384212 580372 384264 580378
rect 384212 580314 384264 580320
rect 388088 580310 388116 587316
rect 391952 583001 391980 587316
rect 391938 582992 391994 583001
rect 391938 582927 391994 582936
rect 395816 580310 395844 587316
rect 399680 580378 399708 587316
rect 403544 583030 403572 587316
rect 407408 583098 407436 587316
rect 411272 583166 411300 587316
rect 415136 583234 415164 587316
rect 418172 587302 419014 587330
rect 415124 583228 415176 583234
rect 415124 583170 415176 583176
rect 411260 583160 411312 583166
rect 411260 583102 411312 583108
rect 407396 583092 407448 583098
rect 407396 583034 407448 583040
rect 403532 583024 403584 583030
rect 403532 582966 403584 582972
rect 399668 580372 399720 580378
rect 399668 580314 399720 580320
rect 388076 580304 388128 580310
rect 388076 580246 388128 580252
rect 395804 580304 395856 580310
rect 395804 580246 395856 580252
rect 418172 572014 418200 587302
rect 422864 583302 422892 587316
rect 426728 583370 426756 587316
rect 430592 585721 430620 587316
rect 433352 587302 434470 587330
rect 437492 587302 438334 587330
rect 430578 585712 430634 585721
rect 430578 585647 430634 585656
rect 426716 583364 426768 583370
rect 426716 583306 426768 583312
rect 422852 583296 422904 583302
rect 422852 583238 422904 583244
rect 433352 572014 433380 587302
rect 437492 572082 437520 587302
rect 442184 583438 442212 587316
rect 446048 585818 446076 587316
rect 449912 585886 449940 587316
rect 453776 585954 453804 587316
rect 457640 586022 457668 587316
rect 461504 586090 461532 587316
rect 465368 586158 465396 587316
rect 465356 586152 465408 586158
rect 465356 586094 465408 586100
rect 461492 586084 461544 586090
rect 461492 586026 461544 586032
rect 457628 586016 457680 586022
rect 457628 585958 457680 585964
rect 453764 585948 453816 585954
rect 453764 585890 453816 585896
rect 449900 585880 449952 585886
rect 469232 585857 469260 587316
rect 449900 585822 449952 585828
rect 469218 585848 469274 585857
rect 446036 585812 446088 585818
rect 469218 585783 469274 585792
rect 446036 585754 446088 585760
rect 473096 585206 473124 587316
rect 473084 585200 473136 585206
rect 476960 585177 476988 587316
rect 477880 586401 477908 702406
rect 485780 700324 485832 700330
rect 485780 700266 485832 700272
rect 477866 586392 477922 586401
rect 477866 586327 477922 586336
rect 479064 586152 479116 586158
rect 479064 586094 479116 586100
rect 478144 586084 478196 586090
rect 478144 586026 478196 586032
rect 477960 585948 478012 585954
rect 477960 585890 478012 585896
rect 477868 585812 477920 585818
rect 477868 585754 477920 585760
rect 473084 585142 473136 585148
rect 476946 585168 477002 585177
rect 476946 585103 477002 585112
rect 442172 583432 442224 583438
rect 442172 583374 442224 583380
rect 437480 572076 437532 572082
rect 437480 572018 437532 572024
rect 418160 572008 418212 572014
rect 418160 571950 418212 571956
rect 433340 572008 433392 572014
rect 433340 571950 433392 571956
rect 373264 570648 373316 570654
rect 373264 570590 373316 570596
rect 392216 462392 392268 462398
rect 391966 462340 392216 462346
rect 391966 462334 392268 462340
rect 391966 462318 392256 462334
rect 303080 461009 303108 461244
rect 303066 461000 303122 461009
rect 303066 460935 303122 460944
rect 306944 460873 306972 461244
rect 306930 460864 306986 460873
rect 306930 460799 306986 460808
rect 310808 459241 310836 461244
rect 314672 459377 314700 461244
rect 318536 459513 318564 461244
rect 318522 459504 318578 459513
rect 318522 459439 318578 459448
rect 314658 459368 314714 459377
rect 314658 459303 314714 459312
rect 310794 459232 310850 459241
rect 310794 459167 310850 459176
rect 302884 458040 302936 458046
rect 302884 457982 302936 457988
rect 302792 456816 302844 456822
rect 302792 456758 302844 456764
rect 302896 451274 302924 457982
rect 322400 457881 322428 461244
rect 326264 458046 326292 461244
rect 330128 458114 330156 461244
rect 333992 458182 334020 461244
rect 333980 458176 334032 458182
rect 333980 458118 334032 458124
rect 330116 458108 330168 458114
rect 330116 458050 330168 458056
rect 326252 458040 326304 458046
rect 337856 458017 337884 461244
rect 341720 459202 341748 461244
rect 345584 459270 345612 461244
rect 345572 459264 345624 459270
rect 345572 459206 345624 459212
rect 341708 459196 341760 459202
rect 341708 459138 341760 459144
rect 349448 458153 349476 461244
rect 353312 459338 353340 461244
rect 357176 461106 357204 461244
rect 357164 461100 357216 461106
rect 357164 461042 357216 461048
rect 361040 461038 361068 461244
rect 364260 461230 364918 461258
rect 364260 461174 364288 461230
rect 364248 461168 364300 461174
rect 364248 461110 364300 461116
rect 361028 461032 361080 461038
rect 361028 460974 361080 460980
rect 368768 459406 368796 461244
rect 372632 459542 372660 461244
rect 376496 459542 376524 461244
rect 372620 459536 372672 459542
rect 372620 459478 372672 459484
rect 373264 459536 373316 459542
rect 373264 459478 373316 459484
rect 376484 459536 376536 459542
rect 376484 459478 376536 459484
rect 368756 459400 368808 459406
rect 368756 459342 368808 459348
rect 353300 459332 353352 459338
rect 353300 459274 353352 459280
rect 349434 458144 349490 458153
rect 349434 458079 349490 458088
rect 326252 457982 326304 457988
rect 337842 458008 337898 458017
rect 337842 457943 337898 457952
rect 322386 457872 322442 457881
rect 322386 457807 322442 457816
rect 302804 451246 302924 451274
rect 302804 332450 302832 451246
rect 373276 445058 373304 459478
rect 380360 459474 380388 461244
rect 384224 460970 384252 461244
rect 384212 460964 384264 460970
rect 384212 460906 384264 460912
rect 380348 459468 380400 459474
rect 380348 459410 380400 459416
rect 388088 459134 388116 461244
rect 388076 459128 388128 459134
rect 388076 459070 388128 459076
rect 395816 458182 395844 461244
rect 395804 458176 395856 458182
rect 395804 458118 395856 458124
rect 399680 458114 399708 461244
rect 403544 459202 403572 461244
rect 407408 459474 407436 461244
rect 407396 459468 407448 459474
rect 407396 459410 407448 459416
rect 411272 459406 411300 461244
rect 415136 459542 415164 461244
rect 415124 459536 415176 459542
rect 415124 459478 415176 459484
rect 418712 459536 418764 459542
rect 418712 459478 418764 459484
rect 411260 459400 411312 459406
rect 411260 459342 411312 459348
rect 403532 459196 403584 459202
rect 403532 459138 403584 459144
rect 399668 458108 399720 458114
rect 399668 458050 399720 458056
rect 418724 458046 418752 459478
rect 419000 458862 419028 461244
rect 418988 458856 419040 458862
rect 418988 458798 419040 458804
rect 418712 458040 418764 458046
rect 418712 457982 418764 457988
rect 422864 457978 422892 461244
rect 422852 457972 422904 457978
rect 422852 457914 422904 457920
rect 426728 457910 426756 461244
rect 430592 459338 430620 461244
rect 430580 459332 430632 459338
rect 430580 459274 430632 459280
rect 434456 458862 434484 461244
rect 438320 459270 438348 461244
rect 442184 460970 442212 461244
rect 446048 461038 446076 461244
rect 449912 461106 449940 461244
rect 453790 461230 453988 461258
rect 453960 461174 453988 461230
rect 453948 461168 454000 461174
rect 453948 461110 454000 461116
rect 449900 461100 449952 461106
rect 449900 461042 449952 461048
rect 446036 461032 446088 461038
rect 446036 460974 446088 460980
rect 442172 460964 442224 460970
rect 442172 460906 442224 460912
rect 457640 459542 457668 461244
rect 461504 460934 461532 461244
rect 461504 460906 461624 460934
rect 461490 459640 461546 459649
rect 461490 459575 461546 459584
rect 461504 459542 461532 459575
rect 461596 459542 461624 460906
rect 465368 459542 465396 461244
rect 457628 459536 457680 459542
rect 457628 459478 457680 459484
rect 461492 459536 461544 459542
rect 461492 459478 461544 459484
rect 461584 459536 461636 459542
rect 461584 459478 461636 459484
rect 463792 459536 463844 459542
rect 463792 459478 463844 459484
rect 465356 459536 465408 459542
rect 465356 459478 465408 459484
rect 438308 459264 438360 459270
rect 438308 459206 438360 459212
rect 434444 458856 434496 458862
rect 463804 458833 463832 459478
rect 469232 458930 469260 461244
rect 473096 460902 473124 461244
rect 473084 460896 473136 460902
rect 473084 460838 473136 460844
rect 469312 459536 469364 459542
rect 469312 459478 469364 459484
rect 469324 458969 469352 459478
rect 469310 458960 469366 458969
rect 469220 458924 469272 458930
rect 469310 458895 469366 458904
rect 469220 458866 469272 458872
rect 434444 458798 434496 458804
rect 463790 458824 463846 458833
rect 463790 458759 463846 458768
rect 476960 458289 476988 461244
rect 477880 461038 477908 585754
rect 477972 461174 478000 585890
rect 478052 585200 478104 585206
rect 478052 585142 478104 585148
rect 477960 461168 478012 461174
rect 477960 461110 478012 461116
rect 477868 461032 477920 461038
rect 477868 460974 477920 460980
rect 476946 458280 477002 458289
rect 476946 458215 477002 458224
rect 426716 457904 426768 457910
rect 426716 457846 426768 457852
rect 373264 445052 373316 445058
rect 373264 444994 373316 445000
rect 442448 334008 442500 334014
rect 442198 333956 442448 333962
rect 442198 333950 442500 333956
rect 442198 333934 442488 333950
rect 302884 332852 302936 332858
rect 302884 332794 302936 332800
rect 302896 332489 302924 332794
rect 303080 332489 303108 333268
rect 306944 332654 306972 333268
rect 306932 332648 306984 332654
rect 306932 332590 306984 332596
rect 302882 332480 302938 332489
rect 302792 332444 302844 332450
rect 302882 332415 302938 332424
rect 303066 332480 303122 332489
rect 303066 332415 303122 332424
rect 302792 332386 302844 332392
rect 302700 332308 302752 332314
rect 302700 332250 302752 332256
rect 302608 315580 302660 315586
rect 302608 315522 302660 315528
rect 302148 315376 302200 315382
rect 302148 315318 302200 315324
rect 302056 203924 302108 203930
rect 302056 203866 302108 203872
rect 301964 78124 302016 78130
rect 301964 78066 302016 78072
rect 302068 77994 302096 203866
rect 302160 187610 302188 315318
rect 302620 314838 302648 315522
rect 302608 314832 302660 314838
rect 302608 314774 302660 314780
rect 302712 204270 302740 332250
rect 302700 204264 302752 204270
rect 302700 204206 302752 204212
rect 302148 187604 302200 187610
rect 302148 187546 302200 187552
rect 302056 77988 302108 77994
rect 302056 77930 302108 77936
rect 300768 69012 300820 69018
rect 300768 68954 300820 68960
rect 302160 67046 302188 187546
rect 302712 78334 302740 204206
rect 302804 204134 302832 332386
rect 310808 332178 310836 333268
rect 314672 332246 314700 333268
rect 318536 332314 318564 333268
rect 322400 332382 322428 333268
rect 326264 332450 326292 333268
rect 330128 332518 330156 333268
rect 330116 332512 330168 332518
rect 330116 332454 330168 332460
rect 326252 332444 326304 332450
rect 326252 332386 326304 332392
rect 322388 332376 322440 332382
rect 322388 332318 322440 332324
rect 318524 332308 318576 332314
rect 318524 332250 318576 332256
rect 314660 332240 314712 332246
rect 314660 332182 314712 332188
rect 310796 332172 310848 332178
rect 310796 332114 310848 332120
rect 303528 315648 303580 315654
rect 303526 315616 303528 315625
rect 303580 315616 303582 315625
rect 333992 315586 334020 333268
rect 336752 333254 337870 333282
rect 340892 333254 341734 333282
rect 336752 315654 336780 333254
rect 340892 315722 340920 333254
rect 345584 332586 345612 333268
rect 349172 333254 349462 333282
rect 345572 332580 345624 332586
rect 345572 332522 345624 332528
rect 349172 315790 349200 333254
rect 350540 332920 350592 332926
rect 350540 332862 350592 332868
rect 350552 332586 350580 332862
rect 353312 332586 353340 333268
rect 356072 333254 357190 333282
rect 360212 333254 361054 333282
rect 350540 332580 350592 332586
rect 350540 332522 350592 332528
rect 353300 332580 353352 332586
rect 353300 332522 353352 332528
rect 356072 315858 356100 333254
rect 360212 315926 360240 333254
rect 361580 332852 361632 332858
rect 361580 332794 361632 332800
rect 361592 332586 361620 332794
rect 364904 332586 364932 333268
rect 368768 332790 368796 333268
rect 368756 332784 368808 332790
rect 368756 332726 368808 332732
rect 372632 332586 372660 333268
rect 376496 332586 376524 333268
rect 379532 333254 380374 333282
rect 361580 332580 361632 332586
rect 361580 332522 361632 332528
rect 364892 332580 364944 332586
rect 364892 332522 364944 332528
rect 372620 332580 372672 332586
rect 372620 332522 372672 332528
rect 376484 332580 376536 332586
rect 376484 332522 376536 332528
rect 372632 331809 372660 332522
rect 372618 331800 372674 331809
rect 372618 331735 372674 331744
rect 379532 315994 379560 333254
rect 384224 332722 384252 333268
rect 387812 333254 388102 333282
rect 384212 332716 384264 332722
rect 384212 332658 384264 332664
rect 379520 315988 379572 315994
rect 379520 315930 379572 315936
rect 360200 315920 360252 315926
rect 360200 315862 360252 315868
rect 356060 315852 356112 315858
rect 356060 315794 356112 315800
rect 349160 315784 349212 315790
rect 349160 315726 349212 315732
rect 340880 315716 340932 315722
rect 340880 315658 340932 315664
rect 336740 315648 336792 315654
rect 336740 315590 336792 315596
rect 303526 315551 303582 315560
rect 333980 315580 334032 315586
rect 333980 315522 334032 315528
rect 387812 315353 387840 333254
rect 391952 315994 391980 333268
rect 395816 332722 395844 333268
rect 395804 332716 395856 332722
rect 395804 332658 395856 332664
rect 399680 331294 399708 333268
rect 403544 331294 403572 333268
rect 399668 331288 399720 331294
rect 399668 331230 399720 331236
rect 400864 331288 400916 331294
rect 400864 331230 400916 331236
rect 403532 331288 403584 331294
rect 403532 331230 403584 331236
rect 405004 331288 405056 331294
rect 405004 331230 405056 331236
rect 391940 315988 391992 315994
rect 391940 315930 391992 315936
rect 400876 315858 400904 331230
rect 405016 315926 405044 331230
rect 407408 329798 407436 333268
rect 407396 329792 407448 329798
rect 407396 329734 407448 329740
rect 411272 329730 411300 333268
rect 415136 331294 415164 333268
rect 418172 333254 419014 333282
rect 422312 333254 422878 333282
rect 426452 333254 426742 333282
rect 415124 331288 415176 331294
rect 415124 331230 415176 331236
rect 411260 329724 411312 329730
rect 411260 329666 411312 329672
rect 418172 318102 418200 333254
rect 418620 331220 418672 331226
rect 418620 331162 418672 331168
rect 418632 329662 418660 331162
rect 418620 329656 418672 329662
rect 418620 329598 418672 329604
rect 418160 318096 418212 318102
rect 418160 318038 418212 318044
rect 405004 315920 405056 315926
rect 405004 315862 405056 315868
rect 400864 315852 400916 315858
rect 400864 315794 400916 315800
rect 422312 315790 422340 333254
rect 422300 315784 422352 315790
rect 422300 315726 422352 315732
rect 426452 315722 426480 333254
rect 430592 332586 430620 333268
rect 433352 333254 434470 333282
rect 438334 333266 438900 333282
rect 438334 333260 438912 333266
rect 438334 333254 438860 333260
rect 433248 332784 433300 332790
rect 433248 332726 433300 332732
rect 433260 332586 433288 332726
rect 430580 332580 430632 332586
rect 430580 332522 430632 332528
rect 433248 332580 433300 332586
rect 433248 332522 433300 332528
rect 426440 315716 426492 315722
rect 426440 315658 426492 315664
rect 433352 315654 433380 333254
rect 438860 333202 438912 333208
rect 446048 332178 446076 333268
rect 449912 332518 449940 333268
rect 449900 332512 449952 332518
rect 449900 332454 449952 332460
rect 453776 332450 453804 333268
rect 453764 332444 453816 332450
rect 453764 332386 453816 332392
rect 457640 332382 457668 333268
rect 457628 332376 457680 332382
rect 457628 332318 457680 332324
rect 461504 332314 461532 333268
rect 461492 332308 461544 332314
rect 461492 332250 461544 332256
rect 465368 332246 465396 333268
rect 465356 332240 465408 332246
rect 465356 332182 465408 332188
rect 446036 332172 446088 332178
rect 446036 332114 446088 332120
rect 469232 331809 469260 333268
rect 473096 332586 473124 333268
rect 473084 332580 473136 332586
rect 473084 332522 473136 332528
rect 469218 331800 469274 331809
rect 469218 331735 469274 331744
rect 476960 331265 476988 333268
rect 477880 332178 477908 460974
rect 477972 332450 478000 461110
rect 478064 460902 478092 585142
rect 478052 460896 478104 460902
rect 478052 460838 478104 460844
rect 478064 332586 478092 460838
rect 478156 458833 478184 586026
rect 478972 586016 479024 586022
rect 478972 585958 479024 585964
rect 478880 583228 478932 583234
rect 478880 583170 478932 583176
rect 478788 462936 478840 462942
rect 478788 462878 478840 462884
rect 478800 462398 478828 462878
rect 478788 462392 478840 462398
rect 478788 462334 478840 462340
rect 478142 458824 478198 458833
rect 478142 458759 478198 458768
rect 478052 332580 478104 332586
rect 478052 332522 478104 332528
rect 477960 332444 478012 332450
rect 477960 332386 478012 332392
rect 477868 332172 477920 332178
rect 477868 332114 477920 332120
rect 477880 331294 477908 332114
rect 477868 331288 477920 331294
rect 476946 331256 477002 331265
rect 477868 331230 477920 331236
rect 476946 331191 477002 331200
rect 477498 329760 477554 329769
rect 477498 329695 477554 329704
rect 477512 329662 477540 329695
rect 477500 329656 477552 329662
rect 477500 329598 477552 329604
rect 476120 315852 476172 315858
rect 476120 315794 476172 315800
rect 433340 315648 433392 315654
rect 433340 315590 433392 315596
rect 476132 315353 476160 315794
rect 387798 315344 387854 315353
rect 387798 315279 387854 315288
rect 476118 315344 476174 315353
rect 476118 315279 476174 315288
rect 302884 314832 302936 314838
rect 302884 314774 302936 314780
rect 302896 204610 302924 314774
rect 477972 229094 478000 332386
rect 478156 332314 478184 458759
rect 478800 456754 478828 462334
rect 478892 458046 478920 583170
rect 478984 459649 479012 585958
rect 478970 459640 479026 459649
rect 478970 459575 479026 459584
rect 478880 458040 478932 458046
rect 478880 457982 478932 457988
rect 478892 456929 478920 457982
rect 478878 456920 478934 456929
rect 478878 456855 478934 456864
rect 478788 456748 478840 456754
rect 478788 456690 478840 456696
rect 478420 333328 478472 333334
rect 478420 333270 478472 333276
rect 478432 332790 478460 333270
rect 478420 332784 478472 332790
rect 478420 332726 478472 332732
rect 478144 332308 478196 332314
rect 478144 332250 478196 332256
rect 477972 229066 478092 229094
rect 442354 206680 442410 206689
rect 442198 206638 442354 206666
rect 442354 206615 442410 206624
rect 476120 206576 476172 206582
rect 476120 206518 476172 206524
rect 313280 206372 313332 206378
rect 313280 206314 313332 206320
rect 302884 204604 302936 204610
rect 302884 204546 302936 204552
rect 302792 204128 302844 204134
rect 302792 204070 302844 204076
rect 302700 78328 302752 78334
rect 302700 78270 302752 78276
rect 302804 78198 302832 204070
rect 302792 78192 302844 78198
rect 302792 78134 302844 78140
rect 302240 68536 302292 68542
rect 302240 68478 302292 68484
rect 302148 67040 302200 67046
rect 302148 66982 302200 66988
rect 300216 57452 300268 57458
rect 300216 57394 300268 57400
rect 298836 57384 298888 57390
rect 298742 57352 298798 57361
rect 298836 57326 298888 57332
rect 298742 57287 298798 57296
rect 300768 57248 300820 57254
rect 300768 57190 300820 57196
rect 298664 55186 298784 55214
rect 298756 54754 298784 55186
rect 292132 54726 292514 54754
rect 293972 54726 294170 54754
rect 295444 54726 295826 54754
rect 297100 54726 297482 54754
rect 298756 54726 299138 54754
rect 300780 54740 300808 57190
rect 302252 54754 302280 68478
rect 302896 67590 302924 204546
rect 303080 204338 303108 205292
rect 306944 204406 306972 205292
rect 306932 204400 306984 204406
rect 306932 204342 306984 204348
rect 303068 204332 303120 204338
rect 303068 204274 303120 204280
rect 310808 203930 310836 205292
rect 313292 203930 313320 206314
rect 387800 206304 387852 206310
rect 387852 206252 388102 206258
rect 387800 206246 388102 206252
rect 387812 206230 388102 206246
rect 438584 205760 438636 205766
rect 391966 205698 392256 205714
rect 438334 205708 438584 205714
rect 476132 205737 476160 206518
rect 438334 205702 438636 205708
rect 476118 205728 476174 205737
rect 391966 205692 392268 205698
rect 391966 205686 392216 205692
rect 438334 205686 438624 205702
rect 476118 205663 476120 205672
rect 392216 205634 392268 205640
rect 476172 205663 476174 205672
rect 476120 205634 476172 205640
rect 476132 205603 476160 205634
rect 314672 203998 314700 205292
rect 318536 204270 318564 205292
rect 318524 204264 318576 204270
rect 318524 204206 318576 204212
rect 322400 204066 322428 205292
rect 326264 204134 326292 205292
rect 330128 204202 330156 205292
rect 333992 204610 334020 205292
rect 333980 204604 334032 204610
rect 333980 204546 334032 204552
rect 337856 204377 337884 205292
rect 341352 205278 341734 205306
rect 341352 204678 341380 205278
rect 341340 204672 341392 204678
rect 341340 204614 341392 204620
rect 337842 204368 337898 204377
rect 337842 204303 337898 204312
rect 330116 204196 330168 204202
rect 330116 204138 330168 204144
rect 326252 204128 326304 204134
rect 345584 204105 345612 205292
rect 349172 205278 349462 205306
rect 326252 204070 326304 204076
rect 345570 204096 345626 204105
rect 322388 204060 322440 204066
rect 345570 204031 345626 204040
rect 322388 204002 322440 204008
rect 314660 203992 314712 203998
rect 314660 203934 314712 203940
rect 310796 203924 310848 203930
rect 310796 203866 310848 203872
rect 312544 203924 312596 203930
rect 312544 203866 312596 203872
rect 313280 203924 313332 203930
rect 313280 203866 313332 203872
rect 312556 186998 312584 203866
rect 349172 187610 349200 205278
rect 349252 204944 349304 204950
rect 349252 204886 349304 204892
rect 349264 204270 349292 204886
rect 353312 204270 353340 205292
rect 357176 204542 357204 205292
rect 360212 205278 361054 205306
rect 357164 204536 357216 204542
rect 357164 204478 357216 204484
rect 349252 204264 349304 204270
rect 349252 204206 349304 204212
rect 353300 204264 353352 204270
rect 353300 204206 353352 204212
rect 360212 187678 360240 205278
rect 364904 204241 364932 205292
rect 364890 204232 364946 204241
rect 364890 204167 364946 204176
rect 368768 201482 368796 205292
rect 372632 204270 372660 205292
rect 376496 204270 376524 205292
rect 380360 204474 380388 205292
rect 380348 204468 380400 204474
rect 380348 204410 380400 204416
rect 372620 204264 372672 204270
rect 372620 204206 372672 204212
rect 376484 204264 376536 204270
rect 376484 204206 376536 204212
rect 372632 203658 372660 204206
rect 384224 203930 384252 205292
rect 384212 203924 384264 203930
rect 384212 203866 384264 203872
rect 372620 203652 372672 203658
rect 372620 203594 372672 203600
rect 395816 201482 395844 205292
rect 399680 202910 399708 205292
rect 403544 204270 403572 205292
rect 407028 204604 407080 204610
rect 407028 204546 407080 204552
rect 407040 204270 407068 204546
rect 403532 204264 403584 204270
rect 403532 204206 403584 204212
rect 407028 204264 407080 204270
rect 407028 204206 407080 204212
rect 407408 202910 407436 205292
rect 411272 204134 411300 205292
rect 415136 204270 415164 205292
rect 418172 205278 419014 205306
rect 415124 204264 415176 204270
rect 415124 204206 415176 204212
rect 411260 204128 411312 204134
rect 411260 204070 411312 204076
rect 413928 204128 413980 204134
rect 413928 204070 413980 204076
rect 399668 202904 399720 202910
rect 399668 202846 399720 202852
rect 407396 202904 407448 202910
rect 407396 202846 407448 202852
rect 410800 202904 410852 202910
rect 410800 202846 410852 202852
rect 368756 201476 368808 201482
rect 368756 201418 368808 201424
rect 395804 201476 395856 201482
rect 395804 201418 395856 201424
rect 410812 201414 410840 202846
rect 410800 201408 410852 201414
rect 410800 201350 410852 201356
rect 413940 201346 413968 204070
rect 413928 201340 413980 201346
rect 413928 201282 413980 201288
rect 418172 189786 418200 205278
rect 418712 204672 418764 204678
rect 418712 204614 418764 204620
rect 418724 204270 418752 204614
rect 422864 204474 422892 205292
rect 426728 204542 426756 205292
rect 426716 204536 426768 204542
rect 426716 204478 426768 204484
rect 422852 204468 422904 204474
rect 422852 204410 422904 204416
rect 418712 204264 418764 204270
rect 430592 204241 430620 205292
rect 434470 205278 434760 205306
rect 434732 204746 434760 205278
rect 434720 204740 434772 204746
rect 434720 204682 434772 204688
rect 418712 204206 418764 204212
rect 430578 204232 430634 204241
rect 430578 204167 430634 204176
rect 446048 204105 446076 205292
rect 446034 204096 446090 204105
rect 446034 204031 446090 204040
rect 449912 203930 449940 205292
rect 453776 204202 453804 205292
rect 453764 204196 453816 204202
rect 453764 204138 453816 204144
rect 457640 204134 457668 205292
rect 457628 204128 457680 204134
rect 457628 204070 457680 204076
rect 461504 204066 461532 205292
rect 461492 204060 461544 204066
rect 461492 204002 461544 204008
rect 465368 203998 465396 205292
rect 465356 203992 465408 203998
rect 465356 203934 465408 203940
rect 449900 203924 449952 203930
rect 449900 203866 449952 203872
rect 469232 203590 469260 205292
rect 473096 203998 473124 205292
rect 475476 204264 475528 204270
rect 475382 204232 475438 204241
rect 475476 204206 475528 204212
rect 475382 204167 475438 204176
rect 473084 203992 473136 203998
rect 475396 203969 475424 204167
rect 475488 204066 475516 204206
rect 476960 204134 476988 205292
rect 477868 204264 477920 204270
rect 477868 204206 477920 204212
rect 477958 204232 478014 204241
rect 476948 204128 477000 204134
rect 476948 204070 477000 204076
rect 475476 204060 475528 204066
rect 475476 204002 475528 204008
rect 476028 203992 476080 203998
rect 473084 203934 473136 203940
rect 475382 203960 475438 203969
rect 476028 203934 476080 203940
rect 475382 203895 475438 203904
rect 476040 203833 476068 203934
rect 476026 203824 476082 203833
rect 476026 203759 476082 203768
rect 469220 203584 469272 203590
rect 469220 203526 469272 203532
rect 477498 202872 477554 202881
rect 477498 202807 477500 202816
rect 477552 202807 477554 202816
rect 477500 202778 477552 202784
rect 418160 189780 418212 189786
rect 418160 189722 418212 189728
rect 360200 187672 360252 187678
rect 360200 187614 360252 187620
rect 349160 187604 349212 187610
rect 349160 187546 349212 187552
rect 312544 186992 312596 186998
rect 312544 186934 312596 186940
rect 314752 78396 314804 78402
rect 314752 78338 314804 78344
rect 307208 78056 307260 78062
rect 306958 78004 307208 78010
rect 306958 77998 307260 78004
rect 306958 77982 307248 77998
rect 310532 77994 310822 78010
rect 310520 77988 310822 77994
rect 310572 77982 310822 77988
rect 311164 77988 311216 77994
rect 310520 77930 310572 77936
rect 311164 77930 311216 77936
rect 303342 77344 303398 77353
rect 303094 77302 303342 77330
rect 303342 77279 303398 77288
rect 307024 74044 307076 74050
rect 307024 73986 307076 73992
rect 305368 72616 305420 72622
rect 305368 72558 305420 72564
rect 303712 69828 303764 69834
rect 303712 69770 303764 69776
rect 302884 67584 302936 67590
rect 302884 67526 302936 67532
rect 303724 54754 303752 69770
rect 305380 54754 305408 72558
rect 307036 54754 307064 73986
rect 308680 58812 308732 58818
rect 308680 58754 308732 58760
rect 308692 54754 308720 58754
rect 310532 57934 310560 77930
rect 311176 77353 311204 77930
rect 311162 77344 311218 77353
rect 314764 77330 314792 78338
rect 317420 78328 317472 78334
rect 317420 78270 317472 78276
rect 318156 78328 318208 78334
rect 318208 78276 318550 78282
rect 318156 78270 318550 78276
rect 316776 78260 316828 78266
rect 316776 78202 316828 78208
rect 314686 77316 314792 77330
rect 311162 77279 311218 77288
rect 314672 77302 314792 77316
rect 311164 74044 311216 74050
rect 311164 73986 311216 73992
rect 310612 58744 310664 58750
rect 310612 58686 310664 58692
rect 310520 57928 310572 57934
rect 310520 57870 310572 57876
rect 310624 54754 310652 58686
rect 311176 57662 311204 73986
rect 314672 57974 314700 77302
rect 316788 75818 316816 78202
rect 316776 75812 316828 75818
rect 316776 75754 316828 75760
rect 316960 75812 317012 75818
rect 316960 75754 317012 75760
rect 314488 57946 314700 57974
rect 312360 57928 312412 57934
rect 312360 57870 312412 57876
rect 311164 57656 311216 57662
rect 311164 57598 311216 57604
rect 302252 54726 302450 54754
rect 303724 54726 304106 54754
rect 305380 54726 305762 54754
rect 307036 54726 307418 54754
rect 308692 54726 309074 54754
rect 310624 54726 310730 54754
rect 312372 54740 312400 57870
rect 314488 54754 314516 57946
rect 315672 56636 315724 56642
rect 315672 56578 315724 56584
rect 314042 54726 314516 54754
rect 315684 54740 315712 56578
rect 316972 54754 317000 75754
rect 317432 56642 317460 78270
rect 318168 78254 318550 78270
rect 318800 78192 318852 78198
rect 430672 78192 430724 78198
rect 393318 78160 393374 78169
rect 318800 78134 318852 78140
rect 318812 75750 318840 78134
rect 329852 78130 330142 78146
rect 329840 78124 330142 78130
rect 329892 78118 330142 78124
rect 329840 78066 329892 78072
rect 322400 75818 322428 77316
rect 326264 75818 326292 77316
rect 322388 75812 322440 75818
rect 322388 75754 322440 75760
rect 326252 75812 326304 75818
rect 326252 75754 326304 75760
rect 318800 75744 318852 75750
rect 318800 75686 318852 75692
rect 317420 56636 317472 56642
rect 317420 56578 317472 56584
rect 318812 54754 318840 75686
rect 322204 75404 322256 75410
rect 322204 75346 322256 75352
rect 322216 67590 322244 75346
rect 327080 75336 327132 75342
rect 327080 75278 327132 75284
rect 327092 69018 327120 75278
rect 329840 71732 329892 71738
rect 329840 71674 329892 71680
rect 327080 69012 327132 69018
rect 327080 68954 327132 68960
rect 322204 67584 322256 67590
rect 322204 67526 322256 67532
rect 322216 64874 322244 67526
rect 321940 64846 322244 64874
rect 320272 63028 320324 63034
rect 320272 62970 320324 62976
rect 320284 54754 320312 62970
rect 321940 54754 321968 64846
rect 323584 59016 323636 59022
rect 323584 58958 323636 58964
rect 323596 54754 323624 58958
rect 325240 58812 325292 58818
rect 325240 58754 325292 58760
rect 325252 54754 325280 58754
rect 327092 54754 327120 68954
rect 328552 67040 328604 67046
rect 328552 66982 328604 66988
rect 328564 54754 328592 66982
rect 329852 55214 329880 71674
rect 329944 63034 329972 78118
rect 430672 78134 430724 78140
rect 393318 78095 393374 78104
rect 394700 78124 394752 78130
rect 390558 78024 390614 78033
rect 390558 77959 390614 77968
rect 336738 77888 336794 77897
rect 336738 77823 336794 77832
rect 337474 77888 337530 77897
rect 389178 77888 389234 77897
rect 337530 77846 337870 77874
rect 337474 77823 337530 77832
rect 389178 77823 389234 77832
rect 333992 75410 334020 77316
rect 333980 75404 334032 75410
rect 333980 75346 334032 75352
rect 331220 75268 331272 75274
rect 331220 75210 331272 75216
rect 331232 74534 331260 75210
rect 331232 74506 331904 74534
rect 330300 72616 330352 72622
rect 330300 72558 330352 72564
rect 330312 71738 330340 72558
rect 330300 71732 330352 71738
rect 330300 71674 330352 71680
rect 329932 63028 329984 63034
rect 329932 62970 329984 62976
rect 329852 55186 330248 55214
rect 330220 54754 330248 55186
rect 331876 54754 331904 74506
rect 333520 64388 333572 64394
rect 333520 64330 333572 64336
rect 332600 64320 332652 64326
rect 332600 64262 332652 64268
rect 332612 57662 332640 64262
rect 332600 57656 332652 57662
rect 332600 57598 332652 57604
rect 333532 54754 333560 64330
rect 335360 62144 335412 62150
rect 335360 62086 335412 62092
rect 335372 54754 335400 62086
rect 336752 59022 336780 77823
rect 340984 77302 341734 77330
rect 340984 75886 341012 77302
rect 340972 75880 341024 75886
rect 340972 75822 341024 75828
rect 336830 75168 336886 75177
rect 336830 75103 336886 75112
rect 336844 63510 336872 75103
rect 340880 72480 340932 72486
rect 340880 72422 340932 72428
rect 338488 65544 338540 65550
rect 338488 65486 338540 65492
rect 336832 63504 336884 63510
rect 336832 63446 336884 63452
rect 336844 62150 336872 63446
rect 336832 62144 336884 62150
rect 336832 62086 336884 62092
rect 336740 59016 336792 59022
rect 336740 58958 336792 58964
rect 336832 58880 336884 58886
rect 336832 58822 336884 58828
rect 336844 54754 336872 58822
rect 338500 54754 338528 65486
rect 340144 62824 340196 62830
rect 340144 62766 340196 62772
rect 340156 54754 340184 62766
rect 340892 55214 340920 72422
rect 340984 58818 341012 75822
rect 345584 75342 345612 77316
rect 349172 77302 349462 77330
rect 345572 75336 345624 75342
rect 345572 75278 345624 75284
rect 349172 67046 349200 77302
rect 353312 72622 353340 77316
rect 357176 75274 357204 77316
rect 360304 77302 361054 77330
rect 364352 77302 364918 77330
rect 368492 77302 368782 77330
rect 357164 75268 357216 75274
rect 357164 75210 357216 75216
rect 356704 73840 356756 73846
rect 356704 73782 356756 73788
rect 353300 72616 353352 72622
rect 353300 72558 353352 72564
rect 349160 67040 349212 67046
rect 349160 66982 349212 66988
rect 355048 66972 355100 66978
rect 355048 66914 355100 66920
rect 348424 66904 348476 66910
rect 348424 66846 348476 66852
rect 345112 65612 345164 65618
rect 345112 65554 345164 65560
rect 343640 62892 343692 62898
rect 343640 62834 343692 62840
rect 341064 62824 341116 62830
rect 341064 62766 341116 62772
rect 340972 58812 341024 58818
rect 340972 58754 341024 58760
rect 341076 57594 341104 62766
rect 341064 57588 341116 57594
rect 341064 57530 341116 57536
rect 340892 55186 341840 55214
rect 341812 54754 341840 55186
rect 343652 54754 343680 62834
rect 345124 54754 345152 65554
rect 346766 58576 346822 58585
rect 346766 58511 346822 58520
rect 346780 54754 346808 58511
rect 348436 54754 348464 66846
rect 353392 64252 353444 64258
rect 353392 64194 353444 64200
rect 351920 64184 351972 64190
rect 351920 64126 351972 64132
rect 350448 57656 350500 57662
rect 350448 57598 350500 57604
rect 316972 54726 317354 54754
rect 318812 54726 319010 54754
rect 320284 54726 320666 54754
rect 321940 54726 322322 54754
rect 323596 54726 323978 54754
rect 325252 54726 325634 54754
rect 327092 54726 327290 54754
rect 328564 54726 328946 54754
rect 330220 54726 330602 54754
rect 331876 54726 332258 54754
rect 333532 54726 333914 54754
rect 335372 54726 335570 54754
rect 336844 54726 337226 54754
rect 338500 54726 338882 54754
rect 340156 54726 340538 54754
rect 341812 54726 342194 54754
rect 343652 54726 343850 54754
rect 345124 54726 345506 54754
rect 346780 54726 347162 54754
rect 348436 54726 348818 54754
rect 350460 54740 350488 57598
rect 351932 54754 351960 64126
rect 353404 54754 353432 64194
rect 355060 54754 355088 66914
rect 356716 54754 356744 73782
rect 360200 71052 360252 71058
rect 360200 70994 360252 71000
rect 358360 69692 358412 69698
rect 358360 69634 358412 69640
rect 358372 54754 358400 69634
rect 360212 54754 360240 70994
rect 360304 64394 360332 77302
rect 363328 71120 363380 71126
rect 363328 71062 363380 71068
rect 361672 68332 361724 68338
rect 361672 68274 361724 68280
rect 360292 64388 360344 64394
rect 360292 64330 360344 64336
rect 361684 54754 361712 68274
rect 363340 54754 363368 71062
rect 364352 63510 364380 77302
rect 364340 63504 364392 63510
rect 364340 63446 364392 63452
rect 364984 60104 365036 60110
rect 364984 60046 365036 60052
rect 364996 54754 365024 60046
rect 368492 58750 368520 77302
rect 369860 76560 369912 76566
rect 369860 76502 369912 76508
rect 369872 74534 369900 76502
rect 372632 75886 372660 77316
rect 372712 77308 372764 77314
rect 372712 77250 372764 77256
rect 372620 75880 372672 75886
rect 372620 75822 372672 75828
rect 369872 74506 369992 74534
rect 368572 68468 368624 68474
rect 368572 68410 368624 68416
rect 368480 58744 368532 58750
rect 368480 58686 368532 58692
rect 367008 57520 367060 57526
rect 367008 57462 367060 57468
rect 351932 54726 352130 54754
rect 353404 54726 353786 54754
rect 355060 54726 355442 54754
rect 356716 54726 357098 54754
rect 358372 54726 358754 54754
rect 360212 54726 360410 54754
rect 361684 54726 362066 54754
rect 363340 54726 363722 54754
rect 364996 54726 365378 54754
rect 367020 54740 367048 57462
rect 368584 54754 368612 68410
rect 369964 54754 369992 74506
rect 372632 71262 372660 75822
rect 372724 74534 372752 77250
rect 376496 75886 376524 77316
rect 379532 77302 380374 77330
rect 383672 77302 384238 77330
rect 387812 77302 388102 77330
rect 376484 75880 376536 75886
rect 376484 75822 376536 75828
rect 375380 75404 375432 75410
rect 375380 75346 375432 75352
rect 373998 75168 374054 75177
rect 373998 75103 374054 75112
rect 374012 74534 374040 75103
rect 372724 74506 373304 74534
rect 374012 74506 374960 74534
rect 372620 71256 372672 71262
rect 372620 71198 372672 71204
rect 371974 57352 372030 57361
rect 371974 57287 372030 57296
rect 368584 54726 368690 54754
rect 369964 54726 370346 54754
rect 371988 54740 372016 57287
rect 373276 54754 373304 74506
rect 374932 54754 374960 74506
rect 375392 72690 375420 75346
rect 376760 75336 376812 75342
rect 376760 75278 376812 75284
rect 375380 72684 375432 72690
rect 375380 72626 375432 72632
rect 376772 54754 376800 75278
rect 378140 75268 378192 75274
rect 378140 75210 378192 75216
rect 378152 74534 378180 75210
rect 378152 74506 378272 74534
rect 378244 54754 378272 74506
rect 379532 60722 379560 77302
rect 383672 62082 383700 77302
rect 387812 64870 387840 77302
rect 389192 74534 389220 77823
rect 390572 74534 390600 77959
rect 391966 77302 392348 77330
rect 392320 74534 392348 77302
rect 389192 74506 389864 74534
rect 390572 74506 391520 74534
rect 392320 74506 392624 74534
rect 387800 64864 387852 64870
rect 387800 64806 387852 64812
rect 383660 62076 383712 62082
rect 383660 62018 383712 62024
rect 379520 60716 379572 60722
rect 379520 60658 379572 60664
rect 386512 60172 386564 60178
rect 386512 60114 386564 60120
rect 379888 60104 379940 60110
rect 379888 60046 379940 60052
rect 379900 54754 379928 60046
rect 381544 58676 381596 58682
rect 381544 58618 381596 58624
rect 381556 54754 381584 58618
rect 383568 57452 383620 57458
rect 383568 57394 383620 57400
rect 373276 54726 373658 54754
rect 374932 54726 375314 54754
rect 376772 54726 376970 54754
rect 378244 54726 378626 54754
rect 379900 54726 380282 54754
rect 381556 54726 381938 54754
rect 383580 54740 383608 57394
rect 385224 57384 385276 57390
rect 385224 57326 385276 57332
rect 385236 54740 385264 57326
rect 386524 54754 386552 60114
rect 388534 57216 388590 57225
rect 388534 57151 388590 57160
rect 386524 54726 386906 54754
rect 388548 54740 388576 57151
rect 389836 54754 389864 74506
rect 391492 54754 391520 74506
rect 392596 74361 392624 74506
rect 392582 74352 392638 74361
rect 392582 74287 392638 74296
rect 392596 61538 392624 74287
rect 392584 61532 392636 61538
rect 392584 61474 392636 61480
rect 393332 54754 393360 78095
rect 394700 78066 394752 78072
rect 394712 74534 394740 78066
rect 430684 77330 430712 78134
rect 394712 74506 394832 74534
rect 394804 54754 394832 74506
rect 395816 74497 395844 77316
rect 399496 77302 399694 77330
rect 403558 77302 403664 77330
rect 407422 77302 407804 77330
rect 395802 74488 395858 74497
rect 395802 74423 395858 74432
rect 395816 73914 395844 74423
rect 395804 73908 395856 73914
rect 395804 73850 395856 73856
rect 399496 73137 399524 77302
rect 403636 73166 403664 77302
rect 403624 73160 403676 73166
rect 399482 73128 399538 73137
rect 403624 73102 403676 73108
rect 399482 73063 399538 73072
rect 399496 61470 399524 73063
rect 399484 61464 399536 61470
rect 399484 61406 399536 61412
rect 403636 60042 403664 73102
rect 407776 73098 407804 77302
rect 407764 73092 407816 73098
rect 407764 73034 407816 73040
rect 407776 61402 407804 73034
rect 411272 73030 411300 77316
rect 415136 75546 415164 77316
rect 414664 75540 414716 75546
rect 414664 75482 414716 75488
rect 415124 75540 415176 75546
rect 415124 75482 415176 75488
rect 411260 73024 411312 73030
rect 411260 72966 411312 72972
rect 411904 73024 411956 73030
rect 411904 72966 411956 72972
rect 411916 62966 411944 72966
rect 414676 65686 414704 75482
rect 419000 72554 419028 77316
rect 422864 75954 422892 77316
rect 426742 77302 427124 77330
rect 430606 77316 430712 77330
rect 422852 75948 422904 75954
rect 422852 75890 422904 75896
rect 422864 74662 422892 75890
rect 422852 74656 422904 74662
rect 422852 74598 422904 74604
rect 427096 74526 427124 77302
rect 430592 77302 430712 77316
rect 430592 74594 430620 77302
rect 434456 75818 434484 77316
rect 433984 75812 434036 75818
rect 433984 75754 434036 75760
rect 434444 75812 434496 75818
rect 434444 75754 434496 75760
rect 430580 74588 430632 74594
rect 430580 74530 430632 74536
rect 427084 74520 427136 74526
rect 427084 74462 427136 74468
rect 427096 74050 427124 74462
rect 427084 74044 427136 74050
rect 427084 73986 427136 73992
rect 418988 72548 419040 72554
rect 418988 72490 419040 72496
rect 414664 65680 414716 65686
rect 414664 65622 414716 65628
rect 411904 62960 411956 62966
rect 411904 62902 411956 62908
rect 433996 62830 434024 75754
rect 438320 75750 438348 77316
rect 442198 77302 442304 77330
rect 446062 77302 446444 77330
rect 438308 75744 438360 75750
rect 438308 75686 438360 75692
rect 438320 75206 438348 75686
rect 442276 75682 442304 77302
rect 442264 75676 442316 75682
rect 442264 75618 442316 75624
rect 438308 75200 438360 75206
rect 438308 75142 438360 75148
rect 433984 62824 434036 62830
rect 433984 62766 434036 62772
rect 407764 61396 407816 61402
rect 407764 61338 407816 61344
rect 403624 60036 403676 60042
rect 403624 59978 403676 59984
rect 396448 58676 396500 58682
rect 396448 58618 396500 58624
rect 396460 54754 396488 58618
rect 442276 57322 442304 75618
rect 446416 74458 446444 77302
rect 449912 75614 449940 77316
rect 449900 75608 449952 75614
rect 449900 75550 449952 75556
rect 449912 75410 449940 75550
rect 449900 75404 449952 75410
rect 449900 75346 449952 75352
rect 446404 74452 446456 74458
rect 446404 74394 446456 74400
rect 446416 65754 446444 74394
rect 453776 74390 453804 77316
rect 453764 74384 453816 74390
rect 453764 74326 453816 74332
rect 453776 68406 453804 74326
rect 457640 74322 457668 77316
rect 457628 74316 457680 74322
rect 457628 74258 457680 74264
rect 457640 69766 457668 74258
rect 461504 74254 461532 77316
rect 465382 77302 465764 77330
rect 461492 74248 461544 74254
rect 461492 74190 461544 74196
rect 461504 73982 461532 74190
rect 465736 74186 465764 77302
rect 465724 74180 465776 74186
rect 465724 74122 465776 74128
rect 461492 73976 461544 73982
rect 461492 73918 461544 73924
rect 457628 69760 457680 69766
rect 457628 69702 457680 69708
rect 453764 68400 453816 68406
rect 453764 68342 453816 68348
rect 446404 65748 446456 65754
rect 446404 65690 446456 65696
rect 442264 57316 442316 57322
rect 442264 57258 442316 57264
rect 465736 57254 465764 74122
rect 469232 60110 469260 77316
rect 473096 74118 473124 77316
rect 476500 77302 476974 77330
rect 473084 74112 473136 74118
rect 473084 74054 473136 74060
rect 473096 71194 473124 74054
rect 473084 71188 473136 71194
rect 473084 71130 473136 71136
rect 476500 64874 476528 77302
rect 477880 74254 477908 204206
rect 478064 204202 478092 229066
rect 478156 204270 478184 332250
rect 478328 331288 478380 331294
rect 478328 331230 478380 331236
rect 478144 204264 478196 204270
rect 478340 204241 478368 331230
rect 478144 204206 478196 204212
rect 478326 204232 478382 204241
rect 477958 204167 478014 204176
rect 478052 204196 478104 204202
rect 477972 74458 478000 204167
rect 478326 204167 478382 204176
rect 478052 204138 478104 204144
rect 477960 74452 478012 74458
rect 477960 74394 478012 74400
rect 478064 74390 478092 204138
rect 478432 203969 478460 332726
rect 478984 332382 479012 459575
rect 479076 458969 479104 586094
rect 479156 585880 479208 585886
rect 479156 585822 479208 585828
rect 479168 462330 479196 585822
rect 481640 583432 481692 583438
rect 481640 583374 481692 583380
rect 480720 583296 480772 583302
rect 480720 583238 480772 583244
rect 480260 583024 480312 583030
rect 480260 582966 480312 582972
rect 480442 582992 480498 583001
rect 479246 533488 479302 533497
rect 479246 533423 479302 533432
rect 479156 462324 479208 462330
rect 479156 462266 479208 462272
rect 479260 460934 479288 533423
rect 479340 462324 479392 462330
rect 479340 462266 479392 462272
rect 479352 461106 479380 462266
rect 479340 461100 479392 461106
rect 479340 461042 479392 461048
rect 479168 460906 479288 460934
rect 479168 459338 479196 460906
rect 479156 459332 479208 459338
rect 479156 459274 479208 459280
rect 479062 458960 479118 458969
rect 479062 458895 479118 458904
rect 478972 332376 479024 332382
rect 478972 332318 479024 332324
rect 478880 331288 478932 331294
rect 478880 331230 478932 331236
rect 478418 203960 478474 203969
rect 478892 203930 478920 331230
rect 478984 203998 479012 332318
rect 479076 332246 479104 458895
rect 479168 333334 479196 459274
rect 479156 333328 479208 333334
rect 479156 333270 479208 333276
rect 479352 332518 479380 461042
rect 480272 459202 480300 582966
rect 480442 582927 480498 582936
rect 480456 462942 480484 582927
rect 480536 572076 480588 572082
rect 480536 572018 480588 572024
rect 480444 462936 480496 462942
rect 480444 462878 480496 462884
rect 480548 459270 480576 572018
rect 480628 462324 480680 462330
rect 480628 462266 480680 462272
rect 480640 461038 480668 462266
rect 480628 461032 480680 461038
rect 480628 460974 480680 460980
rect 480536 459264 480588 459270
rect 480536 459206 480588 459212
rect 480260 459196 480312 459202
rect 480260 459138 480312 459144
rect 480352 458856 480404 458862
rect 480352 458798 480404 458804
rect 479524 364404 479576 364410
rect 479524 364346 479576 364352
rect 479340 332512 479392 332518
rect 479340 332454 479392 332460
rect 479064 332240 479116 332246
rect 479064 332182 479116 332188
rect 479076 331294 479104 332182
rect 479064 331288 479116 331294
rect 479064 331230 479116 331236
rect 479062 329760 479118 329769
rect 479062 329695 479118 329704
rect 479076 204678 479104 329695
rect 479352 316034 479380 332454
rect 479168 316006 479380 316034
rect 479064 204672 479116 204678
rect 479064 204614 479116 204620
rect 478972 203992 479024 203998
rect 478972 203934 479024 203940
rect 478418 203895 478474 203904
rect 478880 203924 478932 203930
rect 478432 200114 478460 203895
rect 478880 203866 478932 203872
rect 478248 200086 478460 200114
rect 478248 78198 478276 200086
rect 478236 78192 478288 78198
rect 478236 78134 478288 78140
rect 478052 74384 478104 74390
rect 478052 74326 478104 74332
rect 477868 74248 477920 74254
rect 477868 74190 477920 74196
rect 478892 74186 478920 203866
rect 478984 74322 479012 203934
rect 479076 75546 479104 204614
rect 479168 203862 479196 316006
rect 479156 203856 479208 203862
rect 479156 203798 479208 203804
rect 479168 75614 479196 203798
rect 479536 78062 479564 364346
rect 480258 331800 480314 331809
rect 480258 331735 480314 331744
rect 480272 93854 480300 331735
rect 480364 315654 480392 458798
rect 480444 456748 480496 456754
rect 480444 456690 480496 456696
rect 480456 315994 480484 456690
rect 480548 333266 480576 459206
rect 480640 334014 480668 460974
rect 480732 457978 480760 583238
rect 480904 470620 480956 470626
rect 480904 470562 480956 470568
rect 480720 457972 480772 457978
rect 480720 457914 480772 457920
rect 480628 334008 480680 334014
rect 480628 333950 480680 333956
rect 480536 333260 480588 333266
rect 480536 333202 480588 333208
rect 480444 315988 480496 315994
rect 480444 315930 480496 315936
rect 480352 315648 480404 315654
rect 480352 315590 480404 315596
rect 480364 204746 480392 315590
rect 480456 206582 480484 315930
rect 480640 207641 480668 333950
rect 480626 207632 480682 207641
rect 480626 207567 480682 207576
rect 480444 206576 480496 206582
rect 480444 206518 480496 206524
rect 480720 205760 480772 205766
rect 480720 205702 480772 205708
rect 480352 204740 480404 204746
rect 480352 204682 480404 204688
rect 480364 200114 480392 204682
rect 480536 204128 480588 204134
rect 480536 204070 480588 204076
rect 480364 200086 480484 200114
rect 480272 93826 480392 93854
rect 479524 78056 479576 78062
rect 479524 77998 479576 78004
rect 480258 77344 480314 77353
rect 480258 77279 480260 77288
rect 480312 77279 480314 77288
rect 480260 77250 480312 77256
rect 479156 75608 479208 75614
rect 479156 75550 479208 75556
rect 479064 75540 479116 75546
rect 479064 75482 479116 75488
rect 480364 75342 480392 93826
rect 480456 75818 480484 200086
rect 480548 78130 480576 204070
rect 480626 149968 480682 149977
rect 480626 149903 480682 149912
rect 480536 78124 480588 78130
rect 480536 78066 480588 78072
rect 480444 75812 480496 75818
rect 480444 75754 480496 75760
rect 480352 75336 480404 75342
rect 480352 75278 480404 75284
rect 480640 74361 480668 149903
rect 480732 75750 480760 205702
rect 480916 204406 480944 470562
rect 481652 462330 481680 583374
rect 481824 583364 481876 583370
rect 481824 583306 481876 583312
rect 481732 572008 481784 572014
rect 481732 571950 481784 571956
rect 481640 462324 481692 462330
rect 481640 462266 481692 462272
rect 481640 458924 481692 458930
rect 481640 458866 481692 458872
rect 481178 207632 481234 207641
rect 481178 207567 481234 207576
rect 481192 207058 481220 207567
rect 481180 207052 481232 207058
rect 481180 206994 481232 207000
rect 480904 204400 480956 204406
rect 480904 204342 480956 204348
rect 480720 75744 480772 75750
rect 480720 75686 480772 75692
rect 481652 75177 481680 458866
rect 481744 458862 481772 571950
rect 481732 458856 481784 458862
rect 481732 458798 481784 458804
rect 481836 457910 481864 583306
rect 484400 583160 484452 583166
rect 484400 583102 484452 583108
rect 483020 583092 483072 583098
rect 483020 583034 483072 583040
rect 483032 459474 483060 583034
rect 483112 580372 483164 580378
rect 483112 580314 483164 580320
rect 483020 459468 483072 459474
rect 483020 459410 483072 459416
rect 482100 459196 482152 459202
rect 482100 459138 482152 459144
rect 481824 457904 481876 457910
rect 481824 457846 481876 457852
rect 481836 315722 481864 457846
rect 482008 333260 482060 333266
rect 482008 333202 482060 333208
rect 481916 332444 481968 332450
rect 481916 332386 481968 332392
rect 481824 315716 481876 315722
rect 481824 315658 481876 315664
rect 481732 315240 481784 315246
rect 481732 315182 481784 315188
rect 481744 204610 481772 315182
rect 481836 314702 481864 315658
rect 481824 314696 481876 314702
rect 481824 314638 481876 314644
rect 481732 204604 481784 204610
rect 481732 204546 481784 204552
rect 481638 75168 481694 75177
rect 481638 75103 481694 75112
rect 480626 74352 480682 74361
rect 478972 74316 479024 74322
rect 480626 74287 480682 74296
rect 478972 74258 479024 74264
rect 478880 74180 478932 74186
rect 478880 74122 478932 74128
rect 481744 73166 481772 204546
rect 481928 203833 481956 332386
rect 482020 205766 482048 333202
rect 482112 315926 482140 459138
rect 483032 458250 483060 459410
rect 483020 458244 483072 458250
rect 483020 458186 483072 458192
rect 483124 458114 483152 580314
rect 483204 580304 483256 580310
rect 483204 580246 483256 580252
rect 483216 460934 483244 580246
rect 483216 460906 483336 460934
rect 483308 458182 483336 460906
rect 484412 459406 484440 583102
rect 484400 459400 484452 459406
rect 484400 459342 484452 459348
rect 483296 458176 483348 458182
rect 483296 458118 483348 458124
rect 483112 458108 483164 458114
rect 483112 458050 483164 458056
rect 483124 456770 483152 458050
rect 483204 457972 483256 457978
rect 483204 457914 483256 457920
rect 483032 456742 483152 456770
rect 482100 315920 482152 315926
rect 482100 315862 482152 315868
rect 482112 315246 482140 315862
rect 483032 315353 483060 456742
rect 483216 456634 483244 457914
rect 483124 456606 483244 456634
rect 483124 315790 483152 456606
rect 483308 451274 483336 458118
rect 483216 451246 483336 451274
rect 483216 332722 483244 451246
rect 483204 332716 483256 332722
rect 483204 332658 483256 332664
rect 483112 315784 483164 315790
rect 483112 315726 483164 315732
rect 483018 315344 483074 315353
rect 483018 315279 483074 315288
rect 482100 315240 482152 315246
rect 482100 315182 482152 315188
rect 483020 207052 483072 207058
rect 483020 206994 483072 207000
rect 482008 205760 482060 205766
rect 482008 205702 482060 205708
rect 481914 203824 481970 203833
rect 481836 203782 481914 203810
rect 481836 74118 481864 203782
rect 481914 203759 481970 203768
rect 481916 203584 481968 203590
rect 481916 203526 481968 203532
rect 481928 75274 481956 203526
rect 483032 75682 483060 206994
rect 483124 204474 483152 315726
rect 483112 204468 483164 204474
rect 483112 204410 483164 204416
rect 483124 200114 483152 204410
rect 483216 201482 483244 332658
rect 484412 329730 484440 459342
rect 484492 458244 484544 458250
rect 484492 458186 484544 458192
rect 484504 329798 484532 458186
rect 484492 329792 484544 329798
rect 484492 329734 484544 329740
rect 484400 329724 484452 329730
rect 484400 329666 484452 329672
rect 484412 329458 484440 329666
rect 484400 329452 484452 329458
rect 484400 329394 484452 329400
rect 483388 314696 483440 314702
rect 483388 314638 483440 314644
rect 483400 204542 483428 314638
rect 484504 209774 484532 329734
rect 484584 329452 484636 329458
rect 484584 329394 484636 329400
rect 484412 209746 484532 209774
rect 483388 204536 483440 204542
rect 483388 204478 483440 204484
rect 483204 201476 483256 201482
rect 483204 201418 483256 201424
rect 483216 200666 483244 201418
rect 483204 200660 483256 200666
rect 483204 200602 483256 200608
rect 483124 200086 483336 200114
rect 483308 75954 483336 200086
rect 483296 75948 483348 75954
rect 483296 75890 483348 75896
rect 483020 75676 483072 75682
rect 483020 75618 483072 75624
rect 481916 75268 481968 75274
rect 481916 75210 481968 75216
rect 483400 74526 483428 204478
rect 484412 201414 484440 209746
rect 484400 201408 484452 201414
rect 484400 201350 484452 201356
rect 483388 74520 483440 74526
rect 483388 74462 483440 74468
rect 481824 74112 481876 74118
rect 481824 74054 481876 74060
rect 481732 73160 481784 73166
rect 481732 73102 481784 73108
rect 484412 73098 484440 201350
rect 484596 201346 484624 329394
rect 484584 201340 484636 201346
rect 484584 201282 484636 201288
rect 484596 200802 484624 201282
rect 484584 200796 484636 200802
rect 484584 200738 484636 200744
rect 484492 200660 484544 200666
rect 484492 200602 484544 200608
rect 484504 74497 484532 200602
rect 484490 74488 484546 74497
rect 484490 74423 484546 74432
rect 484400 73092 484452 73098
rect 484400 73034 484452 73040
rect 476132 64846 476528 64874
rect 469220 60104 469272 60110
rect 469220 60046 469272 60052
rect 476132 58682 476160 64846
rect 476120 58676 476172 58682
rect 476120 58618 476172 58624
rect 465724 57248 465776 57254
rect 465724 57190 465776 57196
rect 389836 54726 390218 54754
rect 391492 54726 391874 54754
rect 393332 54726 393530 54754
rect 394804 54726 395186 54754
rect 396460 54726 396842 54754
rect 335556 24274 335846 24290
rect 335544 24268 335846 24274
rect 335596 24262 335846 24268
rect 335544 24210 335596 24216
rect 364432 24200 364484 24206
rect 364484 24148 364550 24154
rect 364432 24142 364550 24148
rect 364444 24126 364550 24142
rect 367848 24138 368138 24154
rect 367836 24132 368138 24138
rect 367888 24126 368138 24132
rect 367836 24074 367888 24080
rect 266360 23520 266412 23526
rect 266360 23462 266412 23468
rect 267372 23520 267424 23526
rect 267424 23468 267674 23474
rect 267372 23462 267674 23468
rect 202892 23310 203090 23338
rect 205652 23310 206678 23338
rect 209792 23310 210266 23338
rect 212552 23310 213854 23338
rect 216692 23310 217442 23338
rect 220832 23310 221030 23338
rect 223592 23310 224618 23338
rect 200028 22092 200080 22098
rect 200028 22034 200080 22040
rect 156604 21548 156656 21554
rect 156604 21490 156656 21496
rect 149060 21480 149112 21486
rect 149060 21422 149112 21428
rect 138020 19984 138072 19990
rect 138020 19926 138072 19932
rect 131120 17332 131172 17338
rect 131120 17274 131172 17280
rect 131132 16574 131160 17274
rect 138032 16574 138060 19926
rect 149072 16574 149100 21422
rect 155960 21412 156012 21418
rect 155960 21354 156012 21360
rect 150440 18760 150492 18766
rect 150440 18702 150492 18708
rect 150452 16574 150480 18702
rect 151820 18692 151872 18698
rect 151820 18634 151872 18640
rect 131132 16546 131344 16574
rect 138032 16546 138888 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 125600 11892 125652 11898
rect 125600 11834 125652 11840
rect 96620 4888 96672 4894
rect 96620 4830 96672 4836
rect 92480 4820 92532 4826
rect 92480 4762 92532 4768
rect 66260 3460 66312 3466
rect 66260 3402 66312 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 11834
rect 128176 7608 128228 7614
rect 128176 7550 128228 7556
rect 128188 480 128216 7550
rect 129372 4956 129424 4962
rect 129372 4898 129424 4904
rect 129384 480 129412 4898
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 135260 15972 135312 15978
rect 135260 15914 135312 15920
rect 132960 7744 133012 7750
rect 132960 7686 133012 7692
rect 132972 480 133000 7686
rect 135272 480 135300 15914
rect 136456 14612 136508 14618
rect 136456 14554 136508 14560
rect 136468 480 136496 14554
rect 138860 480 138888 16546
rect 139584 13252 139636 13258
rect 139584 13194 139636 13200
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 13194
rect 142160 11756 142212 11762
rect 142160 11698 142212 11704
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 11698
rect 147128 10464 147180 10470
rect 147128 10406 147180 10412
rect 143540 6316 143592 6322
rect 143540 6258 143592 6264
rect 143552 480 143580 6258
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 145944 480 145972 3538
rect 147140 480 147168 10406
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 3534 151860 18634
rect 155972 16574 156000 21354
rect 155972 16546 156184 16574
rect 153752 11960 153804 11966
rect 153752 11902 153804 11908
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 153028 480 153056 3470
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 11902
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156616 10402 156644 21490
rect 178040 20120 178092 20126
rect 178040 20062 178092 20068
rect 169760 20052 169812 20058
rect 169760 19994 169812 20000
rect 169772 16574 169800 19994
rect 175280 18828 175332 18834
rect 175280 18770 175332 18776
rect 171140 17400 171192 17406
rect 171140 17342 171192 17348
rect 171152 16574 171180 17342
rect 175292 16574 175320 18770
rect 178052 16574 178080 20062
rect 184940 18624 184992 18630
rect 184940 18566 184992 18572
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 175292 16546 175504 16574
rect 178052 16546 178632 16574
rect 168380 16040 168432 16046
rect 168380 15982 168432 15988
rect 164424 14544 164476 14550
rect 164424 14486 164476 14492
rect 160100 13184 160152 13190
rect 160100 13126 160152 13132
rect 156604 10396 156656 10402
rect 156604 10338 156656 10344
rect 157800 7812 157852 7818
rect 157800 7754 157852 7760
rect 157812 480 157840 7754
rect 160112 3534 160140 13126
rect 163688 9104 163740 9110
rect 163688 9046 163740 9052
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 160100 2848 160152 2854
rect 160100 2790 160152 2796
rect 160112 480 160140 2790
rect 161308 480 161336 3470
rect 161400 2854 161428 3470
rect 161388 2848 161440 2854
rect 161388 2790 161440 2796
rect 163700 480 163728 9046
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14486
rect 167184 9036 167236 9042
rect 167184 8978 167236 8984
rect 167196 480 167224 8978
rect 168392 480 168420 15982
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 173900 14476 173952 14482
rect 173900 14418 173952 14424
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 14418
rect 175476 480 175504 16546
rect 176660 13116 176712 13122
rect 176660 13058 176712 13064
rect 176672 3398 176700 13058
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177868 480 177896 3334
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 181444 6248 181496 6254
rect 181444 6190 181496 6196
rect 181456 480 181484 6190
rect 182548 5024 182600 5030
rect 182548 4966 182600 4972
rect 182560 480 182588 4966
rect 184952 480 184980 18566
rect 202892 11898 202920 23310
rect 202880 11892 202932 11898
rect 202880 11834 202932 11840
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 186148 480 186176 11766
rect 188528 7676 188580 7682
rect 188528 7618 188580 7624
rect 188540 480 188568 7618
rect 205652 4962 205680 23310
rect 209792 7750 209820 23310
rect 212552 14618 212580 23310
rect 212540 14612 212592 14618
rect 212540 14554 212592 14560
rect 216692 13258 216720 23310
rect 216680 13252 216732 13258
rect 216680 13194 216732 13200
rect 217324 13252 217376 13258
rect 217324 13194 217376 13200
rect 209780 7744 209832 7750
rect 209780 7686 209832 7692
rect 205640 4956 205692 4962
rect 205640 4898 205692 4904
rect 217336 3602 217364 13194
rect 220832 6322 220860 23310
rect 223592 10470 223620 23310
rect 228192 18766 228220 23324
rect 230492 23310 231794 23338
rect 234632 23310 235382 23338
rect 238772 23310 238970 23338
rect 241532 23310 242558 23338
rect 245672 23310 246146 23338
rect 228180 18760 228232 18766
rect 228180 18702 228232 18708
rect 230492 11966 230520 23310
rect 230480 11960 230532 11966
rect 230480 11902 230532 11908
rect 223580 10464 223632 10470
rect 223580 10406 223632 10412
rect 234632 7818 234660 23310
rect 238772 13190 238800 23310
rect 241532 14550 241560 23310
rect 242900 17264 242952 17270
rect 242900 17206 242952 17212
rect 241520 14544 241572 14550
rect 241520 14486 241572 14492
rect 238760 13184 238812 13190
rect 238760 13126 238812 13132
rect 241704 8968 241756 8974
rect 241704 8910 241756 8916
rect 234620 7812 234672 7818
rect 234620 7754 234672 7760
rect 220820 6316 220872 6322
rect 220820 6258 220872 6264
rect 217324 3596 217376 3602
rect 217324 3538 217376 3544
rect 239312 3460 239364 3466
rect 239312 3402 239364 3408
rect 239324 480 239352 3402
rect 241716 480 241744 8910
rect 242912 480 242940 17206
rect 245672 16046 245700 23310
rect 249720 17406 249748 23324
rect 253308 18834 253336 23324
rect 256896 20126 256924 23324
rect 259472 23310 260498 23338
rect 263612 23310 264086 23338
rect 256884 20120 256936 20126
rect 256884 20062 256936 20068
rect 253296 18828 253348 18834
rect 253296 18770 253348 18776
rect 249708 17400 249760 17406
rect 249708 17342 249760 17348
rect 245660 16040 245712 16046
rect 245660 15982 245712 15988
rect 245936 15904 245988 15910
rect 245936 15846 245988 15852
rect 245200 10396 245252 10402
rect 245200 10338 245252 10344
rect 245212 480 245240 10338
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 15846
rect 249984 6180 250036 6186
rect 249984 6122 250036 6128
rect 248788 4820 248840 4826
rect 248788 4762 248840 4768
rect 248800 480 248828 4762
rect 249996 480 250024 6122
rect 259472 5030 259500 23310
rect 263612 11830 263640 23310
rect 263600 11824 263652 11830
rect 263600 11766 263652 11772
rect 259460 5024 259512 5030
rect 259460 4966 259512 4972
rect 252376 4888 252428 4894
rect 252376 4830 252428 4836
rect 252388 480 252416 4830
rect 266372 3466 266400 23462
rect 267384 23446 267674 23462
rect 270512 23310 271262 23338
rect 270512 7614 270540 23310
rect 274836 17338 274864 23324
rect 277412 23310 278438 23338
rect 274824 17332 274876 17338
rect 274824 17274 274876 17280
rect 277412 15978 277440 23310
rect 282012 19990 282040 23324
rect 284312 23310 285614 23338
rect 288452 23310 289202 23338
rect 282000 19984 282052 19990
rect 282000 19926 282052 19932
rect 277400 15972 277452 15978
rect 277400 15914 277452 15920
rect 284312 11762 284340 23310
rect 288452 13258 288480 23310
rect 292580 22772 292632 22778
rect 292580 22714 292632 22720
rect 292592 21826 292620 22714
rect 292580 21820 292632 21826
rect 292580 21762 292632 21768
rect 292776 21486 292804 23324
rect 292764 21480 292816 21486
rect 292764 21422 292816 21428
rect 296364 18698 296392 23324
rect 299952 21418 299980 23324
rect 302252 23310 303554 23338
rect 306392 23310 307142 23338
rect 310532 23310 310730 23338
rect 299940 21412 299992 21418
rect 299940 21354 299992 21360
rect 296352 18692 296404 18698
rect 296352 18634 296404 18640
rect 288440 13252 288492 13258
rect 288440 13194 288492 13200
rect 284300 11756 284352 11762
rect 284300 11698 284352 11704
rect 270500 7608 270552 7614
rect 270500 7550 270552 7556
rect 302252 3534 302280 23310
rect 306392 9110 306420 23310
rect 306380 9104 306432 9110
rect 306380 9046 306432 9052
rect 310532 9042 310560 23310
rect 314304 20058 314332 23324
rect 317432 23310 317906 23338
rect 320192 23310 321494 23338
rect 324332 23310 325082 23338
rect 314292 20052 314344 20058
rect 314292 19994 314344 20000
rect 317432 14482 317460 23310
rect 317420 14476 317472 14482
rect 317420 14418 317472 14424
rect 320192 13122 320220 23310
rect 320180 13116 320232 13122
rect 320180 13058 320232 13064
rect 310520 9036 310572 9042
rect 310520 8978 310572 8984
rect 324332 6254 324360 23310
rect 328656 18630 328684 23324
rect 331232 23310 332258 23338
rect 338132 23310 339434 23338
rect 328644 18624 328696 18630
rect 328644 18566 328696 18572
rect 331232 7682 331260 23310
rect 338132 10334 338160 23310
rect 343008 21894 343036 23324
rect 346596 21962 346624 23324
rect 350184 22166 350212 23324
rect 350172 22160 350224 22166
rect 350172 22102 350224 22108
rect 346584 21956 346636 21962
rect 346584 21898 346636 21904
rect 342996 21888 343048 21894
rect 342996 21830 343048 21836
rect 353772 21826 353800 23324
rect 357360 22001 357388 23324
rect 360948 22030 360976 23324
rect 371712 22137 371740 23324
rect 371698 22128 371754 22137
rect 371698 22063 371754 22072
rect 360936 22024 360988 22030
rect 357346 21992 357402 22001
rect 360936 21966 360988 21972
rect 357346 21927 357402 21936
rect 375300 21865 375328 23324
rect 378888 22098 378916 23324
rect 378876 22092 378928 22098
rect 378876 22034 378928 22040
rect 375286 21856 375342 21865
rect 353760 21820 353812 21826
rect 382476 21826 382504 23324
rect 386064 21894 386092 23324
rect 389652 22098 389680 23324
rect 389640 22092 389692 22098
rect 389640 22034 389692 22040
rect 393240 22030 393268 23324
rect 393228 22024 393280 22030
rect 393228 21966 393280 21972
rect 396828 21962 396856 23324
rect 396816 21956 396868 21962
rect 396816 21898 396868 21904
rect 386052 21888 386104 21894
rect 386052 21830 386104 21836
rect 485792 21826 485820 700266
rect 527192 697610 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 697604 527232 697610
rect 527180 697546 527232 697552
rect 527824 697604 527876 697610
rect 527824 697546 527876 697552
rect 485872 200796 485924 200802
rect 485872 200738 485924 200744
rect 485884 73030 485912 200738
rect 485872 73024 485924 73030
rect 485872 72966 485924 72972
rect 527836 21894 527864 697546
rect 542372 461009 542400 702406
rect 580172 697604 580224 697610
rect 580172 697546 580224 697552
rect 580184 697241 580212 697546
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580630 630864 580686 630873
rect 580630 630799 580686 630808
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 577318 579660 577623
rect 577504 577312 577556 577318
rect 577504 577254 577556 577260
rect 579620 577312 579672 577318
rect 579620 577254 579672 577260
rect 542358 461000 542414 461009
rect 542358 460935 542414 460944
rect 577516 332654 577544 577254
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 577504 332648 577556 332654
rect 577504 332590 577556 332596
rect 579618 78432 579674 78441
rect 579618 78367 579674 78376
rect 579632 77994 579660 78367
rect 579620 77988 579672 77994
rect 579620 77930 579672 77936
rect 580276 22098 580304 590951
rect 580538 524512 580594 524521
rect 580538 524447 580594 524456
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 580264 22092 580316 22098
rect 580264 22034 580316 22040
rect 580368 22030 580396 484599
rect 580446 378448 580502 378457
rect 580446 378383 580502 378392
rect 580356 22024 580408 22030
rect 580356 21966 580408 21972
rect 580460 21962 580488 378383
rect 580552 204338 580580 524447
rect 580644 332489 580672 630799
rect 580920 591025 580948 643991
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 484673 580948 537775
rect 580906 484664 580962 484673
rect 580906 484599 580962 484608
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 378457 580948 431559
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580630 332480 580686 332489
rect 580630 332415 580686 332424
rect 580540 204332 580592 204338
rect 580540 204274 580592 204280
rect 580448 21956 580500 21962
rect 580448 21898 580500 21904
rect 527824 21888 527876 21894
rect 527824 21830 527876 21836
rect 375286 21791 375342 21800
rect 382464 21820 382516 21826
rect 353760 21762 353812 21768
rect 382464 21762 382516 21768
rect 485780 21820 485832 21826
rect 485780 21762 485832 21768
rect 338120 10328 338172 10334
rect 338120 10270 338172 10276
rect 331220 7676 331272 7682
rect 331220 7618 331272 7624
rect 324320 6248 324372 6254
rect 324320 6190 324372 6196
rect 302240 3528 302292 3534
rect 302240 3470 302292 3476
rect 266360 3460 266412 3466
rect 266360 3402 266412 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 671220 3478 671256
rect 3422 671200 3424 671220
rect 3424 671200 3476 671220
rect 3476 671200 3478 671220
rect 2778 658144 2834 658200
rect 3606 619112 3662 619168
rect 2778 607144 2834 607200
rect 2778 566888 2834 566944
rect 2778 553832 2834 553888
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 2778 502288 2834 502344
rect 3422 502288 3478 502344
rect 2778 501744 2834 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 2778 449520 2834 449576
rect 2870 410488 2926 410544
rect 2778 398792 2834 398848
rect 3330 345344 3386 345400
rect 2778 293120 2834 293176
rect 3330 241032 3386 241088
rect 2778 188808 2834 188864
rect 3330 149776 3386 149832
rect 2778 136740 2834 136776
rect 2778 136720 2780 136740
rect 2780 136720 2832 136740
rect 2832 136720 2834 136740
rect 3330 110608 3386 110664
rect 3330 84632 3386 84688
rect 3330 32408 3386 32464
rect 3514 398792 3570 398848
rect 3514 397432 3570 397488
rect 3606 319232 3662 319288
rect 3606 267144 3662 267200
rect 3698 214920 3754 214976
rect 3606 45464 3662 45520
rect 4894 204040 4950 204096
rect 4802 75656 4858 75712
rect 3790 71576 3846 71632
rect 19246 585656 19302 585712
rect 18878 204176 18934 204232
rect 21638 460808 21694 460864
rect 20350 205692 20406 205728
rect 20350 205672 20352 205692
rect 20352 205672 20404 205692
rect 20404 205672 20406 205692
rect 20902 110336 20958 110392
rect 72974 700304 73030 700360
rect 27250 586336 27306 586392
rect 22650 459448 22706 459504
rect 57518 585792 57574 585848
rect 61382 585656 61438 585712
rect 96158 585656 96214 585712
rect 84566 582936 84622 582992
rect 112258 582936 112314 582992
rect 133878 572056 133934 572112
rect 69018 571920 69074 571976
rect 195978 571920 196034 571976
rect 23478 458768 23534 458824
rect 42062 460808 42118 460864
rect 38198 459448 38254 459504
rect 69110 458904 69166 458960
rect 84566 458768 84622 458824
rect 57518 458088 57574 458144
rect 112258 458088 112314 458144
rect 181810 460808 181866 460864
rect 185674 460672 185730 460728
rect 193126 459448 193182 459504
rect 197358 459348 197360 459368
rect 197360 459348 197412 459368
rect 197412 459348 197414 459368
rect 197358 459312 197414 459348
rect 197266 458904 197322 458960
rect 189538 458768 189594 458824
rect 173806 457952 173862 458008
rect 198186 460808 198242 460864
rect 198002 457952 198058 458008
rect 21546 110336 21602 110392
rect 57518 332288 57574 332344
rect 69110 332424 69166 332480
rect 96434 331744 96490 331800
rect 189538 331880 189594 331936
rect 197358 332732 197360 332752
rect 197360 332732 197412 332752
rect 197412 332732 197414 332752
rect 197358 332696 197414 332732
rect 22834 203496 22890 203552
rect 22374 202852 22376 202872
rect 22376 202852 22428 202872
rect 22428 202852 22430 202872
rect 22374 202816 22430 202852
rect 26606 204040 26662 204096
rect 30470 203496 30526 203552
rect 88430 204176 88486 204232
rect 69110 202816 69166 202872
rect 57518 202680 57574 202736
rect 115754 204176 115810 204232
rect 183466 204312 183522 204368
rect 179878 203496 179934 203552
rect 195886 203904 195942 203960
rect 197818 202952 197874 203008
rect 198002 204312 198058 204368
rect 26606 75656 26662 75712
rect 50342 75112 50398 75168
rect 57242 74432 57298 74488
rect 81254 75792 81310 75848
rect 57058 61512 57114 61568
rect 103058 59608 103114 59664
rect 102782 58520 102838 58576
rect 102598 56616 102654 56672
rect 57518 56344 57574 56400
rect 102230 54168 102286 54224
rect 102138 53488 102194 53544
rect 102138 52556 102194 52592
rect 102138 52536 102140 52556
rect 102140 52536 102192 52556
rect 102192 52536 102194 52556
rect 57058 51720 57114 51776
rect 102966 55528 103022 55584
rect 198922 203496 198978 203552
rect 198738 201320 198794 201376
rect 197818 63452 197820 63472
rect 197820 63452 197872 63472
rect 197872 63452 197874 63472
rect 197818 63416 197874 63452
rect 103242 51040 103298 51096
rect 103058 49816 103114 49872
rect 102690 46960 102746 47016
rect 57518 46860 57520 46880
rect 57520 46860 57572 46880
rect 57572 46860 57574 46880
rect 57518 46824 57574 46860
rect 102506 44376 102562 44432
rect 102322 43288 102378 43344
rect 57150 42064 57206 42120
rect 102138 41384 102194 41440
rect 102230 40024 102286 40080
rect 102138 37848 102194 37904
rect 57058 36896 57114 36952
rect 102414 42880 102470 42936
rect 102782 45736 102838 45792
rect 103426 48728 103482 48784
rect 195978 51312 196034 51368
rect 195978 50904 196034 50960
rect 195978 49408 196034 49464
rect 195978 48220 195980 48240
rect 195980 48220 196032 48240
rect 196032 48220 196034 48240
rect 195978 48184 196034 48220
rect 196070 47640 196126 47696
rect 195978 46860 195980 46880
rect 195980 46860 196032 46880
rect 196032 46860 196034 46880
rect 195978 46824 196034 46860
rect 196162 46144 196218 46200
rect 195978 45192 196034 45248
rect 195978 43968 196034 44024
rect 196070 43560 196126 43616
rect 195978 41520 196034 41576
rect 195978 41112 196034 41168
rect 195978 39888 196034 39944
rect 196070 39480 196126 39536
rect 102874 38936 102930 38992
rect 102598 37304 102654 37360
rect 102138 34584 102194 34640
rect 102782 36080 102838 36136
rect 195978 38392 196034 38448
rect 196070 37984 196126 38040
rect 195978 37032 196034 37088
rect 195978 35844 195980 35864
rect 195980 35844 196032 35864
rect 196032 35844 196034 35864
rect 195978 35808 196034 35844
rect 196070 35400 196126 35456
rect 195978 34312 196034 34368
rect 196070 33768 196126 33824
rect 102322 33496 102378 33552
rect 102138 32408 102194 32464
rect 57610 31592 57666 31648
rect 57242 27104 57298 27160
rect 102230 31728 102286 31784
rect 195978 32952 196034 33008
rect 102138 30504 102194 30560
rect 195978 31592 196034 31648
rect 196070 31184 196126 31240
rect 195978 30268 195980 30288
rect 195980 30268 196032 30288
rect 196032 30268 196034 30288
rect 195978 30232 196034 30268
rect 196070 29688 196126 29744
rect 102138 29280 102194 29336
rect 195978 28908 195980 28928
rect 195980 28908 196032 28928
rect 196032 28908 196034 28928
rect 195978 28872 196034 28908
rect 102138 28464 102194 28520
rect 195978 28056 196034 28112
rect 102138 27648 102194 27704
rect 195978 27240 196034 27296
rect 102782 26288 102838 26344
rect 195978 26188 195980 26208
rect 195980 26188 196032 26208
rect 196032 26188 196034 26208
rect 195978 26152 196034 26188
rect 3422 6432 3478 6488
rect 218058 586336 218114 586392
rect 306930 586336 306986 586392
rect 258722 585656 258778 585712
rect 200302 460672 200358 460728
rect 200302 459584 200358 459640
rect 200210 459448 200266 459504
rect 200486 459448 200542 459504
rect 200670 459584 200726 459640
rect 200486 315968 200542 316024
rect 200394 203904 200450 203960
rect 200578 203904 200634 203960
rect 202970 204176 203026 204232
rect 233882 331880 233938 331936
rect 258078 331744 258134 331800
rect 283654 458904 283710 458960
rect 266358 331744 266414 331800
rect 283838 458768 283894 458824
rect 299294 314744 299350 314800
rect 299478 315288 299534 315344
rect 300582 462168 300638 462224
rect 300306 332424 300362 332480
rect 300214 205672 300270 205728
rect 300582 315868 300584 315888
rect 300584 315868 300636 315888
rect 300636 315868 300638 315888
rect 300582 315832 300638 315868
rect 301870 459312 301926 459368
rect 301686 459176 301742 459232
rect 301502 458224 301558 458280
rect 301594 457000 301650 457056
rect 301870 458224 301926 458280
rect 302054 585656 302110 585712
rect 302054 458088 302110 458144
rect 301870 456864 301926 456920
rect 302698 459448 302754 459504
rect 302146 457816 302202 457872
rect 302054 457000 302110 457056
rect 302146 456864 302202 456920
rect 300490 204176 300546 204232
rect 300030 64812 300032 64832
rect 300032 64812 300084 64832
rect 300084 64812 300086 64832
rect 300030 64776 300086 64812
rect 300766 204176 300822 204232
rect 337842 582936 337898 582992
rect 349434 585656 349490 585712
rect 391938 582936 391994 582992
rect 430578 585656 430634 585712
rect 469218 585792 469274 585848
rect 477866 586336 477922 586392
rect 476946 585112 477002 585168
rect 303066 460944 303122 461000
rect 306930 460808 306986 460864
rect 318522 459448 318578 459504
rect 314658 459312 314714 459368
rect 310794 459176 310850 459232
rect 349434 458088 349490 458144
rect 337842 457952 337898 458008
rect 322386 457816 322442 457872
rect 461490 459584 461546 459640
rect 469310 458904 469366 458960
rect 463790 458768 463846 458824
rect 476946 458224 477002 458280
rect 302882 332424 302938 332480
rect 303066 332424 303122 332480
rect 303526 315596 303528 315616
rect 303528 315596 303580 315616
rect 303580 315596 303582 315616
rect 303526 315560 303582 315596
rect 372618 331744 372674 331800
rect 469218 331744 469274 331800
rect 478142 458768 478198 458824
rect 476946 331200 477002 331256
rect 477498 329704 477554 329760
rect 387798 315288 387854 315344
rect 476118 315288 476174 315344
rect 478970 459584 479026 459640
rect 478878 456864 478934 456920
rect 442354 206624 442410 206680
rect 298742 57296 298798 57352
rect 476118 205692 476174 205728
rect 476118 205672 476120 205692
rect 476120 205672 476172 205692
rect 476172 205672 476174 205692
rect 337842 204312 337898 204368
rect 345570 204040 345626 204096
rect 364890 204176 364946 204232
rect 430578 204176 430634 204232
rect 446034 204040 446090 204096
rect 475382 204176 475438 204232
rect 475382 203904 475438 203960
rect 476026 203768 476082 203824
rect 477498 202836 477554 202872
rect 477498 202816 477500 202836
rect 477500 202816 477552 202836
rect 477552 202816 477554 202836
rect 303342 77288 303398 77344
rect 311162 77288 311218 77344
rect 393318 78104 393374 78160
rect 390558 77968 390614 78024
rect 336738 77832 336794 77888
rect 337474 77832 337530 77888
rect 389178 77832 389234 77888
rect 336830 75112 336886 75168
rect 346766 58520 346822 58576
rect 373998 75112 374054 75168
rect 371974 57296 372030 57352
rect 388534 57160 388590 57216
rect 392582 74296 392638 74352
rect 395802 74432 395858 74488
rect 399482 73072 399538 73128
rect 477958 204176 478014 204232
rect 478326 204176 478382 204232
rect 479246 533432 479302 533488
rect 479062 458904 479118 458960
rect 478418 203904 478474 203960
rect 480442 582936 480498 582992
rect 479062 329704 479118 329760
rect 480258 331744 480314 331800
rect 480626 207576 480682 207632
rect 480258 77308 480314 77344
rect 480258 77288 480260 77308
rect 480260 77288 480312 77308
rect 480312 77288 480314 77308
rect 480626 149912 480682 149968
rect 481178 207576 481234 207632
rect 481638 75112 481694 75168
rect 480626 74296 480682 74352
rect 483018 315288 483074 315344
rect 481914 203768 481970 203824
rect 484490 74432 484546 74488
rect 371698 22072 371754 22128
rect 357346 21936 357402 21992
rect 375286 21800 375342 21856
rect 580170 697176 580226 697232
rect 580906 644000 580962 644056
rect 580630 630808 580686 630864
rect 580262 590960 580318 591016
rect 579618 577632 579674 577688
rect 542358 460944 542414 461000
rect 580170 471416 580226 471472
rect 580170 365064 580226 365120
rect 579618 78376 579674 78432
rect 580538 524456 580594 524512
rect 580354 484608 580410 484664
rect 580446 378392 580502 378448
rect 580906 590960 580962 591016
rect 580906 537784 580962 537840
rect 580906 484608 580962 484664
rect 580906 431568 580962 431624
rect 580906 378392 580962 378448
rect 580630 332424 580686 332480
<< metal3 >>
rect 72969 700362 73035 700365
rect 199326 700362 199332 700364
rect 72969 700360 199332 700362
rect 72969 700304 72974 700360
rect 73030 700304 199332 700360
rect 72969 700302 199332 700304
rect 72969 700299 73035 700302
rect 199326 700300 199332 700302
rect 199396 700300 199402 700364
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 583520 683906 584960 683996
rect 583342 683846 584960 683906
rect 583342 683770 583402 683846
rect 583520 683770 584960 683846
rect 583342 683756 584960 683770
rect 583342 683710 583586 683756
rect 479374 683164 479380 683228
rect 479444 683226 479450 683228
rect 583526 683226 583586 683710
rect 479444 683166 583586 683226
rect 479444 683164 479450 683166
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580625 630866 580691 630869
rect 583520 630866 584960 630956
rect 580625 630864 584960 630866
rect 580625 630808 580630 630864
rect 580686 630808 584960 630864
rect 580625 630806 584960 630808
rect 580625 630803 580691 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 583520 617388 584960 617628
rect 2773 607202 2839 607205
rect 3366 607202 3372 607204
rect 2773 607200 3372 607202
rect 2773 607144 2778 607200
rect 2834 607144 3372 607200
rect 2773 607142 3372 607144
rect 2773 607139 2839 607142
rect 3366 607140 3372 607142
rect 3436 607140 3442 607204
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580257 591018 580323 591021
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 580906 591016
rect 580962 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect 27245 586394 27311 586397
rect 218053 586394 218119 586397
rect 27245 586392 218119 586394
rect 27245 586336 27250 586392
rect 27306 586336 218058 586392
rect 218114 586336 218119 586392
rect 27245 586334 218119 586336
rect 27245 586331 27311 586334
rect 218053 586331 218119 586334
rect 306925 586394 306991 586397
rect 477861 586394 477927 586397
rect 306925 586392 477927 586394
rect 306925 586336 306930 586392
rect 306986 586336 477866 586392
rect 477922 586336 477927 586392
rect 306925 586334 477927 586336
rect 306925 586331 306991 586334
rect 477861 586331 477927 586334
rect 23238 585788 23244 585852
rect 23308 585850 23314 585852
rect 57513 585850 57579 585853
rect 23308 585848 57579 585850
rect 23308 585792 57518 585848
rect 57574 585792 57579 585848
rect 23308 585790 57579 585792
rect 23308 585788 23314 585790
rect 57513 585787 57579 585790
rect 469213 585850 469279 585853
rect 480294 585850 480300 585852
rect 469213 585848 480300 585850
rect 469213 585792 469218 585848
rect 469274 585792 480300 585848
rect 469213 585790 480300 585792
rect 469213 585787 469279 585790
rect 480294 585788 480300 585790
rect 480364 585788 480370 585852
rect 19241 585714 19307 585717
rect 61377 585714 61443 585717
rect 19241 585712 61443 585714
rect 19241 585656 19246 585712
rect 19302 585656 61382 585712
rect 61438 585656 61443 585712
rect 19241 585654 61443 585656
rect 19241 585651 19307 585654
rect 61377 585651 61443 585654
rect 96153 585714 96219 585717
rect 258717 585714 258783 585717
rect 96153 585712 258783 585714
rect 96153 585656 96158 585712
rect 96214 585656 258722 585712
rect 258778 585656 258783 585712
rect 96153 585654 258783 585656
rect 96153 585651 96219 585654
rect 258717 585651 258783 585654
rect 302049 585714 302115 585717
rect 349429 585714 349495 585717
rect 302049 585712 349495 585714
rect 302049 585656 302054 585712
rect 302110 585656 349434 585712
rect 349490 585656 349495 585712
rect 302049 585654 349495 585656
rect 302049 585651 302115 585654
rect 349429 585651 349495 585654
rect 430573 585714 430639 585717
rect 476614 585714 476620 585716
rect 430573 585712 476620 585714
rect 430573 585656 430578 585712
rect 430634 585656 476620 585712
rect 430573 585654 476620 585656
rect 430573 585651 430639 585654
rect 476614 585652 476620 585654
rect 476684 585652 476690 585716
rect 476941 585170 477007 585173
rect 481582 585170 481588 585172
rect 476941 585168 481588 585170
rect 476941 585112 476946 585168
rect 477002 585112 481588 585168
rect 476941 585110 481588 585112
rect 476941 585107 477007 585110
rect 481582 585108 481588 585110
rect 481652 585108 481658 585172
rect 23054 582932 23060 582996
rect 23124 582994 23130 582996
rect 84561 582994 84627 582997
rect 23124 582992 84627 582994
rect 23124 582936 84566 582992
rect 84622 582936 84627 582992
rect 23124 582934 84627 582936
rect 23124 582932 23130 582934
rect 84561 582931 84627 582934
rect 112253 582994 112319 582997
rect 199878 582994 199884 582996
rect 112253 582992 199884 582994
rect 112253 582936 112258 582992
rect 112314 582936 199884 582992
rect 112253 582934 199884 582936
rect 112253 582931 112319 582934
rect 199878 582932 199884 582934
rect 199948 582932 199954 582996
rect 303470 582932 303476 582996
rect 303540 582994 303546 582996
rect 337837 582994 337903 582997
rect 303540 582992 337903 582994
rect 303540 582936 337842 582992
rect 337898 582936 337903 582992
rect 303540 582934 337903 582936
rect 303540 582932 303546 582934
rect 337837 582931 337903 582934
rect 391933 582994 391999 582997
rect 480437 582994 480503 582997
rect 391933 582992 480503 582994
rect 391933 582936 391938 582992
rect 391994 582936 480442 582992
rect 480498 582936 480503 582992
rect 391933 582934 480503 582936
rect 391933 582931 391999 582934
rect 480437 582931 480503 582934
rect -960 579852 480 580092
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect 133873 572114 133939 572117
rect 197302 572114 197308 572116
rect 133873 572112 197308 572114
rect 133873 572056 133878 572112
rect 133934 572056 197308 572112
rect 133873 572054 197308 572056
rect 133873 572051 133939 572054
rect 197302 572052 197308 572054
rect 197372 572052 197378 572116
rect 21950 571916 21956 571980
rect 22020 571978 22026 571980
rect 69013 571978 69079 571981
rect 22020 571976 69079 571978
rect 22020 571920 69018 571976
rect 69074 571920 69079 571976
rect 22020 571918 69079 571920
rect 22020 571916 22026 571918
rect 69013 571915 69079 571918
rect 195973 571978 196039 571981
rect 298870 571978 298876 571980
rect 195973 571976 298876 571978
rect 195973 571920 195978 571976
rect 196034 571920 298876 571976
rect 195973 571918 298876 571920
rect 195973 571915 196039 571918
rect 298870 571916 298876 571918
rect 298940 571916 298946 571980
rect -960 566946 480 567036
rect 2773 566946 2839 566949
rect -960 566944 2839 566946
rect -960 566888 2778 566944
rect 2834 566888 2839 566944
rect -960 566886 2839 566888
rect -960 566796 480 566886
rect 2773 566883 2839 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect 477534 533428 477540 533492
rect 477604 533490 477610 533492
rect 479241 533490 479307 533493
rect 477604 533488 479307 533490
rect 477604 533432 479246 533488
rect 479302 533432 479307 533488
rect 477604 533430 479307 533432
rect 477604 533428 477610 533430
rect 479241 533427 479307 533430
rect -960 527764 480 528004
rect 580533 524514 580599 524517
rect 583520 524514 584960 524604
rect 580533 524512 584960 524514
rect 580533 524456 580538 524512
rect 580594 524456 584960 524512
rect 580533 524454 584960 524456
rect 580533 524451 580599 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 583520 511172 584960 511412
rect 2773 502346 2839 502349
rect 3417 502346 3483 502349
rect 2773 502344 3483 502346
rect 2773 502288 2778 502344
rect 2834 502288 3422 502344
rect 3478 502288 3483 502344
rect 2773 502286 3483 502288
rect 2773 502283 2839 502286
rect 3417 502283 3483 502286
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580349 484666 580415 484669
rect 580901 484666 580967 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 580906 484664
rect 580962 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 580901 484603 580967 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 299974 462164 299980 462228
rect 300044 462226 300050 462228
rect 300577 462226 300643 462229
rect 300044 462224 300643 462226
rect 300044 462168 300582 462224
rect 300638 462168 300643 462224
rect 300044 462166 300643 462168
rect 300044 462164 300050 462166
rect 300577 462163 300643 462166
rect 303061 461002 303127 461005
rect 542353 461002 542419 461005
rect 303061 461000 542419 461002
rect 303061 460944 303066 461000
rect 303122 460944 542358 461000
rect 542414 460944 542419 461000
rect 303061 460942 542419 460944
rect 303061 460939 303127 460942
rect 542353 460939 542419 460942
rect 21633 460866 21699 460869
rect 42057 460866 42123 460869
rect 21633 460864 42123 460866
rect 21633 460808 21638 460864
rect 21694 460808 42062 460864
rect 42118 460808 42123 460864
rect 21633 460806 42123 460808
rect 21633 460803 21699 460806
rect 42057 460803 42123 460806
rect 181805 460866 181871 460869
rect 198181 460866 198247 460869
rect 181805 460864 198247 460866
rect 181805 460808 181810 460864
rect 181866 460808 198186 460864
rect 198242 460808 198247 460864
rect 181805 460806 198247 460808
rect 181805 460803 181871 460806
rect 198181 460803 198247 460806
rect 306925 460866 306991 460869
rect 479374 460866 479380 460868
rect 306925 460864 479380 460866
rect 306925 460808 306930 460864
rect 306986 460808 479380 460864
rect 306925 460806 479380 460808
rect 306925 460803 306991 460806
rect 479374 460804 479380 460806
rect 479444 460804 479450 460868
rect 185669 460730 185735 460733
rect 200297 460730 200363 460733
rect 185669 460728 200363 460730
rect 185669 460672 185674 460728
rect 185730 460672 200302 460728
rect 200358 460672 200363 460728
rect 185669 460670 200363 460672
rect 185669 460667 185735 460670
rect 200297 460667 200363 460670
rect 200297 459642 200363 459645
rect 200665 459642 200731 459645
rect 200297 459640 200731 459642
rect 200297 459584 200302 459640
rect 200358 459584 200670 459640
rect 200726 459584 200731 459640
rect 200297 459582 200731 459584
rect 200297 459579 200363 459582
rect 200665 459579 200731 459582
rect 461485 459642 461551 459645
rect 478965 459642 479031 459645
rect 461485 459640 479031 459642
rect 461485 459584 461490 459640
rect 461546 459584 478970 459640
rect 479026 459584 479031 459640
rect 461485 459582 479031 459584
rect 461485 459579 461551 459582
rect 478965 459579 479031 459582
rect 22645 459506 22711 459509
rect 38193 459506 38259 459509
rect 22645 459504 38259 459506
rect 22645 459448 22650 459504
rect 22706 459448 38198 459504
rect 38254 459448 38259 459504
rect 22645 459446 38259 459448
rect 22645 459443 22711 459446
rect 38193 459443 38259 459446
rect 193121 459506 193187 459509
rect 200205 459506 200271 459509
rect 200481 459506 200547 459509
rect 193121 459504 200547 459506
rect 193121 459448 193126 459504
rect 193182 459448 200210 459504
rect 200266 459448 200486 459504
rect 200542 459448 200547 459504
rect 193121 459446 200547 459448
rect 193121 459443 193187 459446
rect 200205 459443 200271 459446
rect 200481 459443 200547 459446
rect 302693 459506 302759 459509
rect 318517 459506 318583 459509
rect 302693 459504 318583 459506
rect 302693 459448 302698 459504
rect 302754 459448 318522 459504
rect 318578 459448 318583 459504
rect 302693 459446 318583 459448
rect 302693 459443 302759 459446
rect 318517 459443 318583 459446
rect 197353 459370 197419 459373
rect 197854 459370 197860 459372
rect 197353 459368 197860 459370
rect 197353 459312 197358 459368
rect 197414 459312 197860 459368
rect 197353 459310 197860 459312
rect 197353 459307 197419 459310
rect 197854 459308 197860 459310
rect 197924 459308 197930 459372
rect 301865 459370 301931 459373
rect 314653 459370 314719 459373
rect 301865 459368 314719 459370
rect 301865 459312 301870 459368
rect 301926 459312 314658 459368
rect 314714 459312 314719 459368
rect 301865 459310 314719 459312
rect 301865 459307 301931 459310
rect 314653 459307 314719 459310
rect 301681 459234 301747 459237
rect 310789 459234 310855 459237
rect 301681 459232 310855 459234
rect 301681 459176 301686 459232
rect 301742 459176 310794 459232
rect 310850 459176 310855 459232
rect 301681 459174 310855 459176
rect 301681 459171 301747 459174
rect 310789 459171 310855 459174
rect 22870 458900 22876 458964
rect 22940 458962 22946 458964
rect 69105 458962 69171 458965
rect 22940 458960 69171 458962
rect 22940 458904 69110 458960
rect 69166 458904 69171 458960
rect 22940 458902 69171 458904
rect 22940 458900 22946 458902
rect 69105 458899 69171 458902
rect 197261 458962 197327 458965
rect 283649 458962 283715 458965
rect 197261 458960 283715 458962
rect 197261 458904 197266 458960
rect 197322 458904 283654 458960
rect 283710 458904 283715 458960
rect 197261 458902 283715 458904
rect 197261 458899 197327 458902
rect 283649 458899 283715 458902
rect 469305 458962 469371 458965
rect 479057 458962 479123 458965
rect 469305 458960 479123 458962
rect 469305 458904 469310 458960
rect 469366 458904 479062 458960
rect 479118 458904 479123 458960
rect 469305 458902 479123 458904
rect 469305 458899 469371 458902
rect 479057 458899 479123 458902
rect 23054 458764 23060 458828
rect 23124 458826 23130 458828
rect 23473 458826 23539 458829
rect 84561 458826 84627 458829
rect 23124 458824 84627 458826
rect 23124 458768 23478 458824
rect 23534 458768 84566 458824
rect 84622 458768 84627 458824
rect 23124 458766 84627 458768
rect 23124 458764 23130 458766
rect 23473 458763 23539 458766
rect 84561 458763 84627 458766
rect 189533 458826 189599 458829
rect 283833 458826 283899 458829
rect 189533 458824 283899 458826
rect 189533 458768 189538 458824
rect 189594 458768 283838 458824
rect 283894 458768 283899 458824
rect 189533 458766 283899 458768
rect 189533 458763 189599 458766
rect 283833 458763 283899 458766
rect 463785 458826 463851 458829
rect 478137 458826 478203 458829
rect 463785 458824 478203 458826
rect 463785 458768 463790 458824
rect 463846 458768 478142 458824
rect 478198 458768 478203 458824
rect 463785 458766 478203 458768
rect 463785 458763 463851 458766
rect 478137 458763 478203 458766
rect 21950 458220 21956 458284
rect 22020 458282 22026 458284
rect 22870 458282 22876 458284
rect 22020 458222 22876 458282
rect 22020 458220 22026 458222
rect 22870 458220 22876 458222
rect 22940 458220 22946 458284
rect 301497 458282 301563 458285
rect 301865 458282 301931 458285
rect 301497 458280 301931 458282
rect 301497 458224 301502 458280
rect 301558 458224 301870 458280
rect 301926 458224 301931 458280
rect 301497 458222 301931 458224
rect 301497 458219 301563 458222
rect 301865 458219 301931 458222
rect 476941 458282 477007 458285
rect 478822 458282 478828 458284
rect 476941 458280 478828 458282
rect 476941 458224 476946 458280
rect 477002 458224 478828 458280
rect 476941 458222 478828 458224
rect 476941 458219 477007 458222
rect 478822 458220 478828 458222
rect 478892 458220 478898 458284
rect 23238 458084 23244 458148
rect 23308 458146 23314 458148
rect 57513 458146 57579 458149
rect 23308 458144 57579 458146
rect 23308 458088 57518 458144
rect 57574 458088 57579 458144
rect 23308 458086 57579 458088
rect 23308 458084 23314 458086
rect 57513 458083 57579 458086
rect 112253 458146 112319 458149
rect 199878 458146 199884 458148
rect 112253 458144 199884 458146
rect 112253 458088 112258 458144
rect 112314 458088 199884 458144
rect 112253 458086 199884 458088
rect 112253 458083 112319 458086
rect 199878 458084 199884 458086
rect 199948 458084 199954 458148
rect 302049 458146 302115 458149
rect 349429 458146 349495 458149
rect 302049 458144 349495 458146
rect 302049 458088 302054 458144
rect 302110 458088 349434 458144
rect 349490 458088 349495 458144
rect 302049 458086 349495 458088
rect 302049 458083 302115 458086
rect 349429 458083 349495 458086
rect 173801 458010 173867 458013
rect 197997 458010 198063 458013
rect 173801 458008 198063 458010
rect 173801 457952 173806 458008
rect 173862 457952 198002 458008
rect 198058 457952 198063 458008
rect 173801 457950 198063 457952
rect 173801 457947 173867 457950
rect 197997 457947 198063 457950
rect 303470 457948 303476 458012
rect 303540 458010 303546 458012
rect 337837 458010 337903 458013
rect 303540 458008 337903 458010
rect 303540 457952 337842 458008
rect 337898 457952 337903 458008
rect 583520 457996 584960 458236
rect 303540 457950 337903 457952
rect 303540 457948 303546 457950
rect 337837 457947 337903 457950
rect 302141 457874 302207 457877
rect 322381 457874 322447 457877
rect 302141 457872 322447 457874
rect 302141 457816 302146 457872
rect 302202 457816 322386 457872
rect 322442 457816 322447 457872
rect 302141 457814 322447 457816
rect 302141 457811 302207 457814
rect 322381 457811 322447 457814
rect 301589 457058 301655 457061
rect 302049 457058 302115 457061
rect 301589 457056 302115 457058
rect 301589 457000 301594 457056
rect 301650 457000 302054 457056
rect 302110 457000 302115 457056
rect 301589 456998 302115 457000
rect 301589 456995 301655 456998
rect 302049 456995 302115 456998
rect 301865 456922 301931 456925
rect 302141 456922 302207 456925
rect 301865 456920 302207 456922
rect 301865 456864 301870 456920
rect 301926 456864 302146 456920
rect 302202 456864 302207 456920
rect 301865 456862 302207 456864
rect 301865 456859 301931 456862
rect 302141 456859 302207 456862
rect 478086 456860 478092 456924
rect 478156 456922 478162 456924
rect 478873 456922 478939 456925
rect 478156 456920 478939 456922
rect 478156 456864 478878 456920
rect 478934 456864 478939 456920
rect 478156 456862 478939 456864
rect 478156 456860 478162 456862
rect 478873 456859 478939 456862
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 580758 418236 580764 418300
rect 580828 418298 580834 418300
rect 583520 418298 584960 418388
rect 580828 418238 584960 418298
rect 580828 418236 580834 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 583520 404820 584960 405060
rect 2773 398850 2839 398853
rect 3509 398850 3575 398853
rect 2773 398848 3575 398850
rect 2773 398792 2778 398848
rect 2834 398792 3514 398848
rect 3570 398792 3575 398848
rect 2773 398790 3575 398792
rect 2773 398787 2839 398790
rect 3509 398787 3575 398790
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580441 378450 580507 378453
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580441 378448 584960 378450
rect 580441 378392 580446 378448
rect 580502 378392 580906 378448
rect 580962 378392 584960 378448
rect 580441 378390 584960 378392
rect 580441 378387 580507 378390
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 674 358458
rect -960 358322 480 358398
rect 614 358322 674 358398
rect -960 358308 674 358322
rect 246 358262 674 358308
rect 246 357778 306 358262
rect 246 357718 6930 357778
rect 6870 357506 6930 357718
rect 21214 357506 21220 357508
rect 6870 357446 21220 357506
rect 21214 357444 21220 357446
rect 21284 357444 21290 357508
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect 197353 332754 197419 332757
rect 198590 332754 198596 332756
rect 197353 332752 198596 332754
rect 197353 332696 197358 332752
rect 197414 332696 198596 332752
rect 197353 332694 198596 332696
rect 197353 332691 197419 332694
rect 198590 332692 198596 332694
rect 198660 332692 198666 332756
rect -960 332196 480 332436
rect 23054 332420 23060 332484
rect 23124 332482 23130 332484
rect 69105 332482 69171 332485
rect 23124 332480 69171 332482
rect 23124 332424 69110 332480
rect 69166 332424 69171 332480
rect 23124 332422 69171 332424
rect 23124 332420 23130 332422
rect 69105 332419 69171 332422
rect 300301 332482 300367 332485
rect 302734 332482 302740 332484
rect 300301 332480 302740 332482
rect 300301 332424 300306 332480
rect 300362 332424 302740 332480
rect 300301 332422 302740 332424
rect 300301 332419 300367 332422
rect 302734 332420 302740 332422
rect 302804 332482 302810 332484
rect 302877 332482 302943 332485
rect 302804 332480 302943 332482
rect 302804 332424 302882 332480
rect 302938 332424 302943 332480
rect 302804 332422 302943 332424
rect 302804 332420 302810 332422
rect 302877 332419 302943 332422
rect 303061 332482 303127 332485
rect 580625 332482 580691 332485
rect 303061 332480 580691 332482
rect 303061 332424 303066 332480
rect 303122 332424 580630 332480
rect 580686 332424 580691 332480
rect 303061 332422 580691 332424
rect 303061 332419 303127 332422
rect 580625 332419 580691 332422
rect 23238 332284 23244 332348
rect 23308 332346 23314 332348
rect 57513 332346 57579 332349
rect 23308 332344 57579 332346
rect 23308 332288 57518 332344
rect 57574 332288 57579 332344
rect 23308 332286 57579 332288
rect 23308 332284 23314 332286
rect 57513 332283 57579 332286
rect 189533 331938 189599 331941
rect 233877 331938 233943 331941
rect 189533 331936 233943 331938
rect 189533 331880 189538 331936
rect 189594 331880 233882 331936
rect 233938 331880 233943 331936
rect 189533 331878 233943 331880
rect 189533 331875 189599 331878
rect 233877 331875 233943 331878
rect 96429 331802 96495 331805
rect 258073 331802 258139 331805
rect 96429 331800 258139 331802
rect 96429 331744 96434 331800
rect 96490 331744 258078 331800
rect 258134 331744 258139 331800
rect 96429 331742 258139 331744
rect 96429 331739 96495 331742
rect 258073 331739 258139 331742
rect 266353 331802 266419 331805
rect 372613 331802 372679 331805
rect 266353 331800 372679 331802
rect 266353 331744 266358 331800
rect 266414 331744 372618 331800
rect 372674 331744 372679 331800
rect 266353 331742 372679 331744
rect 266353 331739 266419 331742
rect 372613 331739 372679 331742
rect 469213 331802 469279 331805
rect 480253 331802 480319 331805
rect 469213 331800 480319 331802
rect 469213 331744 469218 331800
rect 469274 331744 480258 331800
rect 480314 331744 480319 331800
rect 469213 331742 480319 331744
rect 469213 331739 469279 331742
rect 480253 331739 480319 331742
rect 476941 331258 477007 331261
rect 477534 331258 477540 331260
rect 476941 331256 477540 331258
rect 476941 331200 476946 331256
rect 477002 331200 477540 331256
rect 476941 331198 477540 331200
rect 476941 331195 477007 331198
rect 477534 331196 477540 331198
rect 477604 331196 477610 331260
rect 477493 329762 477559 329765
rect 478086 329762 478092 329764
rect 477493 329760 478092 329762
rect 477493 329704 477498 329760
rect 477554 329704 478092 329760
rect 477493 329702 478092 329704
rect 477493 329699 477559 329702
rect 478086 329700 478092 329702
rect 478156 329762 478162 329764
rect 479057 329762 479123 329765
rect 478156 329760 479123 329762
rect 478156 329704 479062 329760
rect 479118 329704 479123 329760
rect 478156 329702 479123 329704
rect 478156 329700 478162 329702
rect 479057 329699 479123 329702
rect 583520 325124 584960 325364
rect -960 319290 480 319380
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 200062 315964 200068 316028
rect 200132 316026 200138 316028
rect 200481 316026 200547 316029
rect 200132 316024 200547 316026
rect 200132 315968 200486 316024
rect 200542 315968 200547 316024
rect 200132 315966 200547 315968
rect 200132 315964 200138 315966
rect 200481 315963 200547 315966
rect 299974 315828 299980 315892
rect 300044 315890 300050 315892
rect 300577 315890 300643 315893
rect 300044 315888 300643 315890
rect 300044 315832 300582 315888
rect 300638 315832 300643 315888
rect 300044 315830 300643 315832
rect 300044 315828 300050 315830
rect 300577 315827 300643 315830
rect 303521 315620 303587 315621
rect 303470 315556 303476 315620
rect 303540 315618 303587 315620
rect 303540 315616 303632 315618
rect 303582 315560 303632 315616
rect 303540 315558 303632 315560
rect 303540 315556 303587 315558
rect 303521 315555 303587 315556
rect 299473 315346 299539 315349
rect 387793 315346 387859 315349
rect 299473 315344 387859 315346
rect 299473 315288 299478 315344
rect 299534 315288 387798 315344
rect 387854 315288 387859 315344
rect 299473 315286 387859 315288
rect 299473 315283 299539 315286
rect 387793 315283 387859 315286
rect 476113 315346 476179 315349
rect 477350 315346 477356 315348
rect 476113 315344 477356 315346
rect 476113 315288 476118 315344
rect 476174 315288 477356 315344
rect 476113 315286 477356 315288
rect 476113 315283 476179 315286
rect 477350 315284 477356 315286
rect 477420 315346 477426 315348
rect 483013 315346 483079 315349
rect 477420 315344 483079 315346
rect 477420 315288 483018 315344
rect 483074 315288 483079 315344
rect 477420 315286 483079 315288
rect 477420 315284 477426 315286
rect 483013 315283 483079 315286
rect 299289 314802 299355 314805
rect 299974 314802 299980 314804
rect 299289 314800 299980 314802
rect 299289 314744 299294 314800
rect 299350 314744 299980 314800
rect 299289 314742 299980 314744
rect 299289 314739 299355 314742
rect 299974 314740 299980 314742
rect 300044 314740 300050 314804
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 477534 275300 477540 275364
rect 477604 275362 477610 275364
rect 477902 275362 477908 275364
rect 477604 275302 477908 275362
rect 477604 275300 477610 275302
rect 477902 275300 477908 275302
rect 477972 275300 477978 275364
rect 583520 272084 584960 272324
rect -960 267202 480 267292
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 3693 214978 3759 214981
rect -960 214976 3759 214978
rect -960 214920 3698 214976
rect 3754 214920 3759 214976
rect -960 214918 3759 214920
rect -960 214828 480 214918
rect 3693 214915 3759 214918
rect 480621 207634 480687 207637
rect 481173 207634 481239 207637
rect 451230 207632 481239 207634
rect 451230 207576 480626 207632
rect 480682 207576 481178 207632
rect 481234 207576 481239 207632
rect 451230 207574 481239 207576
rect 451230 207090 451290 207574
rect 480621 207571 480687 207574
rect 481173 207571 481239 207574
rect 442398 207030 451290 207090
rect 442398 206685 442458 207030
rect 442349 206680 442458 206685
rect 442349 206624 442354 206680
rect 442410 206624 442458 206680
rect 442349 206622 442458 206624
rect 442349 206619 442415 206622
rect 19558 205668 19564 205732
rect 19628 205730 19634 205732
rect 20345 205730 20411 205733
rect 19628 205728 20411 205730
rect 19628 205672 20350 205728
rect 20406 205672 20411 205728
rect 19628 205670 20411 205672
rect 19628 205668 19634 205670
rect 20345 205667 20411 205670
rect 299974 205668 299980 205732
rect 300044 205730 300050 205732
rect 300209 205730 300275 205733
rect 300044 205728 300275 205730
rect 300044 205672 300214 205728
rect 300270 205672 300275 205728
rect 300044 205670 300275 205672
rect 300044 205668 300050 205670
rect 300209 205667 300275 205670
rect 476113 205730 476179 205733
rect 477350 205730 477356 205732
rect 476113 205728 477356 205730
rect 476113 205672 476118 205728
rect 476174 205672 477356 205728
rect 476113 205670 477356 205672
rect 476113 205667 476179 205670
rect 477350 205668 477356 205670
rect 477420 205668 477426 205732
rect 583520 205580 584960 205820
rect 183461 204370 183527 204373
rect 197997 204370 198063 204373
rect 183461 204368 198063 204370
rect 183461 204312 183466 204368
rect 183522 204312 198002 204368
rect 198058 204312 198063 204368
rect 183461 204310 198063 204312
rect 183461 204307 183527 204310
rect 197997 204307 198063 204310
rect 303470 204308 303476 204372
rect 303540 204370 303546 204372
rect 337837 204370 337903 204373
rect 303540 204368 337903 204370
rect 303540 204312 337842 204368
rect 337898 204312 337903 204368
rect 303540 204310 337903 204312
rect 303540 204308 303546 204310
rect 337837 204307 337903 204310
rect 18873 204234 18939 204237
rect 88425 204234 88491 204237
rect 18873 204232 88491 204234
rect 18873 204176 18878 204232
rect 18934 204176 88430 204232
rect 88486 204176 88491 204232
rect 18873 204174 88491 204176
rect 18873 204171 18939 204174
rect 88425 204171 88491 204174
rect 115749 204234 115815 204237
rect 202965 204234 203031 204237
rect 115749 204232 203031 204234
rect 115749 204176 115754 204232
rect 115810 204176 202970 204232
rect 203026 204176 203031 204232
rect 115749 204174 203031 204176
rect 115749 204171 115815 204174
rect 202965 204171 203031 204174
rect 300485 204234 300551 204237
rect 300761 204234 300827 204237
rect 300485 204232 302618 204234
rect 300485 204176 300490 204232
rect 300546 204176 300766 204232
rect 300822 204176 302618 204232
rect 300485 204174 302618 204176
rect 300485 204171 300551 204174
rect 300761 204171 300827 204174
rect 4889 204098 4955 204101
rect 26601 204098 26667 204101
rect 4889 204096 26667 204098
rect 4889 204040 4894 204096
rect 4950 204040 26606 204096
rect 26662 204040 26667 204096
rect 4889 204038 26667 204040
rect 302558 204098 302618 204174
rect 302734 204172 302740 204236
rect 302804 204234 302810 204236
rect 303470 204234 303476 204236
rect 302804 204174 303476 204234
rect 302804 204172 302810 204174
rect 303470 204172 303476 204174
rect 303540 204234 303546 204236
rect 364885 204234 364951 204237
rect 303540 204232 364951 204234
rect 303540 204176 364890 204232
rect 364946 204176 364951 204232
rect 303540 204174 364951 204176
rect 303540 204172 303546 204174
rect 364885 204171 364951 204174
rect 430573 204234 430639 204237
rect 475377 204234 475443 204237
rect 477953 204234 478019 204237
rect 478321 204234 478387 204237
rect 430573 204232 475443 204234
rect 430573 204176 430578 204232
rect 430634 204176 475382 204232
rect 475438 204176 475443 204232
rect 430573 204174 475443 204176
rect 430573 204171 430639 204174
rect 475377 204171 475443 204174
rect 475518 204232 478387 204234
rect 475518 204176 477958 204232
rect 478014 204176 478326 204232
rect 478382 204176 478387 204232
rect 475518 204174 478387 204176
rect 345565 204098 345631 204101
rect 302558 204096 345631 204098
rect 302558 204040 345570 204096
rect 345626 204040 345631 204096
rect 302558 204038 345631 204040
rect 4889 204035 4955 204038
rect 26601 204035 26667 204038
rect 345565 204035 345631 204038
rect 446029 204098 446095 204101
rect 475518 204098 475578 204174
rect 477953 204171 478019 204174
rect 478321 204171 478387 204174
rect 446029 204096 475578 204098
rect 446029 204040 446034 204096
rect 446090 204040 475578 204096
rect 446029 204038 475578 204040
rect 446029 204035 446095 204038
rect 195881 203962 195947 203965
rect 200389 203962 200455 203965
rect 200573 203962 200639 203965
rect 195881 203960 200639 203962
rect 195881 203904 195886 203960
rect 195942 203904 200394 203960
rect 200450 203904 200578 203960
rect 200634 203904 200639 203960
rect 195881 203902 200639 203904
rect 195881 203899 195947 203902
rect 200389 203899 200455 203902
rect 200573 203899 200639 203902
rect 475377 203962 475443 203965
rect 478413 203962 478479 203965
rect 475377 203960 478479 203962
rect 475377 203904 475382 203960
rect 475438 203904 478418 203960
rect 478474 203904 478479 203960
rect 475377 203902 478479 203904
rect 475377 203899 475443 203902
rect 478413 203899 478479 203902
rect 476021 203826 476087 203829
rect 481909 203826 481975 203829
rect 476021 203824 481975 203826
rect 476021 203768 476026 203824
rect 476082 203768 481914 203824
rect 481970 203768 481975 203824
rect 476021 203766 481975 203768
rect 476021 203763 476087 203766
rect 481909 203763 481975 203766
rect 22829 203554 22895 203557
rect 30465 203554 30531 203557
rect 22829 203552 30531 203554
rect 22829 203496 22834 203552
rect 22890 203496 30470 203552
rect 30526 203496 30531 203552
rect 22829 203494 30531 203496
rect 22829 203491 22895 203494
rect 30465 203491 30531 203494
rect 179873 203554 179939 203557
rect 198917 203554 198983 203557
rect 179873 203552 198983 203554
rect 179873 203496 179878 203552
rect 179934 203496 198922 203552
rect 198978 203496 198983 203552
rect 179873 203494 198983 203496
rect 179873 203491 179939 203494
rect 198917 203491 198983 203494
rect 197813 203012 197879 203013
rect 23054 202948 23060 203012
rect 23124 202948 23130 203012
rect 197813 203008 197860 203012
rect 197924 203010 197930 203012
rect 197813 202952 197818 203008
rect 197813 202948 197860 202952
rect 197924 202950 197970 203010
rect 197924 202948 197930 202950
rect 22369 202874 22435 202877
rect 23062 202874 23122 202948
rect 197813 202947 197879 202948
rect 69105 202874 69171 202877
rect 22369 202872 69171 202874
rect 22369 202816 22374 202872
rect 22430 202816 69110 202872
rect 69166 202816 69171 202872
rect 22369 202814 69171 202816
rect 22369 202811 22435 202814
rect 69105 202811 69171 202814
rect 477493 202874 477559 202877
rect 477718 202874 477724 202876
rect 477493 202872 477724 202874
rect 477493 202816 477498 202872
rect 477554 202816 477724 202872
rect 477493 202814 477724 202816
rect 477493 202811 477559 202814
rect 477718 202812 477724 202814
rect 477788 202812 477794 202876
rect 23238 202676 23244 202740
rect 23308 202738 23314 202740
rect 57513 202738 57579 202741
rect 23308 202736 57579 202738
rect 23308 202680 57518 202736
rect 57574 202680 57579 202736
rect 23308 202678 57579 202680
rect 23308 202676 23314 202678
rect 57513 202675 57579 202678
rect -960 201772 480 202012
rect 198590 201316 198596 201380
rect 198660 201378 198666 201380
rect 198733 201378 198799 201381
rect 198660 201376 198799 201378
rect 198660 201320 198738 201376
rect 198794 201320 198799 201376
rect 198660 201318 198799 201320
rect 198660 201316 198666 201318
rect 198733 201315 198799 201318
rect 583520 192388 584960 192628
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 477534 149908 477540 149972
rect 477604 149970 477610 149972
rect 480621 149970 480687 149973
rect 477604 149968 480687 149970
rect 477604 149912 480626 149968
rect 480682 149912 480687 149968
rect 477604 149910 480687 149912
rect 477604 149908 477610 149910
rect 480621 149907 480687 149910
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 20897 110394 20963 110397
rect 21541 110394 21607 110397
rect 20897 110392 21607 110394
rect 20897 110336 20902 110392
rect 20958 110336 21546 110392
rect 21602 110336 21607 110392
rect 20897 110334 21607 110336
rect 20897 110331 20963 110334
rect 21541 110331 21607 110334
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 477534 81908 477540 81972
rect 477604 81970 477610 81972
rect 477902 81970 477908 81972
rect 477604 81910 477908 81970
rect 477604 81908 477610 81910
rect 477902 81908 477908 81910
rect 477972 81908 477978 81972
rect 579613 78434 579679 78437
rect 580758 78434 580764 78436
rect 579613 78432 580764 78434
rect 579613 78376 579618 78432
rect 579674 78376 580764 78432
rect 579613 78374 580764 78376
rect 579613 78371 579679 78374
rect 580758 78372 580764 78374
rect 580828 78372 580834 78436
rect 393313 78162 393379 78165
rect 477718 78162 477724 78164
rect 393313 78160 477724 78162
rect 393313 78104 393318 78160
rect 393374 78104 477724 78160
rect 393313 78102 477724 78104
rect 393313 78099 393379 78102
rect 477718 78100 477724 78102
rect 477788 78100 477794 78164
rect 390553 78026 390619 78029
rect 478822 78026 478828 78028
rect 390553 78024 478828 78026
rect 390553 77968 390558 78024
rect 390614 77968 478828 78024
rect 390553 77966 478828 77968
rect 390553 77963 390619 77966
rect 478822 77964 478828 77966
rect 478892 77964 478898 78028
rect 303286 77828 303292 77892
rect 303356 77890 303362 77892
rect 336733 77890 336799 77893
rect 337469 77890 337535 77893
rect 303356 77888 337535 77890
rect 303356 77832 336738 77888
rect 336794 77832 337474 77888
rect 337530 77832 337535 77888
rect 303356 77830 337535 77832
rect 303356 77828 303362 77830
rect 336733 77827 336799 77830
rect 337469 77827 337535 77830
rect 389173 77890 389239 77893
rect 481582 77890 481588 77892
rect 389173 77888 481588 77890
rect 389173 77832 389178 77888
rect 389234 77832 481588 77888
rect 389173 77830 481588 77832
rect 389173 77827 389239 77830
rect 481582 77828 481588 77830
rect 481652 77828 481658 77892
rect 303337 77346 303403 77349
rect 311157 77346 311223 77349
rect 303337 77344 311223 77346
rect 303337 77288 303342 77344
rect 303398 77288 311162 77344
rect 311218 77288 311223 77344
rect 303337 77286 311223 77288
rect 303337 77283 303403 77286
rect 311157 77283 311223 77286
rect 480253 77348 480319 77349
rect 480253 77344 480300 77348
rect 480364 77346 480370 77348
rect 480253 77288 480258 77344
rect 480253 77284 480300 77288
rect 480364 77286 480410 77346
rect 480364 77284 480370 77286
rect 480253 77283 480319 77284
rect 19558 75788 19564 75852
rect 19628 75850 19634 75852
rect 81249 75850 81315 75853
rect 19628 75848 81315 75850
rect 19628 75792 81254 75848
rect 81310 75792 81315 75848
rect 19628 75790 81315 75792
rect 19628 75788 19634 75790
rect 81249 75787 81315 75790
rect 4797 75714 4863 75717
rect 26601 75714 26667 75717
rect 4797 75712 26667 75714
rect 4797 75656 4802 75712
rect 4858 75656 26606 75712
rect 26662 75656 26667 75712
rect 4797 75654 26667 75656
rect 4797 75651 4863 75654
rect 26601 75651 26667 75654
rect 50337 75170 50403 75173
rect 98494 75170 98500 75172
rect 50337 75168 98500 75170
rect 50337 75112 50342 75168
rect 50398 75112 98500 75168
rect 50337 75110 98500 75112
rect 50337 75107 50403 75110
rect 98494 75108 98500 75110
rect 98564 75108 98570 75172
rect 303470 75108 303476 75172
rect 303540 75170 303546 75172
rect 336825 75170 336891 75173
rect 303540 75168 336891 75170
rect 303540 75112 336830 75168
rect 336886 75112 336891 75168
rect 303540 75110 336891 75112
rect 303540 75108 303546 75110
rect 336825 75107 336891 75110
rect 373993 75170 374059 75173
rect 481633 75170 481699 75173
rect 373993 75168 481699 75170
rect 373993 75112 373998 75168
rect 374054 75112 481638 75168
rect 481694 75112 481699 75168
rect 373993 75110 481699 75112
rect 373993 75107 374059 75110
rect 481633 75107 481699 75110
rect 23238 74428 23244 74492
rect 23308 74490 23314 74492
rect 57237 74490 57303 74493
rect 23308 74488 57303 74490
rect 23308 74432 57242 74488
rect 57298 74432 57303 74488
rect 23308 74430 57303 74432
rect 23308 74428 23314 74430
rect 57237 74427 57303 74430
rect 395797 74490 395863 74493
rect 484485 74490 484551 74493
rect 395797 74488 484551 74490
rect 395797 74432 395802 74488
rect 395858 74432 484490 74488
rect 484546 74432 484551 74488
rect 395797 74430 484551 74432
rect 395797 74427 395863 74430
rect 484485 74427 484551 74430
rect 392577 74354 392643 74357
rect 480621 74354 480687 74357
rect 392577 74352 480687 74354
rect 392577 74296 392582 74352
rect 392638 74296 480626 74352
rect 480682 74296 480687 74352
rect 392577 74294 480687 74296
rect 392577 74291 392643 74294
rect 480621 74291 480687 74294
rect 399477 73130 399543 73133
rect 476614 73130 476620 73132
rect 399477 73128 476620 73130
rect 399477 73072 399482 73128
rect 399538 73072 476620 73128
rect 399477 73070 476620 73072
rect 399477 73067 399543 73070
rect 476614 73068 476620 73070
rect 476684 73068 476690 73132
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 3785 71634 3851 71637
rect -960 71632 3851 71634
rect -960 71576 3790 71632
rect 3846 71576 3851 71632
rect -960 71574 3851 71576
rect -960 71484 480 71574
rect 3785 71571 3851 71574
rect 300025 64836 300091 64837
rect 299974 64834 299980 64836
rect 299934 64774 299980 64834
rect 300044 64832 300091 64836
rect 300086 64776 300091 64832
rect 299974 64772 299980 64774
rect 300044 64772 300091 64776
rect 300025 64771 300091 64772
rect 197813 63476 197879 63477
rect 197813 63472 197860 63476
rect 197924 63474 197930 63476
rect 197813 63416 197818 63472
rect 197813 63412 197860 63416
rect 197924 63414 197970 63474
rect 197924 63412 197930 63414
rect 197813 63411 197879 63412
rect 57053 61570 57119 61573
rect 57053 61568 60106 61570
rect 57053 61512 57058 61568
rect 57114 61512 60106 61568
rect 57053 61510 60106 61512
rect 57053 61507 57119 61510
rect 60046 61064 60106 61510
rect 99790 60754 99850 61336
rect 102726 60754 102732 60756
rect 99790 60694 102732 60754
rect 102726 60692 102732 60694
rect 102796 60692 102802 60756
rect 99790 59666 99850 60248
rect 103053 59666 103119 59669
rect 99790 59664 103119 59666
rect 99790 59608 103058 59664
rect 103114 59608 103119 59664
rect 99790 59606 103119 59608
rect 103053 59603 103119 59606
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 99790 58578 99850 59160
rect 99966 58652 99972 58716
rect 100036 58714 100042 58716
rect 100036 58654 103530 58714
rect 100036 58652 100042 58654
rect 102777 58578 102843 58581
rect 99790 58576 102843 58578
rect 99790 58520 102782 58576
rect 102838 58520 102843 58576
rect 99790 58518 102843 58520
rect 103470 58578 103530 58654
rect 346761 58578 346827 58581
rect 103470 58576 346827 58578
rect 103470 58520 346766 58576
rect 346822 58520 346827 58576
rect 103470 58518 346827 58520
rect 102777 58515 102843 58518
rect 346761 58515 346827 58518
rect 99790 58034 99850 58072
rect 102910 58034 102916 58036
rect 99790 57974 102916 58034
rect 102910 57972 102916 57974
rect 102980 57972 102986 58036
rect 298737 57354 298803 57357
rect 371969 57354 372035 57357
rect 298737 57352 372035 57354
rect 298737 57296 298742 57352
rect 298798 57296 371974 57352
rect 372030 57296 372035 57352
rect 298737 57294 372035 57296
rect 298737 57291 298803 57294
rect 371969 57291 372035 57294
rect 298870 57156 298876 57220
rect 298940 57218 298946 57220
rect 388529 57218 388595 57221
rect 298940 57216 388595 57218
rect 298940 57160 388534 57216
rect 388590 57160 388595 57216
rect 298940 57158 388595 57160
rect 298940 57156 298946 57158
rect 388529 57155 388595 57158
rect 99790 56674 99850 56984
rect 102593 56674 102659 56677
rect 99790 56672 102659 56674
rect 99790 56616 102598 56672
rect 102654 56616 102659 56672
rect 99790 56614 102659 56616
rect 102593 56611 102659 56614
rect 57513 56402 57579 56405
rect 57513 56400 60106 56402
rect 57513 56344 57518 56400
rect 57574 56344 60106 56400
rect 57513 56342 60106 56344
rect 57513 56339 57579 56342
rect 60046 56168 60106 56342
rect 99790 55586 99850 55896
rect 102961 55586 103027 55589
rect 99790 55584 103027 55586
rect 99790 55528 102966 55584
rect 103022 55528 103027 55584
rect 99790 55526 103027 55528
rect 102961 55523 103027 55526
rect 99790 54226 99850 54808
rect 102225 54226 102291 54229
rect 99790 54224 102291 54226
rect 99790 54168 102230 54224
rect 102286 54168 102291 54224
rect 99790 54166 102291 54168
rect 102225 54163 102291 54166
rect 99790 53546 99850 53720
rect 102133 53546 102199 53549
rect 99790 53544 102199 53546
rect 99790 53488 102138 53544
rect 102194 53488 102199 53544
rect 99790 53486 102199 53488
rect 102133 53483 102199 53486
rect 99790 52594 99850 52632
rect 102133 52594 102199 52597
rect 99790 52592 102199 52594
rect 99790 52536 102138 52592
rect 102194 52536 102199 52592
rect 99790 52534 102199 52536
rect 102133 52531 102199 52534
rect 57053 51778 57119 51781
rect 57053 51776 60106 51778
rect 57053 51720 57058 51776
rect 57114 51720 60106 51776
rect 57053 51718 60106 51720
rect 57053 51715 57119 51718
rect 60046 51272 60106 51718
rect 99790 51098 99850 51544
rect 102726 51444 102732 51508
rect 102796 51506 102802 51508
rect 199334 51506 199394 52088
rect 102796 51446 199394 51506
rect 102796 51444 102802 51446
rect 195973 51370 196039 51373
rect 195973 51368 199394 51370
rect 195973 51312 195978 51368
rect 196034 51312 199394 51368
rect 195973 51310 199394 51312
rect 195973 51307 196039 51310
rect 199334 51272 199394 51310
rect 103237 51098 103303 51101
rect 99790 51096 103303 51098
rect 99790 51040 103242 51096
rect 103298 51040 103303 51096
rect 99790 51038 103303 51040
rect 103237 51035 103303 51038
rect 195973 50962 196039 50965
rect 195973 50960 199394 50962
rect 195973 50904 195978 50960
rect 196034 50904 199394 50960
rect 195973 50902 199394 50904
rect 195973 50899 196039 50902
rect 199334 50456 199394 50902
rect 99790 49874 99850 50456
rect 103053 49874 103119 49877
rect 99790 49872 103119 49874
rect 99790 49816 103058 49872
rect 103114 49816 103119 49872
rect 99790 49814 103119 49816
rect 103053 49811 103119 49814
rect 199334 49602 199394 49640
rect 180750 49542 199394 49602
rect 99790 48786 99850 49368
rect 103421 48786 103487 48789
rect 99790 48784 103487 48786
rect 99790 48728 103426 48784
rect 103482 48728 103487 48784
rect 99790 48726 103487 48728
rect 103421 48723 103487 48726
rect 102910 48588 102916 48652
rect 102980 48650 102986 48652
rect 180750 48650 180810 49542
rect 195973 49466 196039 49469
rect 195973 49464 199394 49466
rect 195973 49408 195978 49464
rect 196034 49408 199394 49464
rect 195973 49406 199394 49408
rect 195973 49403 196039 49406
rect 199334 48824 199394 49406
rect 102980 48590 180810 48650
rect 102980 48588 102986 48590
rect 99790 47698 99850 48280
rect 195973 48242 196039 48245
rect 195973 48240 199394 48242
rect 195973 48184 195978 48240
rect 196034 48184 199394 48240
rect 195973 48182 199394 48184
rect 195973 48179 196039 48182
rect 199334 48008 199394 48182
rect 102726 47698 102732 47700
rect 99790 47638 102732 47698
rect 102726 47636 102732 47638
rect 102796 47636 102802 47700
rect 196065 47698 196131 47701
rect 196065 47696 199394 47698
rect 196065 47640 196070 47696
rect 196126 47640 199394 47696
rect 196065 47638 199394 47640
rect 196065 47635 196131 47638
rect 199334 47192 199394 47638
rect 99790 47018 99850 47192
rect 102685 47018 102751 47021
rect 99790 47016 102751 47018
rect 99790 46960 102690 47016
rect 102746 46960 102751 47016
rect 99790 46958 102751 46960
rect 102685 46955 102751 46958
rect 57513 46882 57579 46885
rect 195973 46882 196039 46885
rect 57513 46880 60106 46882
rect 57513 46824 57518 46880
rect 57574 46824 60106 46880
rect 57513 46822 60106 46824
rect 57513 46819 57579 46822
rect 60046 46376 60106 46822
rect 195973 46880 199394 46882
rect 195973 46824 195978 46880
rect 196034 46824 199394 46880
rect 195973 46822 199394 46824
rect 195973 46819 196039 46822
rect 199334 46376 199394 46822
rect 196157 46202 196223 46205
rect 196157 46200 199394 46202
rect 196157 46144 196162 46200
rect 196218 46144 199394 46200
rect 583520 46188 584960 46428
rect 196157 46142 199394 46144
rect 196157 46139 196223 46142
rect 99790 45794 99850 46104
rect 102777 45794 102843 45797
rect 99790 45792 102843 45794
rect 99790 45736 102782 45792
rect 102838 45736 102843 45792
rect 99790 45734 102843 45736
rect 102777 45731 102843 45734
rect -960 45522 480 45612
rect 199334 45560 199394 46142
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 195973 45250 196039 45253
rect 195973 45248 199394 45250
rect 195973 45192 195978 45248
rect 196034 45192 199394 45248
rect 195973 45190 199394 45192
rect 195973 45187 196039 45190
rect 99790 44434 99850 45016
rect 199334 44744 199394 45190
rect 102501 44434 102567 44437
rect 99790 44432 102567 44434
rect 99790 44376 102506 44432
rect 102562 44376 102567 44432
rect 99790 44374 102567 44376
rect 102501 44371 102567 44374
rect 195973 44026 196039 44029
rect 195973 44024 199394 44026
rect 195973 43968 195978 44024
rect 196034 43968 199394 44024
rect 195973 43966 199394 43968
rect 195973 43963 196039 43966
rect 199334 43928 199394 43966
rect 99790 43346 99850 43928
rect 196065 43618 196131 43621
rect 196065 43616 199394 43618
rect 196065 43560 196070 43616
rect 196126 43560 199394 43616
rect 196065 43558 199394 43560
rect 196065 43555 196131 43558
rect 102317 43346 102383 43349
rect 99790 43344 102383 43346
rect 99790 43288 102322 43344
rect 102378 43288 102383 43344
rect 99790 43286 102383 43288
rect 102317 43283 102383 43286
rect 199334 43112 199394 43558
rect 102409 42938 102475 42941
rect 99790 42936 102475 42938
rect 99790 42880 102414 42936
rect 102470 42880 102475 42936
rect 99790 42878 102475 42880
rect 99790 42840 99850 42878
rect 102409 42875 102475 42878
rect 57145 42122 57211 42125
rect 57145 42120 60106 42122
rect 57145 42064 57150 42120
rect 57206 42064 60106 42120
rect 57145 42062 60106 42064
rect 57145 42059 57211 42062
rect 60046 41480 60106 42062
rect 99790 41442 99850 41752
rect 102726 41652 102732 41716
rect 102796 41714 102802 41716
rect 199334 41714 199394 42296
rect 102796 41654 199394 41714
rect 102796 41652 102802 41654
rect 195973 41578 196039 41581
rect 195973 41576 199394 41578
rect 195973 41520 195978 41576
rect 196034 41520 199394 41576
rect 195973 41518 199394 41520
rect 195973 41515 196039 41518
rect 199334 41480 199394 41518
rect 102133 41442 102199 41445
rect 99790 41440 102199 41442
rect 99790 41384 102138 41440
rect 102194 41384 102199 41440
rect 99790 41382 102199 41384
rect 102133 41379 102199 41382
rect 195973 41170 196039 41173
rect 195973 41168 199394 41170
rect 195973 41112 195978 41168
rect 196034 41112 199394 41168
rect 195973 41110 199394 41112
rect 195973 41107 196039 41110
rect 199334 40664 199394 41110
rect 99790 40082 99850 40664
rect 102225 40082 102291 40085
rect 99790 40080 102291 40082
rect 99790 40024 102230 40080
rect 102286 40024 102291 40080
rect 99790 40022 102291 40024
rect 102225 40019 102291 40022
rect 195973 39946 196039 39949
rect 195973 39944 199394 39946
rect 195973 39888 195978 39944
rect 196034 39888 199394 39944
rect 195973 39886 199394 39888
rect 195973 39883 196039 39886
rect 199334 39848 199394 39886
rect 99790 38994 99850 39576
rect 196065 39538 196131 39541
rect 196065 39536 199394 39538
rect 196065 39480 196070 39536
rect 196126 39480 199394 39536
rect 196065 39478 199394 39480
rect 196065 39475 196131 39478
rect 199334 39032 199394 39478
rect 102869 38994 102935 38997
rect 99790 38992 102935 38994
rect 99790 38936 102874 38992
rect 102930 38936 102935 38992
rect 99790 38934 102935 38936
rect 102869 38931 102935 38934
rect 99790 37906 99850 38488
rect 195973 38450 196039 38453
rect 195973 38448 199394 38450
rect 195973 38392 195978 38448
rect 196034 38392 199394 38448
rect 195973 38390 199394 38392
rect 195973 38387 196039 38390
rect 199334 38216 199394 38390
rect 196065 38042 196131 38045
rect 196065 38040 199394 38042
rect 196065 37984 196070 38040
rect 196126 37984 199394 38040
rect 196065 37982 199394 37984
rect 196065 37979 196131 37982
rect 102133 37906 102199 37909
rect 99790 37904 102199 37906
rect 99790 37848 102138 37904
rect 102194 37848 102199 37904
rect 99790 37846 102199 37848
rect 102133 37843 102199 37846
rect 199334 37400 199394 37982
rect 99790 37362 99850 37400
rect 102593 37362 102659 37365
rect 99790 37360 102659 37362
rect 99790 37304 102598 37360
rect 102654 37304 102659 37360
rect 99790 37302 102659 37304
rect 102593 37299 102659 37302
rect 195973 37090 196039 37093
rect 195973 37088 199394 37090
rect 195973 37032 195978 37088
rect 196034 37032 199394 37088
rect 195973 37030 199394 37032
rect 195973 37027 196039 37030
rect 57053 36954 57119 36957
rect 57053 36952 60106 36954
rect 57053 36896 57058 36952
rect 57114 36896 60106 36952
rect 57053 36894 60106 36896
rect 57053 36891 57119 36894
rect 60046 36584 60106 36894
rect 199334 36584 199394 37030
rect 99790 36138 99850 36312
rect 102777 36138 102843 36141
rect 99790 36136 102843 36138
rect 99790 36080 102782 36136
rect 102838 36080 102843 36136
rect 99790 36078 102843 36080
rect 102777 36075 102843 36078
rect 195973 35866 196039 35869
rect 195973 35864 199394 35866
rect 195973 35808 195978 35864
rect 196034 35808 199394 35864
rect 195973 35806 199394 35808
rect 195973 35803 196039 35806
rect 199334 35768 199394 35806
rect 196065 35458 196131 35461
rect 196065 35456 199394 35458
rect 196065 35400 196070 35456
rect 196126 35400 199394 35456
rect 196065 35398 199394 35400
rect 196065 35395 196131 35398
rect 99790 34642 99850 35224
rect 199334 34952 199394 35398
rect 102133 34642 102199 34645
rect 99790 34640 102199 34642
rect 99790 34584 102138 34640
rect 102194 34584 102199 34640
rect 99790 34582 102199 34584
rect 102133 34579 102199 34582
rect 195973 34370 196039 34373
rect 195973 34368 199394 34370
rect 195973 34312 195978 34368
rect 196034 34312 199394 34368
rect 195973 34310 199394 34312
rect 195973 34307 196039 34310
rect 199334 34136 199394 34310
rect 99790 33554 99850 34136
rect 196065 33826 196131 33829
rect 196065 33824 199394 33826
rect 196065 33768 196070 33824
rect 196126 33768 199394 33824
rect 196065 33766 199394 33768
rect 196065 33763 196131 33766
rect 102317 33554 102383 33557
rect 99790 33552 102383 33554
rect 99790 33496 102322 33552
rect 102378 33496 102383 33552
rect 99790 33494 102383 33496
rect 102317 33491 102383 33494
rect 199334 33320 199394 33766
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect 99790 32466 99850 33048
rect 195973 33010 196039 33013
rect 195973 33008 199394 33010
rect 195973 32952 195978 33008
rect 196034 32952 199394 33008
rect 583520 32996 584960 33236
rect 195973 32950 199394 32952
rect 195973 32947 196039 32950
rect 199334 32504 199394 32950
rect 102133 32466 102199 32469
rect 99790 32464 102199 32466
rect 99790 32408 102138 32464
rect 102194 32408 102199 32464
rect 99790 32406 102199 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 102133 32403 102199 32406
rect 99790 31786 99850 31960
rect 102225 31786 102291 31789
rect 99790 31784 102291 31786
rect 99790 31728 102230 31784
rect 102286 31728 102291 31784
rect 99790 31726 102291 31728
rect 102225 31723 102291 31726
rect 57605 31650 57671 31653
rect 60046 31650 60106 31688
rect 57605 31648 60106 31650
rect 57605 31592 57610 31648
rect 57666 31592 60106 31648
rect 57605 31590 60106 31592
rect 195973 31650 196039 31653
rect 199334 31650 199394 31688
rect 195973 31648 199394 31650
rect 195973 31592 195978 31648
rect 196034 31592 199394 31648
rect 195973 31590 199394 31592
rect 57605 31587 57671 31590
rect 195973 31587 196039 31590
rect 196065 31242 196131 31245
rect 196065 31240 199394 31242
rect 196065 31184 196070 31240
rect 196126 31184 199394 31240
rect 196065 31182 199394 31184
rect 196065 31179 196131 31182
rect 199334 30872 199394 31182
rect 99790 30562 99850 30872
rect 102133 30562 102199 30565
rect 99790 30560 102199 30562
rect 99790 30504 102138 30560
rect 102194 30504 102199 30560
rect 99790 30502 102199 30504
rect 102133 30499 102199 30502
rect 195973 30290 196039 30293
rect 195973 30288 199394 30290
rect 195973 30232 195978 30288
rect 196034 30232 199394 30288
rect 195973 30230 199394 30232
rect 195973 30227 196039 30230
rect 199334 30056 199394 30230
rect 99790 29338 99850 29784
rect 196065 29746 196131 29749
rect 196065 29744 199394 29746
rect 196065 29688 196070 29744
rect 196126 29688 199394 29744
rect 196065 29686 199394 29688
rect 196065 29683 196131 29686
rect 102133 29338 102199 29341
rect 99790 29336 102199 29338
rect 99790 29280 102138 29336
rect 102194 29280 102199 29336
rect 99790 29278 102199 29280
rect 102133 29275 102199 29278
rect 199334 29240 199394 29686
rect 195973 28930 196039 28933
rect 195973 28928 199394 28930
rect 195973 28872 195978 28928
rect 196034 28872 199394 28928
rect 195973 28870 199394 28872
rect 195973 28867 196039 28870
rect 99790 28522 99850 28696
rect 102133 28522 102199 28525
rect 99790 28520 102199 28522
rect 99790 28464 102138 28520
rect 102194 28464 102199 28520
rect 99790 28462 102199 28464
rect 102133 28459 102199 28462
rect 199334 28424 199394 28870
rect 195973 28114 196039 28117
rect 195973 28112 199394 28114
rect 195973 28056 195978 28112
rect 196034 28056 199394 28112
rect 195973 28054 199394 28056
rect 195973 28051 196039 28054
rect 102133 27706 102199 27709
rect 99790 27704 102199 27706
rect 99790 27648 102138 27704
rect 102194 27648 102199 27704
rect 99790 27646 102199 27648
rect 99790 27608 99850 27646
rect 102133 27643 102199 27646
rect 199334 27608 199394 28054
rect 195973 27298 196039 27301
rect 195973 27296 199394 27298
rect 195973 27240 195978 27296
rect 196034 27240 199394 27296
rect 195973 27238 199394 27240
rect 195973 27235 196039 27238
rect 57237 27162 57303 27165
rect 57237 27160 60106 27162
rect 57237 27104 57242 27160
rect 57298 27104 60106 27160
rect 57237 27102 60106 27104
rect 57237 27099 57303 27102
rect 60046 26792 60106 27102
rect 199334 26792 199394 27238
rect 99790 26346 99850 26520
rect 102777 26346 102843 26349
rect 99790 26344 102843 26346
rect 99790 26288 102782 26344
rect 102838 26288 102843 26344
rect 99790 26286 102843 26288
rect 102777 26283 102843 26286
rect 195973 26210 196039 26213
rect 195973 26208 199394 26210
rect 195973 26152 195978 26208
rect 196034 26152 199394 26208
rect 195973 26150 199394 26152
rect 195973 26147 196039 26150
rect 199334 25976 199394 26150
rect 3366 22068 3372 22132
rect 3436 22130 3442 22132
rect 371693 22130 371759 22133
rect 3436 22128 371759 22130
rect 3436 22072 371698 22128
rect 371754 22072 371759 22128
rect 3436 22070 371759 22072
rect 3436 22068 3442 22070
rect 371693 22067 371759 22070
rect 21214 21932 21220 21996
rect 21284 21994 21290 21996
rect 357341 21994 357407 21997
rect 21284 21992 357407 21994
rect 21284 21936 357346 21992
rect 357402 21936 357407 21992
rect 21284 21934 357407 21936
rect 21284 21932 21290 21934
rect 357341 21931 357407 21934
rect 199326 21796 199332 21860
rect 199396 21858 199402 21860
rect 375281 21858 375347 21861
rect 199396 21856 375347 21858
rect 199396 21800 375286 21856
rect 375342 21800 375347 21856
rect 199396 21798 375347 21800
rect 199396 21796 199402 21798
rect 375281 21795 375347 21798
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 199332 700300 199396 700364
rect 479380 683164 479444 683228
rect 3372 607140 3436 607204
rect 3372 606052 3436 606116
rect 23244 585788 23308 585852
rect 480300 585788 480364 585852
rect 476620 585652 476684 585716
rect 481588 585108 481652 585172
rect 23060 582932 23124 582996
rect 199884 582932 199948 582996
rect 303476 582932 303540 582996
rect 197308 572052 197372 572116
rect 21956 571916 22020 571980
rect 298876 571916 298940 571980
rect 477540 533428 477604 533492
rect 299980 462164 300044 462228
rect 479380 460804 479444 460868
rect 197860 459308 197924 459372
rect 22876 458900 22940 458964
rect 23060 458764 23124 458828
rect 21956 458220 22020 458284
rect 22876 458220 22940 458284
rect 478828 458220 478892 458284
rect 23244 458084 23308 458148
rect 199884 458084 199948 458148
rect 303476 457948 303540 458012
rect 478092 456860 478156 456924
rect 580764 418236 580828 418300
rect 21220 357444 21284 357508
rect 198596 332692 198660 332756
rect 23060 332420 23124 332484
rect 302740 332420 302804 332484
rect 23244 332284 23308 332348
rect 477540 331196 477604 331260
rect 478092 329700 478156 329764
rect 200068 315964 200132 316028
rect 299980 315828 300044 315892
rect 303476 315616 303540 315620
rect 303476 315560 303526 315616
rect 303526 315560 303540 315616
rect 303476 315556 303540 315560
rect 477356 315284 477420 315348
rect 299980 314740 300044 314804
rect 477540 275300 477604 275364
rect 477908 275300 477972 275364
rect 19564 205668 19628 205732
rect 299980 205668 300044 205732
rect 477356 205668 477420 205732
rect 303476 204308 303540 204372
rect 302740 204172 302804 204236
rect 303476 204172 303540 204236
rect 23060 202948 23124 203012
rect 197860 203008 197924 203012
rect 197860 202952 197874 203008
rect 197874 202952 197924 203008
rect 197860 202948 197924 202952
rect 477724 202812 477788 202876
rect 23244 202676 23308 202740
rect 198596 201316 198660 201380
rect 477540 149908 477604 149972
rect 477540 81908 477604 81972
rect 477908 81908 477972 81972
rect 580764 78372 580828 78436
rect 477724 78100 477788 78164
rect 478828 77964 478892 78028
rect 303292 77828 303356 77892
rect 481588 77828 481652 77892
rect 480300 77344 480364 77348
rect 480300 77288 480314 77344
rect 480314 77288 480364 77344
rect 480300 77284 480364 77288
rect 19564 75788 19628 75852
rect 98500 75108 98564 75172
rect 303476 75108 303540 75172
rect 23244 74428 23308 74492
rect 476620 73068 476684 73132
rect 299980 64832 300044 64836
rect 299980 64776 300030 64832
rect 300030 64776 300044 64832
rect 299980 64772 300044 64776
rect 197860 63472 197924 63476
rect 197860 63416 197874 63472
rect 197874 63416 197924 63472
rect 197860 63412 197924 63416
rect 102732 60692 102796 60756
rect 99972 58652 100036 58716
rect 102916 57972 102980 58036
rect 298876 57156 298940 57220
rect 102732 51444 102796 51508
rect 102916 48588 102980 48652
rect 102732 47636 102796 47700
rect 102732 41652 102796 41716
rect 3372 22068 3436 22132
rect 21220 21932 21284 21996
rect 199332 21796 199396 21860
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 3371 607204 3437 607205
rect 3371 607140 3372 607204
rect 3436 607140 3437 607204
rect 3371 607139 3437 607140
rect 3374 606117 3434 607139
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 22133 3434 606051
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 3371 22132 3437 22133
rect 3371 22068 3372 22132
rect 3436 22068 3437 22132
rect 3371 22067 3437 22068
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 700000 51914 700398
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 700000 87914 700398
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 700000 123914 700398
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 700000 159914 700398
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 700000 195914 700398
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 199331 700364 199397 700365
rect 199331 700300 199332 700364
rect 199396 700300 199397 700364
rect 199331 700299 199397 700300
rect 33868 691954 34868 691986
rect 33868 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 34868 691954
rect 33868 691634 34868 691718
rect 33868 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 34868 691634
rect 33868 691366 34868 691398
rect 53868 691954 54868 691986
rect 53868 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 54868 691954
rect 53868 691634 54868 691718
rect 53868 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 54868 691634
rect 53868 691366 54868 691398
rect 73868 691954 74868 691986
rect 73868 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 74868 691954
rect 73868 691634 74868 691718
rect 73868 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 74868 691634
rect 73868 691366 74868 691398
rect 93868 691954 94868 691986
rect 93868 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 94868 691954
rect 93868 691634 94868 691718
rect 93868 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 94868 691634
rect 93868 691366 94868 691398
rect 113868 691954 114868 691986
rect 113868 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 114868 691954
rect 113868 691634 114868 691718
rect 113868 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 114868 691634
rect 113868 691366 114868 691398
rect 133868 691954 134868 691986
rect 133868 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 134868 691954
rect 133868 691634 134868 691718
rect 133868 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 134868 691634
rect 133868 691366 134868 691398
rect 153868 691954 154868 691986
rect 153868 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 154868 691954
rect 153868 691634 154868 691718
rect 153868 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 154868 691634
rect 153868 691366 154868 691398
rect 173868 691954 174868 691986
rect 173868 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 174868 691954
rect 173868 691634 174868 691718
rect 173868 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 174868 691634
rect 173868 691366 174868 691398
rect 193868 691954 194868 691986
rect 193868 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 194868 691954
rect 193868 691634 194868 691718
rect 193868 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 194868 691634
rect 193868 691366 194868 691398
rect 23868 687454 24868 687486
rect 23868 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 24868 687454
rect 23868 687134 24868 687218
rect 23868 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 24868 687134
rect 23868 686866 24868 686898
rect 43868 687454 44868 687486
rect 43868 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 44868 687454
rect 43868 687134 44868 687218
rect 43868 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 44868 687134
rect 43868 686866 44868 686898
rect 63868 687454 64868 687486
rect 63868 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 64868 687454
rect 63868 687134 64868 687218
rect 63868 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 64868 687134
rect 63868 686866 64868 686898
rect 83868 687454 84868 687486
rect 83868 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 84868 687454
rect 83868 687134 84868 687218
rect 83868 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 84868 687134
rect 83868 686866 84868 686898
rect 103868 687454 104868 687486
rect 103868 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 104868 687454
rect 103868 687134 104868 687218
rect 103868 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 104868 687134
rect 103868 686866 104868 686898
rect 123868 687454 124868 687486
rect 123868 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 124868 687454
rect 123868 687134 124868 687218
rect 123868 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 124868 687134
rect 123868 686866 124868 686898
rect 143868 687454 144868 687486
rect 143868 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 144868 687454
rect 143868 687134 144868 687218
rect 143868 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 144868 687134
rect 143868 686866 144868 686898
rect 163868 687454 164868 687486
rect 163868 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 164868 687454
rect 163868 687134 164868 687218
rect 163868 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 164868 687134
rect 163868 686866 164868 686898
rect 183868 687454 184868 687486
rect 183868 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 184868 687454
rect 183868 687134 184868 687218
rect 183868 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 184868 687134
rect 183868 686866 184868 686898
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 33868 655954 34868 655986
rect 33868 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 34868 655954
rect 33868 655634 34868 655718
rect 33868 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 34868 655634
rect 33868 655366 34868 655398
rect 53868 655954 54868 655986
rect 53868 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 54868 655954
rect 53868 655634 54868 655718
rect 53868 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 54868 655634
rect 53868 655366 54868 655398
rect 73868 655954 74868 655986
rect 73868 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 74868 655954
rect 73868 655634 74868 655718
rect 73868 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 74868 655634
rect 73868 655366 74868 655398
rect 93868 655954 94868 655986
rect 93868 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 94868 655954
rect 93868 655634 94868 655718
rect 93868 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 94868 655634
rect 93868 655366 94868 655398
rect 113868 655954 114868 655986
rect 113868 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 114868 655954
rect 113868 655634 114868 655718
rect 113868 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 114868 655634
rect 113868 655366 114868 655398
rect 133868 655954 134868 655986
rect 133868 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 134868 655954
rect 133868 655634 134868 655718
rect 133868 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 134868 655634
rect 133868 655366 134868 655398
rect 153868 655954 154868 655986
rect 153868 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 154868 655954
rect 153868 655634 154868 655718
rect 153868 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 154868 655634
rect 153868 655366 154868 655398
rect 173868 655954 174868 655986
rect 173868 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 174868 655954
rect 173868 655634 174868 655718
rect 173868 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 174868 655634
rect 173868 655366 174868 655398
rect 193868 655954 194868 655986
rect 193868 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 194868 655954
rect 193868 655634 194868 655718
rect 193868 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 194868 655634
rect 193868 655366 194868 655398
rect 23868 651454 24868 651486
rect 23868 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 24868 651454
rect 23868 651134 24868 651218
rect 23868 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 24868 651134
rect 23868 650866 24868 650898
rect 43868 651454 44868 651486
rect 43868 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 44868 651454
rect 43868 651134 44868 651218
rect 43868 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 44868 651134
rect 43868 650866 44868 650898
rect 63868 651454 64868 651486
rect 63868 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 64868 651454
rect 63868 651134 64868 651218
rect 63868 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 64868 651134
rect 63868 650866 64868 650898
rect 83868 651454 84868 651486
rect 83868 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 84868 651454
rect 83868 651134 84868 651218
rect 83868 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 84868 651134
rect 83868 650866 84868 650898
rect 103868 651454 104868 651486
rect 103868 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 104868 651454
rect 103868 651134 104868 651218
rect 103868 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 104868 651134
rect 103868 650866 104868 650898
rect 123868 651454 124868 651486
rect 123868 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 124868 651454
rect 123868 651134 124868 651218
rect 123868 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 124868 651134
rect 123868 650866 124868 650898
rect 143868 651454 144868 651486
rect 143868 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 144868 651454
rect 143868 651134 144868 651218
rect 143868 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 144868 651134
rect 143868 650866 144868 650898
rect 163868 651454 164868 651486
rect 163868 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 164868 651454
rect 163868 651134 164868 651218
rect 163868 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 164868 651134
rect 163868 650866 164868 650898
rect 183868 651454 184868 651486
rect 183868 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 184868 651454
rect 183868 651134 184868 651218
rect 183868 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 184868 651134
rect 183868 650866 184868 650898
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 33868 619954 34868 619986
rect 33868 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 34868 619954
rect 33868 619634 34868 619718
rect 33868 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 34868 619634
rect 33868 619366 34868 619398
rect 53868 619954 54868 619986
rect 53868 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 54868 619954
rect 53868 619634 54868 619718
rect 53868 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 54868 619634
rect 53868 619366 54868 619398
rect 73868 619954 74868 619986
rect 73868 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 74868 619954
rect 73868 619634 74868 619718
rect 73868 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 74868 619634
rect 73868 619366 74868 619398
rect 93868 619954 94868 619986
rect 93868 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 94868 619954
rect 93868 619634 94868 619718
rect 93868 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 94868 619634
rect 93868 619366 94868 619398
rect 113868 619954 114868 619986
rect 113868 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 114868 619954
rect 113868 619634 114868 619718
rect 113868 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 114868 619634
rect 113868 619366 114868 619398
rect 133868 619954 134868 619986
rect 133868 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 134868 619954
rect 133868 619634 134868 619718
rect 133868 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 134868 619634
rect 133868 619366 134868 619398
rect 153868 619954 154868 619986
rect 153868 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 154868 619954
rect 153868 619634 154868 619718
rect 153868 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 154868 619634
rect 153868 619366 154868 619398
rect 173868 619954 174868 619986
rect 173868 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 174868 619954
rect 173868 619634 174868 619718
rect 173868 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 174868 619634
rect 173868 619366 174868 619398
rect 193868 619954 194868 619986
rect 193868 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 194868 619954
rect 193868 619634 194868 619718
rect 193868 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 194868 619634
rect 193868 619366 194868 619398
rect 23868 615454 24868 615486
rect 23868 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 24868 615454
rect 23868 615134 24868 615218
rect 23868 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 24868 615134
rect 23868 614866 24868 614898
rect 43868 615454 44868 615486
rect 43868 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 44868 615454
rect 43868 615134 44868 615218
rect 43868 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 44868 615134
rect 43868 614866 44868 614898
rect 63868 615454 64868 615486
rect 63868 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 64868 615454
rect 63868 615134 64868 615218
rect 63868 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 64868 615134
rect 63868 614866 64868 614898
rect 83868 615454 84868 615486
rect 83868 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 84868 615454
rect 83868 615134 84868 615218
rect 83868 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 84868 615134
rect 83868 614866 84868 614898
rect 103868 615454 104868 615486
rect 103868 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 104868 615454
rect 103868 615134 104868 615218
rect 103868 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 104868 615134
rect 103868 614866 104868 614898
rect 123868 615454 124868 615486
rect 123868 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 124868 615454
rect 123868 615134 124868 615218
rect 123868 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 124868 615134
rect 123868 614866 124868 614898
rect 143868 615454 144868 615486
rect 143868 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 144868 615454
rect 143868 615134 144868 615218
rect 143868 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 144868 615134
rect 143868 614866 144868 614898
rect 163868 615454 164868 615486
rect 163868 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 164868 615454
rect 163868 615134 164868 615218
rect 163868 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 164868 615134
rect 163868 614866 164868 614898
rect 183868 615454 184868 615486
rect 183868 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 184868 615454
rect 183868 615134 184868 615218
rect 183868 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 184868 615134
rect 183868 614866 184868 614898
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 23243 585852 23309 585853
rect 23243 585788 23244 585852
rect 23308 585788 23309 585852
rect 23243 585787 23309 585788
rect 23059 582996 23125 582997
rect 23059 582932 23060 582996
rect 23124 582932 23125 582996
rect 23059 582931 23125 582932
rect 21955 571980 22021 571981
rect 21955 571916 21956 571980
rect 22020 571916 22021 571980
rect 21955 571915 22021 571916
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 21958 458285 22018 571915
rect 22875 458964 22941 458965
rect 22875 458900 22876 458964
rect 22940 458900 22941 458964
rect 22875 458899 22941 458900
rect 22878 458285 22938 458899
rect 23062 458829 23122 582931
rect 23059 458828 23125 458829
rect 23059 458764 23060 458828
rect 23124 458764 23125 458828
rect 23059 458763 23125 458764
rect 21955 458284 22021 458285
rect 21955 458220 21956 458284
rect 22020 458220 22021 458284
rect 21955 458219 22021 458220
rect 22875 458284 22941 458285
rect 22875 458220 22876 458284
rect 22940 458220 22941 458284
rect 22875 458219 22941 458220
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 21219 357508 21285 357509
rect 21219 357444 21220 357508
rect 21284 357444 21285 357508
rect 21219 357443 21285 357444
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 19563 205732 19629 205733
rect 19563 205668 19564 205732
rect 19628 205668 19629 205732
rect 19563 205667 19629 205668
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 19566 75853 19626 205667
rect 19563 75852 19629 75853
rect 19563 75788 19564 75852
rect 19628 75788 19629 75852
rect 19563 75787 19629 75788
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 57454 20414 76000
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 21222 21997 21282 357443
rect 22878 345030 22938 458219
rect 23246 458149 23306 585787
rect 197307 572116 197373 572117
rect 197307 572052 197308 572116
rect 197372 572052 197373 572116
rect 197307 572051 197373 572052
rect 33868 547954 34868 547986
rect 33868 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 34868 547954
rect 33868 547634 34868 547718
rect 33868 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 34868 547634
rect 33868 547366 34868 547398
rect 53868 547954 54868 547986
rect 53868 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 54868 547954
rect 53868 547634 54868 547718
rect 53868 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 54868 547634
rect 53868 547366 54868 547398
rect 73868 547954 74868 547986
rect 73868 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 74868 547954
rect 73868 547634 74868 547718
rect 73868 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 74868 547634
rect 73868 547366 74868 547398
rect 93868 547954 94868 547986
rect 93868 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 94868 547954
rect 93868 547634 94868 547718
rect 93868 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 94868 547634
rect 93868 547366 94868 547398
rect 113868 547954 114868 547986
rect 113868 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 114868 547954
rect 113868 547634 114868 547718
rect 113868 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 114868 547634
rect 113868 547366 114868 547398
rect 133868 547954 134868 547986
rect 133868 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 134868 547954
rect 133868 547634 134868 547718
rect 133868 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 134868 547634
rect 133868 547366 134868 547398
rect 153868 547954 154868 547986
rect 153868 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 154868 547954
rect 153868 547634 154868 547718
rect 153868 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 154868 547634
rect 153868 547366 154868 547398
rect 173868 547954 174868 547986
rect 173868 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 174868 547954
rect 173868 547634 174868 547718
rect 173868 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 174868 547634
rect 173868 547366 174868 547398
rect 193868 547954 194868 547986
rect 193868 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 194868 547954
rect 193868 547634 194868 547718
rect 193868 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 194868 547634
rect 193868 547366 194868 547398
rect 23868 543454 24868 543486
rect 23868 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 24868 543454
rect 23868 543134 24868 543218
rect 23868 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 24868 543134
rect 23868 542866 24868 542898
rect 43868 543454 44868 543486
rect 43868 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 44868 543454
rect 43868 543134 44868 543218
rect 43868 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 44868 543134
rect 43868 542866 44868 542898
rect 63868 543454 64868 543486
rect 63868 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 64868 543454
rect 63868 543134 64868 543218
rect 63868 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 64868 543134
rect 63868 542866 64868 542898
rect 83868 543454 84868 543486
rect 83868 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 84868 543454
rect 83868 543134 84868 543218
rect 83868 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 84868 543134
rect 83868 542866 84868 542898
rect 103868 543454 104868 543486
rect 103868 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 104868 543454
rect 103868 543134 104868 543218
rect 103868 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 104868 543134
rect 103868 542866 104868 542898
rect 123868 543454 124868 543486
rect 123868 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 124868 543454
rect 123868 543134 124868 543218
rect 123868 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 124868 543134
rect 123868 542866 124868 542898
rect 143868 543454 144868 543486
rect 143868 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 144868 543454
rect 143868 543134 144868 543218
rect 143868 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 144868 543134
rect 143868 542866 144868 542898
rect 163868 543454 164868 543486
rect 163868 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 164868 543454
rect 163868 543134 164868 543218
rect 163868 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 164868 543134
rect 163868 542866 164868 542898
rect 183868 543454 184868 543486
rect 183868 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 184868 543454
rect 183868 543134 184868 543218
rect 183868 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 184868 543134
rect 183868 542866 184868 542898
rect 33868 511954 34868 511986
rect 33868 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 34868 511954
rect 33868 511634 34868 511718
rect 33868 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 34868 511634
rect 33868 511366 34868 511398
rect 53868 511954 54868 511986
rect 53868 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 54868 511954
rect 53868 511634 54868 511718
rect 53868 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 54868 511634
rect 53868 511366 54868 511398
rect 73868 511954 74868 511986
rect 73868 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 74868 511954
rect 73868 511634 74868 511718
rect 73868 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 74868 511634
rect 73868 511366 74868 511398
rect 93868 511954 94868 511986
rect 93868 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 94868 511954
rect 93868 511634 94868 511718
rect 93868 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 94868 511634
rect 93868 511366 94868 511398
rect 113868 511954 114868 511986
rect 113868 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 114868 511954
rect 113868 511634 114868 511718
rect 113868 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 114868 511634
rect 113868 511366 114868 511398
rect 133868 511954 134868 511986
rect 133868 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 134868 511954
rect 133868 511634 134868 511718
rect 133868 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 134868 511634
rect 133868 511366 134868 511398
rect 153868 511954 154868 511986
rect 153868 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 154868 511954
rect 153868 511634 154868 511718
rect 153868 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 154868 511634
rect 153868 511366 154868 511398
rect 173868 511954 174868 511986
rect 173868 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 174868 511954
rect 173868 511634 174868 511718
rect 173868 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 174868 511634
rect 173868 511366 174868 511398
rect 193868 511954 194868 511986
rect 193868 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 194868 511954
rect 193868 511634 194868 511718
rect 193868 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 194868 511634
rect 193868 511366 194868 511398
rect 23868 507454 24868 507486
rect 23868 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 24868 507454
rect 23868 507134 24868 507218
rect 23868 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 24868 507134
rect 23868 506866 24868 506898
rect 43868 507454 44868 507486
rect 43868 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 44868 507454
rect 43868 507134 44868 507218
rect 43868 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 44868 507134
rect 43868 506866 44868 506898
rect 63868 507454 64868 507486
rect 63868 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 64868 507454
rect 63868 507134 64868 507218
rect 63868 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 64868 507134
rect 63868 506866 64868 506898
rect 83868 507454 84868 507486
rect 83868 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 84868 507454
rect 83868 507134 84868 507218
rect 83868 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 84868 507134
rect 83868 506866 84868 506898
rect 103868 507454 104868 507486
rect 103868 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 104868 507454
rect 103868 507134 104868 507218
rect 103868 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 104868 507134
rect 103868 506866 104868 506898
rect 123868 507454 124868 507486
rect 123868 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 124868 507454
rect 123868 507134 124868 507218
rect 123868 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 124868 507134
rect 123868 506866 124868 506898
rect 143868 507454 144868 507486
rect 143868 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 144868 507454
rect 143868 507134 144868 507218
rect 143868 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 144868 507134
rect 143868 506866 144868 506898
rect 163868 507454 164868 507486
rect 163868 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 164868 507454
rect 163868 507134 164868 507218
rect 163868 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 164868 507134
rect 163868 506866 164868 506898
rect 183868 507454 184868 507486
rect 183868 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 184868 507454
rect 183868 507134 184868 507218
rect 183868 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 184868 507134
rect 183868 506866 184868 506898
rect 197310 480270 197370 572051
rect 197310 480210 197922 480270
rect 33868 475954 34868 475986
rect 33868 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 34868 475954
rect 33868 475634 34868 475718
rect 33868 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 34868 475634
rect 33868 475366 34868 475398
rect 53868 475954 54868 475986
rect 53868 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 54868 475954
rect 53868 475634 54868 475718
rect 53868 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 54868 475634
rect 53868 475366 54868 475398
rect 73868 475954 74868 475986
rect 73868 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 74868 475954
rect 73868 475634 74868 475718
rect 73868 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 74868 475634
rect 73868 475366 74868 475398
rect 93868 475954 94868 475986
rect 93868 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 94868 475954
rect 93868 475634 94868 475718
rect 93868 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 94868 475634
rect 93868 475366 94868 475398
rect 113868 475954 114868 475986
rect 113868 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 114868 475954
rect 113868 475634 114868 475718
rect 113868 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 114868 475634
rect 113868 475366 114868 475398
rect 133868 475954 134868 475986
rect 133868 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 134868 475954
rect 133868 475634 134868 475718
rect 133868 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 134868 475634
rect 133868 475366 134868 475398
rect 153868 475954 154868 475986
rect 153868 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 154868 475954
rect 153868 475634 154868 475718
rect 153868 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 154868 475634
rect 153868 475366 154868 475398
rect 173868 475954 174868 475986
rect 173868 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 174868 475954
rect 173868 475634 174868 475718
rect 173868 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 174868 475634
rect 173868 475366 174868 475398
rect 193868 475954 194868 475986
rect 193868 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 194868 475954
rect 193868 475634 194868 475718
rect 193868 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 194868 475634
rect 193868 475366 194868 475398
rect 23868 471454 24868 471486
rect 23868 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 24868 471454
rect 23868 471134 24868 471218
rect 23868 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 24868 471134
rect 23868 470866 24868 470898
rect 43868 471454 44868 471486
rect 43868 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 44868 471454
rect 43868 471134 44868 471218
rect 43868 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 44868 471134
rect 43868 470866 44868 470898
rect 63868 471454 64868 471486
rect 63868 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 64868 471454
rect 63868 471134 64868 471218
rect 63868 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 64868 471134
rect 63868 470866 64868 470898
rect 83868 471454 84868 471486
rect 83868 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 84868 471454
rect 83868 471134 84868 471218
rect 83868 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 84868 471134
rect 83868 470866 84868 470898
rect 103868 471454 104868 471486
rect 103868 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 104868 471454
rect 103868 471134 104868 471218
rect 103868 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 104868 471134
rect 103868 470866 104868 470898
rect 123868 471454 124868 471486
rect 123868 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 124868 471454
rect 123868 471134 124868 471218
rect 123868 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 124868 471134
rect 123868 470866 124868 470898
rect 143868 471454 144868 471486
rect 143868 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 144868 471454
rect 143868 471134 144868 471218
rect 143868 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 144868 471134
rect 143868 470866 144868 470898
rect 163868 471454 164868 471486
rect 163868 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 164868 471454
rect 163868 471134 164868 471218
rect 163868 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 164868 471134
rect 163868 470866 164868 470898
rect 183868 471454 184868 471486
rect 183868 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 184868 471454
rect 183868 471134 184868 471218
rect 183868 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 184868 471134
rect 183868 470866 184868 470898
rect 197862 459373 197922 480210
rect 197859 459372 197925 459373
rect 197859 459308 197860 459372
rect 197924 459308 197925 459372
rect 197859 459307 197925 459308
rect 23243 458148 23309 458149
rect 23243 458084 23244 458148
rect 23308 458084 23309 458148
rect 23243 458083 23309 458084
rect 22878 344970 23122 345030
rect 23062 332485 23122 344970
rect 23059 332484 23125 332485
rect 23059 332420 23060 332484
rect 23124 332420 23125 332484
rect 23059 332419 23125 332420
rect 23062 203013 23122 332419
rect 23246 332349 23306 458083
rect 33868 439954 34868 439986
rect 33868 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 34868 439954
rect 33868 439634 34868 439718
rect 33868 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 34868 439634
rect 33868 439366 34868 439398
rect 53868 439954 54868 439986
rect 53868 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 54868 439954
rect 53868 439634 54868 439718
rect 53868 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 54868 439634
rect 53868 439366 54868 439398
rect 73868 439954 74868 439986
rect 73868 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 74868 439954
rect 73868 439634 74868 439718
rect 73868 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 74868 439634
rect 73868 439366 74868 439398
rect 93868 439954 94868 439986
rect 93868 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 94868 439954
rect 93868 439634 94868 439718
rect 93868 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 94868 439634
rect 93868 439366 94868 439398
rect 113868 439954 114868 439986
rect 113868 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 114868 439954
rect 113868 439634 114868 439718
rect 113868 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 114868 439634
rect 113868 439366 114868 439398
rect 133868 439954 134868 439986
rect 133868 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 134868 439954
rect 133868 439634 134868 439718
rect 133868 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 134868 439634
rect 133868 439366 134868 439398
rect 153868 439954 154868 439986
rect 153868 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 154868 439954
rect 153868 439634 154868 439718
rect 153868 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 154868 439634
rect 153868 439366 154868 439398
rect 173868 439954 174868 439986
rect 173868 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 174868 439954
rect 173868 439634 174868 439718
rect 173868 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 174868 439634
rect 173868 439366 174868 439398
rect 193868 439954 194868 439986
rect 193868 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 194868 439954
rect 193868 439634 194868 439718
rect 193868 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 194868 439634
rect 193868 439366 194868 439398
rect 23868 435454 24868 435486
rect 23868 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 24868 435454
rect 23868 435134 24868 435218
rect 23868 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 24868 435134
rect 23868 434866 24868 434898
rect 43868 435454 44868 435486
rect 43868 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 44868 435454
rect 43868 435134 44868 435218
rect 43868 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 44868 435134
rect 43868 434866 44868 434898
rect 63868 435454 64868 435486
rect 63868 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 64868 435454
rect 63868 435134 64868 435218
rect 63868 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 64868 435134
rect 63868 434866 64868 434898
rect 83868 435454 84868 435486
rect 83868 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 84868 435454
rect 83868 435134 84868 435218
rect 83868 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 84868 435134
rect 83868 434866 84868 434898
rect 103868 435454 104868 435486
rect 103868 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 104868 435454
rect 103868 435134 104868 435218
rect 103868 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 104868 435134
rect 103868 434866 104868 434898
rect 123868 435454 124868 435486
rect 123868 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 124868 435454
rect 123868 435134 124868 435218
rect 123868 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 124868 435134
rect 123868 434866 124868 434898
rect 143868 435454 144868 435486
rect 143868 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 144868 435454
rect 143868 435134 144868 435218
rect 143868 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 144868 435134
rect 143868 434866 144868 434898
rect 163868 435454 164868 435486
rect 163868 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 164868 435454
rect 163868 435134 164868 435218
rect 163868 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 164868 435134
rect 163868 434866 164868 434898
rect 183868 435454 184868 435486
rect 183868 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 184868 435454
rect 183868 435134 184868 435218
rect 183868 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 184868 435134
rect 183868 434866 184868 434898
rect 33868 403954 34868 403986
rect 33868 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 34868 403954
rect 33868 403634 34868 403718
rect 33868 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 34868 403634
rect 33868 403366 34868 403398
rect 53868 403954 54868 403986
rect 53868 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 54868 403954
rect 53868 403634 54868 403718
rect 53868 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 54868 403634
rect 53868 403366 54868 403398
rect 73868 403954 74868 403986
rect 73868 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 74868 403954
rect 73868 403634 74868 403718
rect 73868 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 74868 403634
rect 73868 403366 74868 403398
rect 93868 403954 94868 403986
rect 93868 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 94868 403954
rect 93868 403634 94868 403718
rect 93868 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 94868 403634
rect 93868 403366 94868 403398
rect 113868 403954 114868 403986
rect 113868 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 114868 403954
rect 113868 403634 114868 403718
rect 113868 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 114868 403634
rect 113868 403366 114868 403398
rect 133868 403954 134868 403986
rect 133868 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 134868 403954
rect 133868 403634 134868 403718
rect 133868 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 134868 403634
rect 133868 403366 134868 403398
rect 153868 403954 154868 403986
rect 153868 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 154868 403954
rect 153868 403634 154868 403718
rect 153868 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 154868 403634
rect 153868 403366 154868 403398
rect 173868 403954 174868 403986
rect 173868 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 174868 403954
rect 173868 403634 174868 403718
rect 173868 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 174868 403634
rect 173868 403366 174868 403398
rect 193868 403954 194868 403986
rect 193868 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 194868 403954
rect 193868 403634 194868 403718
rect 193868 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 194868 403634
rect 193868 403366 194868 403398
rect 23868 399454 24868 399486
rect 23868 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 24868 399454
rect 23868 399134 24868 399218
rect 23868 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 24868 399134
rect 23868 398866 24868 398898
rect 43868 399454 44868 399486
rect 43868 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 44868 399454
rect 43868 399134 44868 399218
rect 43868 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 44868 399134
rect 43868 398866 44868 398898
rect 63868 399454 64868 399486
rect 63868 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 64868 399454
rect 63868 399134 64868 399218
rect 63868 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 64868 399134
rect 63868 398866 64868 398898
rect 83868 399454 84868 399486
rect 83868 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 84868 399454
rect 83868 399134 84868 399218
rect 83868 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 84868 399134
rect 83868 398866 84868 398898
rect 103868 399454 104868 399486
rect 103868 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 104868 399454
rect 103868 399134 104868 399218
rect 103868 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 104868 399134
rect 103868 398866 104868 398898
rect 123868 399454 124868 399486
rect 123868 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 124868 399454
rect 123868 399134 124868 399218
rect 123868 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 124868 399134
rect 123868 398866 124868 398898
rect 143868 399454 144868 399486
rect 143868 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 144868 399454
rect 143868 399134 144868 399218
rect 143868 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 144868 399134
rect 143868 398866 144868 398898
rect 163868 399454 164868 399486
rect 163868 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 164868 399454
rect 163868 399134 164868 399218
rect 163868 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 164868 399134
rect 163868 398866 164868 398898
rect 183868 399454 184868 399486
rect 183868 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 184868 399454
rect 183868 399134 184868 399218
rect 183868 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 184868 399134
rect 183868 398866 184868 398898
rect 33868 367954 34868 367986
rect 33868 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 34868 367954
rect 33868 367634 34868 367718
rect 33868 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 34868 367634
rect 33868 367366 34868 367398
rect 53868 367954 54868 367986
rect 53868 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 54868 367954
rect 53868 367634 54868 367718
rect 53868 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 54868 367634
rect 53868 367366 54868 367398
rect 73868 367954 74868 367986
rect 73868 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 74868 367954
rect 73868 367634 74868 367718
rect 73868 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 74868 367634
rect 73868 367366 74868 367398
rect 93868 367954 94868 367986
rect 93868 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 94868 367954
rect 93868 367634 94868 367718
rect 93868 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 94868 367634
rect 93868 367366 94868 367398
rect 113868 367954 114868 367986
rect 113868 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 114868 367954
rect 113868 367634 114868 367718
rect 113868 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 114868 367634
rect 113868 367366 114868 367398
rect 133868 367954 134868 367986
rect 133868 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 134868 367954
rect 133868 367634 134868 367718
rect 133868 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 134868 367634
rect 133868 367366 134868 367398
rect 153868 367954 154868 367986
rect 153868 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 154868 367954
rect 153868 367634 154868 367718
rect 153868 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 154868 367634
rect 153868 367366 154868 367398
rect 173868 367954 174868 367986
rect 173868 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 174868 367954
rect 173868 367634 174868 367718
rect 173868 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 174868 367634
rect 173868 367366 174868 367398
rect 193868 367954 194868 367986
rect 193868 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 194868 367954
rect 193868 367634 194868 367718
rect 193868 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 194868 367634
rect 193868 367366 194868 367398
rect 23868 363454 24868 363486
rect 23868 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 24868 363454
rect 23868 363134 24868 363218
rect 23868 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 24868 363134
rect 23868 362866 24868 362898
rect 43868 363454 44868 363486
rect 43868 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 44868 363454
rect 43868 363134 44868 363218
rect 43868 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 44868 363134
rect 43868 362866 44868 362898
rect 63868 363454 64868 363486
rect 63868 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 64868 363454
rect 63868 363134 64868 363218
rect 63868 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 64868 363134
rect 63868 362866 64868 362898
rect 83868 363454 84868 363486
rect 83868 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 84868 363454
rect 83868 363134 84868 363218
rect 83868 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 84868 363134
rect 83868 362866 84868 362898
rect 103868 363454 104868 363486
rect 103868 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 104868 363454
rect 103868 363134 104868 363218
rect 103868 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 104868 363134
rect 103868 362866 104868 362898
rect 123868 363454 124868 363486
rect 123868 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 124868 363454
rect 123868 363134 124868 363218
rect 123868 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 124868 363134
rect 123868 362866 124868 362898
rect 143868 363454 144868 363486
rect 143868 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 144868 363454
rect 143868 363134 144868 363218
rect 143868 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 144868 363134
rect 143868 362866 144868 362898
rect 163868 363454 164868 363486
rect 163868 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 164868 363454
rect 163868 363134 164868 363218
rect 163868 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 164868 363134
rect 163868 362866 164868 362898
rect 183868 363454 184868 363486
rect 183868 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 184868 363454
rect 183868 363134 184868 363218
rect 183868 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 184868 363134
rect 183868 362866 184868 362898
rect 197862 345030 197922 459307
rect 197862 344970 198658 345030
rect 198598 332757 198658 344970
rect 198595 332756 198661 332757
rect 198595 332692 198596 332756
rect 198660 332692 198661 332756
rect 198595 332691 198661 332692
rect 23243 332348 23309 332349
rect 23243 332284 23244 332348
rect 23308 332284 23309 332348
rect 23243 332283 23309 332284
rect 23059 203012 23125 203013
rect 23059 202948 23060 203012
rect 23124 202948 23125 203012
rect 23059 202947 23125 202948
rect 23246 202741 23306 332283
rect 33868 295954 34868 295986
rect 33868 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 34868 295954
rect 33868 295634 34868 295718
rect 33868 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 34868 295634
rect 33868 295366 34868 295398
rect 53868 295954 54868 295986
rect 53868 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 54868 295954
rect 53868 295634 54868 295718
rect 53868 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 54868 295634
rect 53868 295366 54868 295398
rect 73868 295954 74868 295986
rect 73868 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 74868 295954
rect 73868 295634 74868 295718
rect 73868 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 74868 295634
rect 73868 295366 74868 295398
rect 93868 295954 94868 295986
rect 93868 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 94868 295954
rect 93868 295634 94868 295718
rect 93868 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 94868 295634
rect 93868 295366 94868 295398
rect 113868 295954 114868 295986
rect 113868 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 114868 295954
rect 113868 295634 114868 295718
rect 113868 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 114868 295634
rect 113868 295366 114868 295398
rect 133868 295954 134868 295986
rect 133868 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 134868 295954
rect 133868 295634 134868 295718
rect 133868 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 134868 295634
rect 133868 295366 134868 295398
rect 153868 295954 154868 295986
rect 153868 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 154868 295954
rect 153868 295634 154868 295718
rect 153868 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 154868 295634
rect 153868 295366 154868 295398
rect 173868 295954 174868 295986
rect 173868 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 174868 295954
rect 173868 295634 174868 295718
rect 173868 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 174868 295634
rect 173868 295366 174868 295398
rect 193868 295954 194868 295986
rect 193868 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 194868 295954
rect 193868 295634 194868 295718
rect 193868 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 194868 295634
rect 193868 295366 194868 295398
rect 23868 291454 24868 291486
rect 23868 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 24868 291454
rect 23868 291134 24868 291218
rect 23868 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 24868 291134
rect 23868 290866 24868 290898
rect 43868 291454 44868 291486
rect 43868 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 44868 291454
rect 43868 291134 44868 291218
rect 43868 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 44868 291134
rect 43868 290866 44868 290898
rect 63868 291454 64868 291486
rect 63868 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 64868 291454
rect 63868 291134 64868 291218
rect 63868 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 64868 291134
rect 63868 290866 64868 290898
rect 83868 291454 84868 291486
rect 83868 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 84868 291454
rect 83868 291134 84868 291218
rect 83868 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 84868 291134
rect 83868 290866 84868 290898
rect 103868 291454 104868 291486
rect 103868 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 104868 291454
rect 103868 291134 104868 291218
rect 103868 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 104868 291134
rect 103868 290866 104868 290898
rect 123868 291454 124868 291486
rect 123868 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 124868 291454
rect 123868 291134 124868 291218
rect 123868 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 124868 291134
rect 123868 290866 124868 290898
rect 143868 291454 144868 291486
rect 143868 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 144868 291454
rect 143868 291134 144868 291218
rect 143868 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 144868 291134
rect 143868 290866 144868 290898
rect 163868 291454 164868 291486
rect 163868 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 164868 291454
rect 163868 291134 164868 291218
rect 163868 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 164868 291134
rect 163868 290866 164868 290898
rect 183868 291454 184868 291486
rect 183868 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 184868 291454
rect 183868 291134 184868 291218
rect 183868 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 184868 291134
rect 183868 290866 184868 290898
rect 33868 259954 34868 259986
rect 33868 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 34868 259954
rect 33868 259634 34868 259718
rect 33868 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 34868 259634
rect 33868 259366 34868 259398
rect 53868 259954 54868 259986
rect 53868 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 54868 259954
rect 53868 259634 54868 259718
rect 53868 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 54868 259634
rect 53868 259366 54868 259398
rect 73868 259954 74868 259986
rect 73868 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 74868 259954
rect 73868 259634 74868 259718
rect 73868 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 74868 259634
rect 73868 259366 74868 259398
rect 93868 259954 94868 259986
rect 93868 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 94868 259954
rect 93868 259634 94868 259718
rect 93868 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 94868 259634
rect 93868 259366 94868 259398
rect 113868 259954 114868 259986
rect 113868 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 114868 259954
rect 113868 259634 114868 259718
rect 113868 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 114868 259634
rect 113868 259366 114868 259398
rect 133868 259954 134868 259986
rect 133868 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 134868 259954
rect 133868 259634 134868 259718
rect 133868 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 134868 259634
rect 133868 259366 134868 259398
rect 153868 259954 154868 259986
rect 153868 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 154868 259954
rect 153868 259634 154868 259718
rect 153868 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 154868 259634
rect 153868 259366 154868 259398
rect 173868 259954 174868 259986
rect 173868 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 174868 259954
rect 173868 259634 174868 259718
rect 173868 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 174868 259634
rect 173868 259366 174868 259398
rect 193868 259954 194868 259986
rect 193868 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 194868 259954
rect 193868 259634 194868 259718
rect 193868 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 194868 259634
rect 193868 259366 194868 259398
rect 23868 255454 24868 255486
rect 23868 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 24868 255454
rect 23868 255134 24868 255218
rect 23868 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 24868 255134
rect 23868 254866 24868 254898
rect 43868 255454 44868 255486
rect 43868 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 44868 255454
rect 43868 255134 44868 255218
rect 43868 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 44868 255134
rect 43868 254866 44868 254898
rect 63868 255454 64868 255486
rect 63868 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 64868 255454
rect 63868 255134 64868 255218
rect 63868 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 64868 255134
rect 63868 254866 64868 254898
rect 83868 255454 84868 255486
rect 83868 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 84868 255454
rect 83868 255134 84868 255218
rect 83868 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 84868 255134
rect 83868 254866 84868 254898
rect 103868 255454 104868 255486
rect 103868 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 104868 255454
rect 103868 255134 104868 255218
rect 103868 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 104868 255134
rect 103868 254866 104868 254898
rect 123868 255454 124868 255486
rect 123868 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 124868 255454
rect 123868 255134 124868 255218
rect 123868 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 124868 255134
rect 123868 254866 124868 254898
rect 143868 255454 144868 255486
rect 143868 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 144868 255454
rect 143868 255134 144868 255218
rect 143868 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 144868 255134
rect 143868 254866 144868 254898
rect 163868 255454 164868 255486
rect 163868 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 164868 255454
rect 163868 255134 164868 255218
rect 163868 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 164868 255134
rect 163868 254866 164868 254898
rect 183868 255454 184868 255486
rect 183868 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 184868 255454
rect 183868 255134 184868 255218
rect 183868 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 184868 255134
rect 183868 254866 184868 254898
rect 33868 223954 34868 223986
rect 33868 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 34868 223954
rect 33868 223634 34868 223718
rect 33868 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 34868 223634
rect 33868 223366 34868 223398
rect 53868 223954 54868 223986
rect 53868 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 54868 223954
rect 53868 223634 54868 223718
rect 53868 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 54868 223634
rect 53868 223366 54868 223398
rect 73868 223954 74868 223986
rect 73868 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 74868 223954
rect 73868 223634 74868 223718
rect 73868 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 74868 223634
rect 73868 223366 74868 223398
rect 93868 223954 94868 223986
rect 93868 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 94868 223954
rect 93868 223634 94868 223718
rect 93868 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 94868 223634
rect 93868 223366 94868 223398
rect 113868 223954 114868 223986
rect 113868 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 114868 223954
rect 113868 223634 114868 223718
rect 113868 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 114868 223634
rect 113868 223366 114868 223398
rect 133868 223954 134868 223986
rect 133868 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 134868 223954
rect 133868 223634 134868 223718
rect 133868 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 134868 223634
rect 133868 223366 134868 223398
rect 153868 223954 154868 223986
rect 153868 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 154868 223954
rect 153868 223634 154868 223718
rect 153868 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 154868 223634
rect 153868 223366 154868 223398
rect 173868 223954 174868 223986
rect 173868 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 174868 223954
rect 173868 223634 174868 223718
rect 173868 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 174868 223634
rect 173868 223366 174868 223398
rect 193868 223954 194868 223986
rect 193868 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 194868 223954
rect 193868 223634 194868 223718
rect 193868 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 194868 223634
rect 193868 223366 194868 223398
rect 23868 219454 24868 219486
rect 23868 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 24868 219454
rect 23868 219134 24868 219218
rect 23868 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 24868 219134
rect 23868 218866 24868 218898
rect 43868 219454 44868 219486
rect 43868 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 44868 219454
rect 43868 219134 44868 219218
rect 43868 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 44868 219134
rect 43868 218866 44868 218898
rect 63868 219454 64868 219486
rect 63868 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 64868 219454
rect 63868 219134 64868 219218
rect 63868 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 64868 219134
rect 63868 218866 64868 218898
rect 83868 219454 84868 219486
rect 83868 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 84868 219454
rect 83868 219134 84868 219218
rect 83868 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 84868 219134
rect 83868 218866 84868 218898
rect 103868 219454 104868 219486
rect 103868 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 104868 219454
rect 103868 219134 104868 219218
rect 103868 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 104868 219134
rect 103868 218866 104868 218898
rect 123868 219454 124868 219486
rect 123868 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 124868 219454
rect 123868 219134 124868 219218
rect 123868 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 124868 219134
rect 123868 218866 124868 218898
rect 143868 219454 144868 219486
rect 143868 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 144868 219454
rect 143868 219134 144868 219218
rect 143868 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 144868 219134
rect 143868 218866 144868 218898
rect 163868 219454 164868 219486
rect 163868 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 164868 219454
rect 163868 219134 164868 219218
rect 163868 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 164868 219134
rect 163868 218866 164868 218898
rect 183868 219454 184868 219486
rect 183868 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 184868 219454
rect 183868 219134 184868 219218
rect 183868 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 184868 219134
rect 183868 218866 184868 218898
rect 197859 203012 197925 203013
rect 197859 202948 197860 203012
rect 197924 202948 197925 203012
rect 197859 202947 197925 202948
rect 23243 202740 23309 202741
rect 23243 202676 23244 202740
rect 23308 202676 23309 202740
rect 23243 202675 23309 202676
rect 23246 74493 23306 202675
rect 23868 183454 24868 183486
rect 23868 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 24868 183454
rect 23868 183134 24868 183218
rect 23868 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 24868 183134
rect 23868 182866 24868 182898
rect 43868 183454 44868 183486
rect 43868 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 44868 183454
rect 43868 183134 44868 183218
rect 43868 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 44868 183134
rect 43868 182866 44868 182898
rect 63868 183454 64868 183486
rect 63868 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 64868 183454
rect 63868 183134 64868 183218
rect 63868 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 64868 183134
rect 63868 182866 64868 182898
rect 83868 183454 84868 183486
rect 83868 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 84868 183454
rect 83868 183134 84868 183218
rect 83868 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 84868 183134
rect 83868 182866 84868 182898
rect 103868 183454 104868 183486
rect 103868 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 104868 183454
rect 103868 183134 104868 183218
rect 103868 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 104868 183134
rect 103868 182866 104868 182898
rect 123868 183454 124868 183486
rect 123868 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 124868 183454
rect 123868 183134 124868 183218
rect 123868 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 124868 183134
rect 123868 182866 124868 182898
rect 143868 183454 144868 183486
rect 143868 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 144868 183454
rect 143868 183134 144868 183218
rect 143868 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 144868 183134
rect 143868 182866 144868 182898
rect 163868 183454 164868 183486
rect 163868 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 164868 183454
rect 163868 183134 164868 183218
rect 163868 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 164868 183134
rect 163868 182866 164868 182898
rect 183868 183454 184868 183486
rect 183868 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 184868 183454
rect 183868 183134 184868 183218
rect 183868 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 184868 183134
rect 183868 182866 184868 182898
rect 33868 151954 34868 151986
rect 33868 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 34868 151954
rect 33868 151634 34868 151718
rect 33868 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 34868 151634
rect 33868 151366 34868 151398
rect 53868 151954 54868 151986
rect 53868 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 54868 151954
rect 53868 151634 54868 151718
rect 53868 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 54868 151634
rect 53868 151366 54868 151398
rect 73868 151954 74868 151986
rect 73868 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 74868 151954
rect 73868 151634 74868 151718
rect 73868 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 74868 151634
rect 73868 151366 74868 151398
rect 93868 151954 94868 151986
rect 93868 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 94868 151954
rect 93868 151634 94868 151718
rect 93868 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 94868 151634
rect 93868 151366 94868 151398
rect 113868 151954 114868 151986
rect 113868 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 114868 151954
rect 113868 151634 114868 151718
rect 113868 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 114868 151634
rect 113868 151366 114868 151398
rect 133868 151954 134868 151986
rect 133868 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 134868 151954
rect 133868 151634 134868 151718
rect 133868 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 134868 151634
rect 133868 151366 134868 151398
rect 153868 151954 154868 151986
rect 153868 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 154868 151954
rect 153868 151634 154868 151718
rect 153868 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 154868 151634
rect 153868 151366 154868 151398
rect 173868 151954 174868 151986
rect 173868 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 174868 151954
rect 173868 151634 174868 151718
rect 173868 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 174868 151634
rect 173868 151366 174868 151398
rect 193868 151954 194868 151986
rect 193868 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 194868 151954
rect 193868 151634 194868 151718
rect 193868 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 194868 151634
rect 193868 151366 194868 151398
rect 23868 147454 24868 147486
rect 23868 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 24868 147454
rect 23868 147134 24868 147218
rect 23868 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 24868 147134
rect 23868 146866 24868 146898
rect 43868 147454 44868 147486
rect 43868 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 44868 147454
rect 43868 147134 44868 147218
rect 43868 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 44868 147134
rect 43868 146866 44868 146898
rect 63868 147454 64868 147486
rect 63868 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 64868 147454
rect 63868 147134 64868 147218
rect 63868 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 64868 147134
rect 63868 146866 64868 146898
rect 83868 147454 84868 147486
rect 83868 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 84868 147454
rect 83868 147134 84868 147218
rect 83868 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 84868 147134
rect 83868 146866 84868 146898
rect 103868 147454 104868 147486
rect 103868 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 104868 147454
rect 103868 147134 104868 147218
rect 103868 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 104868 147134
rect 103868 146866 104868 146898
rect 123868 147454 124868 147486
rect 123868 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 124868 147454
rect 123868 147134 124868 147218
rect 123868 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 124868 147134
rect 123868 146866 124868 146898
rect 143868 147454 144868 147486
rect 143868 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 144868 147454
rect 143868 147134 144868 147218
rect 143868 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 144868 147134
rect 143868 146866 144868 146898
rect 163868 147454 164868 147486
rect 163868 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 164868 147454
rect 163868 147134 164868 147218
rect 163868 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 164868 147134
rect 163868 146866 164868 146898
rect 183868 147454 184868 147486
rect 183868 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 184868 147454
rect 183868 147134 184868 147218
rect 183868 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 184868 147134
rect 183868 146866 184868 146898
rect 33868 115954 34868 115986
rect 33868 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 34868 115954
rect 33868 115634 34868 115718
rect 33868 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 34868 115634
rect 33868 115366 34868 115398
rect 53868 115954 54868 115986
rect 53868 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 54868 115954
rect 53868 115634 54868 115718
rect 53868 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 54868 115634
rect 53868 115366 54868 115398
rect 73868 115954 74868 115986
rect 73868 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 74868 115954
rect 73868 115634 74868 115718
rect 73868 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 74868 115634
rect 73868 115366 74868 115398
rect 93868 115954 94868 115986
rect 93868 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 94868 115954
rect 93868 115634 94868 115718
rect 93868 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 94868 115634
rect 93868 115366 94868 115398
rect 113868 115954 114868 115986
rect 113868 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 114868 115954
rect 113868 115634 114868 115718
rect 113868 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 114868 115634
rect 113868 115366 114868 115398
rect 133868 115954 134868 115986
rect 133868 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 134868 115954
rect 133868 115634 134868 115718
rect 133868 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 134868 115634
rect 133868 115366 134868 115398
rect 153868 115954 154868 115986
rect 153868 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 154868 115954
rect 153868 115634 154868 115718
rect 153868 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 154868 115634
rect 153868 115366 154868 115398
rect 173868 115954 174868 115986
rect 173868 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 174868 115954
rect 173868 115634 174868 115718
rect 173868 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 174868 115634
rect 173868 115366 174868 115398
rect 193868 115954 194868 115986
rect 193868 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 194868 115954
rect 193868 115634 194868 115718
rect 193868 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 194868 115634
rect 193868 115366 194868 115398
rect 23868 111454 24868 111486
rect 23868 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 24868 111454
rect 23868 111134 24868 111218
rect 23868 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 24868 111134
rect 23868 110866 24868 110898
rect 43868 111454 44868 111486
rect 43868 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 44868 111454
rect 43868 111134 44868 111218
rect 43868 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 44868 111134
rect 43868 110866 44868 110898
rect 63868 111454 64868 111486
rect 63868 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 64868 111454
rect 63868 111134 64868 111218
rect 63868 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 64868 111134
rect 63868 110866 64868 110898
rect 83868 111454 84868 111486
rect 83868 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 84868 111454
rect 83868 111134 84868 111218
rect 83868 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 84868 111134
rect 83868 110866 84868 110898
rect 103868 111454 104868 111486
rect 103868 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 104868 111454
rect 103868 111134 104868 111218
rect 103868 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 104868 111134
rect 103868 110866 104868 110898
rect 123868 111454 124868 111486
rect 123868 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 124868 111454
rect 123868 111134 124868 111218
rect 123868 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 124868 111134
rect 123868 110866 124868 110898
rect 143868 111454 144868 111486
rect 143868 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 144868 111454
rect 143868 111134 144868 111218
rect 143868 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 144868 111134
rect 143868 110866 144868 110898
rect 163868 111454 164868 111486
rect 163868 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 164868 111454
rect 163868 111134 164868 111218
rect 163868 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 164868 111134
rect 163868 110866 164868 110898
rect 183868 111454 184868 111486
rect 183868 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 184868 111454
rect 183868 111134 184868 111218
rect 183868 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 184868 111134
rect 183868 110866 184868 110898
rect 23243 74492 23309 74493
rect 23243 74428 23244 74492
rect 23308 74428 23309 74492
rect 23243 74427 23309 74428
rect 24294 61954 24914 76000
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 21219 21996 21285 21997
rect 21219 21932 21220 21996
rect 21284 21932 21285 21996
rect 21219 21931 21285 21932
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 66454 29414 76000
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 70954 33914 76000
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 75454 38414 76000
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 43954 42914 76000
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 48454 47414 76000
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 52954 51914 76000
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 76000
rect 98499 75172 98565 75173
rect 98499 75108 98500 75172
rect 98564 75108 98565 75172
rect 98499 75107 98565 75108
rect 98502 58850 98562 75107
rect 105294 70954 105914 76000
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 102731 60756 102797 60757
rect 102731 60692 102732 60756
rect 102796 60692 102797 60756
rect 102731 60691 102797 60692
rect 98502 58790 100034 58850
rect 99974 58717 100034 58790
rect 99971 58716 100037 58717
rect 99971 58652 99972 58716
rect 100036 58652 100037 58716
rect 99971 58651 100037 58652
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 102734 51509 102794 60691
rect 102915 58036 102981 58037
rect 102915 57972 102916 58036
rect 102980 57972 102981 58036
rect 102915 57971 102981 57972
rect 102731 51508 102797 51509
rect 102731 51444 102732 51508
rect 102796 51444 102797 51508
rect 102731 51443 102797 51444
rect 102918 48653 102978 57971
rect 102915 48652 102981 48653
rect 102915 48588 102916 48652
rect 102980 48588 102981 48652
rect 102915 48587 102981 48588
rect 102731 47700 102797 47701
rect 102731 47636 102732 47700
rect 102796 47636 102797 47700
rect 102731 47635 102797 47636
rect 79568 43954 79888 43986
rect 79568 43718 79610 43954
rect 79846 43718 79888 43954
rect 79568 43634 79888 43718
rect 79568 43398 79610 43634
rect 79846 43398 79888 43634
rect 79568 43366 79888 43398
rect 102734 41717 102794 47635
rect 102731 41716 102797 41717
rect 102731 41652 102732 41716
rect 102796 41652 102797 41716
rect 102731 41651 102797 41652
rect 64208 39454 64528 39486
rect 64208 39218 64250 39454
rect 64486 39218 64528 39454
rect 64208 39134 64528 39218
rect 64208 38898 64250 39134
rect 64486 38898 64528 39134
rect 64208 38866 64528 38898
rect 94928 39454 95248 39486
rect 94928 39218 94970 39454
rect 95206 39218 95248 39454
rect 94928 39134 95248 39218
rect 94928 38898 94970 39134
rect 95206 38898 95248 39134
rect 94928 38866 95248 38898
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 73794 3454 74414 22000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 22000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 22000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 22000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 21454 92414 22000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 76000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 76000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 76000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 76000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 76000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 76000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 76000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 76000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 76000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 76000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 76000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 76000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 76000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 76000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 76000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 76000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 76000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 76000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 76000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 76000
rect 197862 63477 197922 202947
rect 198598 201381 198658 332691
rect 198595 201380 198661 201381
rect 198595 201316 198596 201380
rect 198660 201316 198661 201380
rect 198595 201315 198661 201316
rect 197859 63476 197925 63477
rect 197859 63412 197860 63476
rect 197924 63412 197925 63476
rect 197859 63411 197925 63412
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 199334 21861 199394 700299
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 199883 582996 199949 582997
rect 199883 582932 199884 582996
rect 199948 582932 199949 582996
rect 199883 582931 199949 582932
rect 199886 458149 199946 582931
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 199883 458148 199949 458149
rect 199883 458084 199884 458148
rect 199948 458084 199949 458148
rect 199883 458083 199949 458084
rect 199886 316050 199946 458083
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 199886 316029 200130 316050
rect 199886 316028 200133 316029
rect 199886 315990 200068 316028
rect 200067 315964 200068 315990
rect 200132 315964 200133 316028
rect 200067 315963 200133 315964
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 56000 204914 61398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 56000 209414 65898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 56000 213914 70398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 56000 218414 74898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 56000 222914 79398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 56000 227414 83898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 56000 231914 88398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 56000 236414 56898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 56000 240914 61398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 56000 245414 65898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 56000 249914 70398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 56000 254414 74898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 56000 258914 79398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 56000 263414 83898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 56000 267914 88398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 56000 272414 56898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 56000 276914 61398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 56000 281414 65898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 56000 285914 70398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 56000 290414 74898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 700000 303914 700398
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 700000 339914 700398
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 700000 375914 700398
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 700000 411914 700398
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 700000 447914 700398
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 313868 691954 314868 691986
rect 313868 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 314868 691954
rect 313868 691634 314868 691718
rect 313868 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 314868 691634
rect 313868 691366 314868 691398
rect 333868 691954 334868 691986
rect 333868 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 334868 691954
rect 333868 691634 334868 691718
rect 333868 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 334868 691634
rect 333868 691366 334868 691398
rect 353868 691954 354868 691986
rect 353868 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 354868 691954
rect 353868 691634 354868 691718
rect 353868 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 354868 691634
rect 353868 691366 354868 691398
rect 373868 691954 374868 691986
rect 373868 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 374868 691954
rect 373868 691634 374868 691718
rect 373868 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 374868 691634
rect 373868 691366 374868 691398
rect 393868 691954 394868 691986
rect 393868 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 394868 691954
rect 393868 691634 394868 691718
rect 393868 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 394868 691634
rect 393868 691366 394868 691398
rect 413868 691954 414868 691986
rect 413868 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 414868 691954
rect 413868 691634 414868 691718
rect 413868 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 414868 691634
rect 413868 691366 414868 691398
rect 433868 691954 434868 691986
rect 433868 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 434868 691954
rect 433868 691634 434868 691718
rect 433868 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 434868 691634
rect 433868 691366 434868 691398
rect 453868 691954 454868 691986
rect 453868 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 454868 691954
rect 453868 691634 454868 691718
rect 453868 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 454868 691634
rect 453868 691366 454868 691398
rect 473868 691954 474868 691986
rect 473868 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 474868 691954
rect 473868 691634 474868 691718
rect 473868 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 474868 691634
rect 473868 691366 474868 691398
rect 303868 687454 304868 687486
rect 303868 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 304868 687454
rect 303868 687134 304868 687218
rect 303868 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 304868 687134
rect 303868 686866 304868 686898
rect 323868 687454 324868 687486
rect 323868 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 324868 687454
rect 323868 687134 324868 687218
rect 323868 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 324868 687134
rect 323868 686866 324868 686898
rect 343868 687454 344868 687486
rect 343868 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 344868 687454
rect 343868 687134 344868 687218
rect 343868 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 344868 687134
rect 343868 686866 344868 686898
rect 363868 687454 364868 687486
rect 363868 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 364868 687454
rect 363868 687134 364868 687218
rect 363868 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 364868 687134
rect 363868 686866 364868 686898
rect 383868 687454 384868 687486
rect 383868 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 384868 687454
rect 383868 687134 384868 687218
rect 383868 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 384868 687134
rect 383868 686866 384868 686898
rect 403868 687454 404868 687486
rect 403868 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 404868 687454
rect 403868 687134 404868 687218
rect 403868 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 404868 687134
rect 403868 686866 404868 686898
rect 423868 687454 424868 687486
rect 423868 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 424868 687454
rect 423868 687134 424868 687218
rect 423868 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 424868 687134
rect 423868 686866 424868 686898
rect 443868 687454 444868 687486
rect 443868 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 444868 687454
rect 443868 687134 444868 687218
rect 443868 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 444868 687134
rect 443868 686866 444868 686898
rect 463868 687454 464868 687486
rect 463868 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 464868 687454
rect 463868 687134 464868 687218
rect 463868 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 464868 687134
rect 463868 686866 464868 686898
rect 479379 683228 479445 683229
rect 479379 683164 479380 683228
rect 479444 683164 479445 683228
rect 479379 683163 479445 683164
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 313868 655954 314868 655986
rect 313868 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 314868 655954
rect 313868 655634 314868 655718
rect 313868 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 314868 655634
rect 313868 655366 314868 655398
rect 333868 655954 334868 655986
rect 333868 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 334868 655954
rect 333868 655634 334868 655718
rect 333868 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 334868 655634
rect 333868 655366 334868 655398
rect 353868 655954 354868 655986
rect 353868 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 354868 655954
rect 353868 655634 354868 655718
rect 353868 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 354868 655634
rect 353868 655366 354868 655398
rect 373868 655954 374868 655986
rect 373868 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 374868 655954
rect 373868 655634 374868 655718
rect 373868 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 374868 655634
rect 373868 655366 374868 655398
rect 393868 655954 394868 655986
rect 393868 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 394868 655954
rect 393868 655634 394868 655718
rect 393868 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 394868 655634
rect 393868 655366 394868 655398
rect 413868 655954 414868 655986
rect 413868 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 414868 655954
rect 413868 655634 414868 655718
rect 413868 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 414868 655634
rect 413868 655366 414868 655398
rect 433868 655954 434868 655986
rect 433868 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 434868 655954
rect 433868 655634 434868 655718
rect 433868 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 434868 655634
rect 433868 655366 434868 655398
rect 453868 655954 454868 655986
rect 453868 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 454868 655954
rect 453868 655634 454868 655718
rect 453868 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 454868 655634
rect 453868 655366 454868 655398
rect 473868 655954 474868 655986
rect 473868 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 474868 655954
rect 473868 655634 474868 655718
rect 473868 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 474868 655634
rect 473868 655366 474868 655398
rect 303868 651454 304868 651486
rect 303868 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 304868 651454
rect 303868 651134 304868 651218
rect 303868 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 304868 651134
rect 303868 650866 304868 650898
rect 323868 651454 324868 651486
rect 323868 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 324868 651454
rect 323868 651134 324868 651218
rect 323868 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 324868 651134
rect 323868 650866 324868 650898
rect 343868 651454 344868 651486
rect 343868 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 344868 651454
rect 343868 651134 344868 651218
rect 343868 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 344868 651134
rect 343868 650866 344868 650898
rect 363868 651454 364868 651486
rect 363868 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 364868 651454
rect 363868 651134 364868 651218
rect 363868 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 364868 651134
rect 363868 650866 364868 650898
rect 383868 651454 384868 651486
rect 383868 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 384868 651454
rect 383868 651134 384868 651218
rect 383868 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 384868 651134
rect 383868 650866 384868 650898
rect 403868 651454 404868 651486
rect 403868 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 404868 651454
rect 403868 651134 404868 651218
rect 403868 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 404868 651134
rect 403868 650866 404868 650898
rect 423868 651454 424868 651486
rect 423868 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 424868 651454
rect 423868 651134 424868 651218
rect 423868 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 424868 651134
rect 423868 650866 424868 650898
rect 443868 651454 444868 651486
rect 443868 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 444868 651454
rect 443868 651134 444868 651218
rect 443868 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 444868 651134
rect 443868 650866 444868 650898
rect 463868 651454 464868 651486
rect 463868 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 464868 651454
rect 463868 651134 464868 651218
rect 463868 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 464868 651134
rect 463868 650866 464868 650898
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 313868 619954 314868 619986
rect 313868 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 314868 619954
rect 313868 619634 314868 619718
rect 313868 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 314868 619634
rect 313868 619366 314868 619398
rect 333868 619954 334868 619986
rect 333868 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 334868 619954
rect 333868 619634 334868 619718
rect 333868 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 334868 619634
rect 333868 619366 334868 619398
rect 353868 619954 354868 619986
rect 353868 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 354868 619954
rect 353868 619634 354868 619718
rect 353868 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 354868 619634
rect 353868 619366 354868 619398
rect 373868 619954 374868 619986
rect 373868 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 374868 619954
rect 373868 619634 374868 619718
rect 373868 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 374868 619634
rect 373868 619366 374868 619398
rect 393868 619954 394868 619986
rect 393868 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 394868 619954
rect 393868 619634 394868 619718
rect 393868 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 394868 619634
rect 393868 619366 394868 619398
rect 413868 619954 414868 619986
rect 413868 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 414868 619954
rect 413868 619634 414868 619718
rect 413868 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 414868 619634
rect 413868 619366 414868 619398
rect 433868 619954 434868 619986
rect 433868 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 434868 619954
rect 433868 619634 434868 619718
rect 433868 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 434868 619634
rect 433868 619366 434868 619398
rect 453868 619954 454868 619986
rect 453868 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 454868 619954
rect 453868 619634 454868 619718
rect 453868 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 454868 619634
rect 453868 619366 454868 619398
rect 473868 619954 474868 619986
rect 473868 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 474868 619954
rect 473868 619634 474868 619718
rect 473868 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 474868 619634
rect 473868 619366 474868 619398
rect 303868 615454 304868 615486
rect 303868 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 304868 615454
rect 303868 615134 304868 615218
rect 303868 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 304868 615134
rect 303868 614866 304868 614898
rect 323868 615454 324868 615486
rect 323868 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 324868 615454
rect 323868 615134 324868 615218
rect 323868 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 324868 615134
rect 323868 614866 324868 614898
rect 343868 615454 344868 615486
rect 343868 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 344868 615454
rect 343868 615134 344868 615218
rect 343868 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 344868 615134
rect 343868 614866 344868 614898
rect 363868 615454 364868 615486
rect 363868 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 364868 615454
rect 363868 615134 364868 615218
rect 363868 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 364868 615134
rect 363868 614866 364868 614898
rect 383868 615454 384868 615486
rect 383868 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 384868 615454
rect 383868 615134 384868 615218
rect 383868 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 384868 615134
rect 383868 614866 384868 614898
rect 403868 615454 404868 615486
rect 403868 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 404868 615454
rect 403868 615134 404868 615218
rect 403868 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 404868 615134
rect 403868 614866 404868 614898
rect 423868 615454 424868 615486
rect 423868 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 424868 615454
rect 423868 615134 424868 615218
rect 423868 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 424868 615134
rect 423868 614866 424868 614898
rect 443868 615454 444868 615486
rect 443868 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 444868 615454
rect 443868 615134 444868 615218
rect 443868 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 444868 615134
rect 443868 614866 444868 614898
rect 463868 615454 464868 615486
rect 463868 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 464868 615454
rect 463868 615134 464868 615218
rect 463868 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 464868 615134
rect 463868 614866 464868 614898
rect 476619 585716 476685 585717
rect 476619 585652 476620 585716
rect 476684 585652 476685 585716
rect 476619 585651 476685 585652
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 303475 582996 303541 582997
rect 303475 582932 303476 582996
rect 303540 582932 303541 582996
rect 303475 582931 303541 582932
rect 298875 571980 298941 571981
rect 298875 571916 298876 571980
rect 298940 571916 298941 571980
rect 298875 571915 298941 571916
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 56000 294914 79398
rect 298878 57221 298938 571915
rect 299979 462228 300045 462229
rect 299979 462164 299980 462228
rect 300044 462164 300045 462228
rect 299979 462163 300045 462164
rect 299982 315893 300042 462163
rect 303478 458013 303538 582931
rect 313868 547954 314868 547986
rect 313868 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 314868 547954
rect 313868 547634 314868 547718
rect 313868 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 314868 547634
rect 313868 547366 314868 547398
rect 333868 547954 334868 547986
rect 333868 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 334868 547954
rect 333868 547634 334868 547718
rect 333868 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 334868 547634
rect 333868 547366 334868 547398
rect 353868 547954 354868 547986
rect 353868 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 354868 547954
rect 353868 547634 354868 547718
rect 353868 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 354868 547634
rect 353868 547366 354868 547398
rect 373868 547954 374868 547986
rect 373868 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 374868 547954
rect 373868 547634 374868 547718
rect 373868 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 374868 547634
rect 373868 547366 374868 547398
rect 393868 547954 394868 547986
rect 393868 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 394868 547954
rect 393868 547634 394868 547718
rect 393868 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 394868 547634
rect 393868 547366 394868 547398
rect 413868 547954 414868 547986
rect 413868 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 414868 547954
rect 413868 547634 414868 547718
rect 413868 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 414868 547634
rect 413868 547366 414868 547398
rect 433868 547954 434868 547986
rect 433868 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 434868 547954
rect 433868 547634 434868 547718
rect 433868 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 434868 547634
rect 433868 547366 434868 547398
rect 453868 547954 454868 547986
rect 453868 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 454868 547954
rect 453868 547634 454868 547718
rect 453868 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 454868 547634
rect 453868 547366 454868 547398
rect 473868 547954 474868 547986
rect 473868 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 474868 547954
rect 473868 547634 474868 547718
rect 473868 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 474868 547634
rect 473868 547366 474868 547398
rect 303868 543454 304868 543486
rect 303868 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 304868 543454
rect 303868 543134 304868 543218
rect 303868 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 304868 543134
rect 303868 542866 304868 542898
rect 323868 543454 324868 543486
rect 323868 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 324868 543454
rect 323868 543134 324868 543218
rect 323868 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 324868 543134
rect 323868 542866 324868 542898
rect 343868 543454 344868 543486
rect 343868 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 344868 543454
rect 343868 543134 344868 543218
rect 343868 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 344868 543134
rect 343868 542866 344868 542898
rect 363868 543454 364868 543486
rect 363868 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 364868 543454
rect 363868 543134 364868 543218
rect 363868 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 364868 543134
rect 363868 542866 364868 542898
rect 383868 543454 384868 543486
rect 383868 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 384868 543454
rect 383868 543134 384868 543218
rect 383868 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 384868 543134
rect 383868 542866 384868 542898
rect 403868 543454 404868 543486
rect 403868 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 404868 543454
rect 403868 543134 404868 543218
rect 403868 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 404868 543134
rect 403868 542866 404868 542898
rect 423868 543454 424868 543486
rect 423868 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 424868 543454
rect 423868 543134 424868 543218
rect 423868 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 424868 543134
rect 423868 542866 424868 542898
rect 443868 543454 444868 543486
rect 443868 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 444868 543454
rect 443868 543134 444868 543218
rect 443868 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 444868 543134
rect 443868 542866 444868 542898
rect 463868 543454 464868 543486
rect 463868 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 464868 543454
rect 463868 543134 464868 543218
rect 463868 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 464868 543134
rect 463868 542866 464868 542898
rect 476622 533490 476682 585651
rect 477539 533492 477605 533493
rect 477539 533490 477540 533492
rect 476622 533430 477540 533490
rect 477539 533428 477540 533430
rect 477604 533428 477605 533492
rect 477539 533427 477605 533428
rect 313868 511954 314868 511986
rect 313868 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 314868 511954
rect 313868 511634 314868 511718
rect 313868 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 314868 511634
rect 313868 511366 314868 511398
rect 333868 511954 334868 511986
rect 333868 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 334868 511954
rect 333868 511634 334868 511718
rect 333868 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 334868 511634
rect 333868 511366 334868 511398
rect 353868 511954 354868 511986
rect 353868 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 354868 511954
rect 353868 511634 354868 511718
rect 353868 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 354868 511634
rect 353868 511366 354868 511398
rect 373868 511954 374868 511986
rect 373868 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 374868 511954
rect 373868 511634 374868 511718
rect 373868 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 374868 511634
rect 373868 511366 374868 511398
rect 393868 511954 394868 511986
rect 393868 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 394868 511954
rect 393868 511634 394868 511718
rect 393868 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 394868 511634
rect 393868 511366 394868 511398
rect 413868 511954 414868 511986
rect 413868 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 414868 511954
rect 413868 511634 414868 511718
rect 413868 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 414868 511634
rect 413868 511366 414868 511398
rect 433868 511954 434868 511986
rect 433868 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 434868 511954
rect 433868 511634 434868 511718
rect 433868 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 434868 511634
rect 433868 511366 434868 511398
rect 453868 511954 454868 511986
rect 453868 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 454868 511954
rect 453868 511634 454868 511718
rect 453868 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 454868 511634
rect 453868 511366 454868 511398
rect 473868 511954 474868 511986
rect 473868 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 474868 511954
rect 473868 511634 474868 511718
rect 473868 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 474868 511634
rect 473868 511366 474868 511398
rect 303868 507454 304868 507486
rect 303868 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 304868 507454
rect 303868 507134 304868 507218
rect 303868 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 304868 507134
rect 303868 506866 304868 506898
rect 323868 507454 324868 507486
rect 323868 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 324868 507454
rect 323868 507134 324868 507218
rect 323868 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 324868 507134
rect 323868 506866 324868 506898
rect 343868 507454 344868 507486
rect 343868 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 344868 507454
rect 343868 507134 344868 507218
rect 343868 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 344868 507134
rect 343868 506866 344868 506898
rect 363868 507454 364868 507486
rect 363868 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 364868 507454
rect 363868 507134 364868 507218
rect 363868 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 364868 507134
rect 363868 506866 364868 506898
rect 383868 507454 384868 507486
rect 383868 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 384868 507454
rect 383868 507134 384868 507218
rect 383868 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 384868 507134
rect 383868 506866 384868 506898
rect 403868 507454 404868 507486
rect 403868 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 404868 507454
rect 403868 507134 404868 507218
rect 403868 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 404868 507134
rect 403868 506866 404868 506898
rect 423868 507454 424868 507486
rect 423868 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 424868 507454
rect 423868 507134 424868 507218
rect 423868 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 424868 507134
rect 423868 506866 424868 506898
rect 443868 507454 444868 507486
rect 443868 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 444868 507454
rect 443868 507134 444868 507218
rect 443868 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 444868 507134
rect 443868 506866 444868 506898
rect 463868 507454 464868 507486
rect 463868 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 464868 507454
rect 463868 507134 464868 507218
rect 463868 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 464868 507134
rect 463868 506866 464868 506898
rect 313868 475954 314868 475986
rect 313868 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 314868 475954
rect 313868 475634 314868 475718
rect 313868 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 314868 475634
rect 313868 475366 314868 475398
rect 333868 475954 334868 475986
rect 333868 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 334868 475954
rect 333868 475634 334868 475718
rect 333868 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 334868 475634
rect 333868 475366 334868 475398
rect 353868 475954 354868 475986
rect 353868 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 354868 475954
rect 353868 475634 354868 475718
rect 353868 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 354868 475634
rect 353868 475366 354868 475398
rect 373868 475954 374868 475986
rect 373868 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 374868 475954
rect 373868 475634 374868 475718
rect 373868 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 374868 475634
rect 373868 475366 374868 475398
rect 393868 475954 394868 475986
rect 393868 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 394868 475954
rect 393868 475634 394868 475718
rect 393868 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 394868 475634
rect 393868 475366 394868 475398
rect 413868 475954 414868 475986
rect 413868 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 414868 475954
rect 413868 475634 414868 475718
rect 413868 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 414868 475634
rect 413868 475366 414868 475398
rect 433868 475954 434868 475986
rect 433868 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 434868 475954
rect 433868 475634 434868 475718
rect 433868 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 434868 475634
rect 433868 475366 434868 475398
rect 453868 475954 454868 475986
rect 453868 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 454868 475954
rect 453868 475634 454868 475718
rect 453868 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 454868 475634
rect 453868 475366 454868 475398
rect 473868 475954 474868 475986
rect 473868 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 474868 475954
rect 473868 475634 474868 475718
rect 473868 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 474868 475634
rect 473868 475366 474868 475398
rect 303868 471454 304868 471486
rect 303868 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 304868 471454
rect 303868 471134 304868 471218
rect 303868 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 304868 471134
rect 303868 470866 304868 470898
rect 323868 471454 324868 471486
rect 323868 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 324868 471454
rect 323868 471134 324868 471218
rect 323868 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 324868 471134
rect 323868 470866 324868 470898
rect 343868 471454 344868 471486
rect 343868 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 344868 471454
rect 343868 471134 344868 471218
rect 343868 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 344868 471134
rect 343868 470866 344868 470898
rect 363868 471454 364868 471486
rect 363868 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 364868 471454
rect 363868 471134 364868 471218
rect 363868 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 364868 471134
rect 363868 470866 364868 470898
rect 383868 471454 384868 471486
rect 383868 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 384868 471454
rect 383868 471134 384868 471218
rect 383868 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 384868 471134
rect 383868 470866 384868 470898
rect 403868 471454 404868 471486
rect 403868 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 404868 471454
rect 403868 471134 404868 471218
rect 403868 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 404868 471134
rect 403868 470866 404868 470898
rect 423868 471454 424868 471486
rect 423868 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 424868 471454
rect 423868 471134 424868 471218
rect 423868 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 424868 471134
rect 423868 470866 424868 470898
rect 443868 471454 444868 471486
rect 443868 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 444868 471454
rect 443868 471134 444868 471218
rect 443868 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 444868 471134
rect 443868 470866 444868 470898
rect 463868 471454 464868 471486
rect 463868 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 464868 471454
rect 463868 471134 464868 471218
rect 463868 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 464868 471134
rect 463868 470866 464868 470898
rect 479382 460869 479442 683163
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 480299 585852 480365 585853
rect 480299 585788 480300 585852
rect 480364 585788 480365 585852
rect 480299 585787 480365 585788
rect 479379 460868 479445 460869
rect 479379 460804 479380 460868
rect 479444 460804 479445 460868
rect 479379 460803 479445 460804
rect 478827 458284 478893 458285
rect 478827 458220 478828 458284
rect 478892 458220 478893 458284
rect 478827 458219 478893 458220
rect 303475 458012 303541 458013
rect 303475 457948 303476 458012
rect 303540 457948 303541 458012
rect 303475 457947 303541 457948
rect 302739 332484 302805 332485
rect 302739 332420 302740 332484
rect 302804 332420 302805 332484
rect 302739 332419 302805 332420
rect 299979 315892 300045 315893
rect 299979 315828 299980 315892
rect 300044 315828 300045 315892
rect 299979 315827 300045 315828
rect 299982 314805 300042 315827
rect 299979 314804 300045 314805
rect 299979 314740 299980 314804
rect 300044 314740 300045 314804
rect 299979 314739 300045 314740
rect 299979 205732 300045 205733
rect 299979 205668 299980 205732
rect 300044 205668 300045 205732
rect 299979 205667 300045 205668
rect 299982 64837 300042 205667
rect 302742 204237 302802 332419
rect 303478 315621 303538 457947
rect 478091 456924 478157 456925
rect 478091 456860 478092 456924
rect 478156 456860 478157 456924
rect 478091 456859 478157 456860
rect 313868 439954 314868 439986
rect 313868 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 314868 439954
rect 313868 439634 314868 439718
rect 313868 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 314868 439634
rect 313868 439366 314868 439398
rect 333868 439954 334868 439986
rect 333868 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 334868 439954
rect 333868 439634 334868 439718
rect 333868 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 334868 439634
rect 333868 439366 334868 439398
rect 353868 439954 354868 439986
rect 353868 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 354868 439954
rect 353868 439634 354868 439718
rect 353868 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 354868 439634
rect 353868 439366 354868 439398
rect 373868 439954 374868 439986
rect 373868 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 374868 439954
rect 373868 439634 374868 439718
rect 373868 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 374868 439634
rect 373868 439366 374868 439398
rect 393868 439954 394868 439986
rect 393868 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 394868 439954
rect 393868 439634 394868 439718
rect 393868 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 394868 439634
rect 393868 439366 394868 439398
rect 413868 439954 414868 439986
rect 413868 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 414868 439954
rect 413868 439634 414868 439718
rect 413868 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 414868 439634
rect 413868 439366 414868 439398
rect 433868 439954 434868 439986
rect 433868 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 434868 439954
rect 433868 439634 434868 439718
rect 433868 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 434868 439634
rect 433868 439366 434868 439398
rect 453868 439954 454868 439986
rect 453868 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 454868 439954
rect 453868 439634 454868 439718
rect 453868 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 454868 439634
rect 453868 439366 454868 439398
rect 473868 439954 474868 439986
rect 473868 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 474868 439954
rect 473868 439634 474868 439718
rect 473868 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 474868 439634
rect 473868 439366 474868 439398
rect 303868 435454 304868 435486
rect 303868 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 304868 435454
rect 303868 435134 304868 435218
rect 303868 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 304868 435134
rect 303868 434866 304868 434898
rect 323868 435454 324868 435486
rect 323868 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 324868 435454
rect 323868 435134 324868 435218
rect 323868 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 324868 435134
rect 323868 434866 324868 434898
rect 343868 435454 344868 435486
rect 343868 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 344868 435454
rect 343868 435134 344868 435218
rect 343868 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 344868 435134
rect 343868 434866 344868 434898
rect 363868 435454 364868 435486
rect 363868 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 364868 435454
rect 363868 435134 364868 435218
rect 363868 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 364868 435134
rect 363868 434866 364868 434898
rect 383868 435454 384868 435486
rect 383868 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 384868 435454
rect 383868 435134 384868 435218
rect 383868 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 384868 435134
rect 383868 434866 384868 434898
rect 403868 435454 404868 435486
rect 403868 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 404868 435454
rect 403868 435134 404868 435218
rect 403868 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 404868 435134
rect 403868 434866 404868 434898
rect 423868 435454 424868 435486
rect 423868 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 424868 435454
rect 423868 435134 424868 435218
rect 423868 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 424868 435134
rect 423868 434866 424868 434898
rect 443868 435454 444868 435486
rect 443868 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 444868 435454
rect 443868 435134 444868 435218
rect 443868 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 444868 435134
rect 443868 434866 444868 434898
rect 463868 435454 464868 435486
rect 463868 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 464868 435454
rect 463868 435134 464868 435218
rect 463868 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 464868 435134
rect 463868 434866 464868 434898
rect 313868 403954 314868 403986
rect 313868 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 314868 403954
rect 313868 403634 314868 403718
rect 313868 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 314868 403634
rect 313868 403366 314868 403398
rect 333868 403954 334868 403986
rect 333868 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 334868 403954
rect 333868 403634 334868 403718
rect 333868 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 334868 403634
rect 333868 403366 334868 403398
rect 353868 403954 354868 403986
rect 353868 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 354868 403954
rect 353868 403634 354868 403718
rect 353868 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 354868 403634
rect 353868 403366 354868 403398
rect 373868 403954 374868 403986
rect 373868 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 374868 403954
rect 373868 403634 374868 403718
rect 373868 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 374868 403634
rect 373868 403366 374868 403398
rect 393868 403954 394868 403986
rect 393868 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 394868 403954
rect 393868 403634 394868 403718
rect 393868 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 394868 403634
rect 393868 403366 394868 403398
rect 413868 403954 414868 403986
rect 413868 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 414868 403954
rect 413868 403634 414868 403718
rect 413868 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 414868 403634
rect 413868 403366 414868 403398
rect 433868 403954 434868 403986
rect 433868 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 434868 403954
rect 433868 403634 434868 403718
rect 433868 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 434868 403634
rect 433868 403366 434868 403398
rect 453868 403954 454868 403986
rect 453868 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 454868 403954
rect 453868 403634 454868 403718
rect 453868 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 454868 403634
rect 453868 403366 454868 403398
rect 473868 403954 474868 403986
rect 473868 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 474868 403954
rect 473868 403634 474868 403718
rect 473868 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 474868 403634
rect 473868 403366 474868 403398
rect 303868 399454 304868 399486
rect 303868 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 304868 399454
rect 303868 399134 304868 399218
rect 303868 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 304868 399134
rect 303868 398866 304868 398898
rect 323868 399454 324868 399486
rect 323868 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 324868 399454
rect 323868 399134 324868 399218
rect 323868 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 324868 399134
rect 323868 398866 324868 398898
rect 343868 399454 344868 399486
rect 343868 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 344868 399454
rect 343868 399134 344868 399218
rect 343868 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 344868 399134
rect 343868 398866 344868 398898
rect 363868 399454 364868 399486
rect 363868 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 364868 399454
rect 363868 399134 364868 399218
rect 363868 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 364868 399134
rect 363868 398866 364868 398898
rect 383868 399454 384868 399486
rect 383868 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 384868 399454
rect 383868 399134 384868 399218
rect 383868 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 384868 399134
rect 383868 398866 384868 398898
rect 403868 399454 404868 399486
rect 403868 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 404868 399454
rect 403868 399134 404868 399218
rect 403868 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 404868 399134
rect 403868 398866 404868 398898
rect 423868 399454 424868 399486
rect 423868 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 424868 399454
rect 423868 399134 424868 399218
rect 423868 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 424868 399134
rect 423868 398866 424868 398898
rect 443868 399454 444868 399486
rect 443868 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 444868 399454
rect 443868 399134 444868 399218
rect 443868 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 444868 399134
rect 443868 398866 444868 398898
rect 463868 399454 464868 399486
rect 463868 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 464868 399454
rect 463868 399134 464868 399218
rect 463868 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 464868 399134
rect 463868 398866 464868 398898
rect 313868 367954 314868 367986
rect 313868 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 314868 367954
rect 313868 367634 314868 367718
rect 313868 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 314868 367634
rect 313868 367366 314868 367398
rect 333868 367954 334868 367986
rect 333868 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 334868 367954
rect 333868 367634 334868 367718
rect 333868 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 334868 367634
rect 333868 367366 334868 367398
rect 353868 367954 354868 367986
rect 353868 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 354868 367954
rect 353868 367634 354868 367718
rect 353868 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 354868 367634
rect 353868 367366 354868 367398
rect 373868 367954 374868 367986
rect 373868 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 374868 367954
rect 373868 367634 374868 367718
rect 373868 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 374868 367634
rect 373868 367366 374868 367398
rect 393868 367954 394868 367986
rect 393868 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 394868 367954
rect 393868 367634 394868 367718
rect 393868 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 394868 367634
rect 393868 367366 394868 367398
rect 413868 367954 414868 367986
rect 413868 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 414868 367954
rect 413868 367634 414868 367718
rect 413868 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 414868 367634
rect 413868 367366 414868 367398
rect 433868 367954 434868 367986
rect 433868 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 434868 367954
rect 433868 367634 434868 367718
rect 433868 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 434868 367634
rect 433868 367366 434868 367398
rect 453868 367954 454868 367986
rect 453868 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 454868 367954
rect 453868 367634 454868 367718
rect 453868 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 454868 367634
rect 453868 367366 454868 367398
rect 473868 367954 474868 367986
rect 473868 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 474868 367954
rect 473868 367634 474868 367718
rect 473868 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 474868 367634
rect 473868 367366 474868 367398
rect 303868 363454 304868 363486
rect 303868 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 304868 363454
rect 303868 363134 304868 363218
rect 303868 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 304868 363134
rect 303868 362866 304868 362898
rect 323868 363454 324868 363486
rect 323868 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 324868 363454
rect 323868 363134 324868 363218
rect 323868 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 324868 363134
rect 323868 362866 324868 362898
rect 343868 363454 344868 363486
rect 343868 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 344868 363454
rect 343868 363134 344868 363218
rect 343868 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 344868 363134
rect 343868 362866 344868 362898
rect 363868 363454 364868 363486
rect 363868 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 364868 363454
rect 363868 363134 364868 363218
rect 363868 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 364868 363134
rect 363868 362866 364868 362898
rect 383868 363454 384868 363486
rect 383868 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 384868 363454
rect 383868 363134 384868 363218
rect 383868 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 384868 363134
rect 383868 362866 384868 362898
rect 403868 363454 404868 363486
rect 403868 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 404868 363454
rect 403868 363134 404868 363218
rect 403868 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 404868 363134
rect 403868 362866 404868 362898
rect 423868 363454 424868 363486
rect 423868 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 424868 363454
rect 423868 363134 424868 363218
rect 423868 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 424868 363134
rect 423868 362866 424868 362898
rect 443868 363454 444868 363486
rect 443868 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 444868 363454
rect 443868 363134 444868 363218
rect 443868 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 444868 363134
rect 443868 362866 444868 362898
rect 463868 363454 464868 363486
rect 463868 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 464868 363454
rect 463868 363134 464868 363218
rect 463868 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 464868 363134
rect 463868 362866 464868 362898
rect 477539 331260 477605 331261
rect 477539 331196 477540 331260
rect 477604 331196 477605 331260
rect 477539 331195 477605 331196
rect 303475 315620 303541 315621
rect 303475 315556 303476 315620
rect 303540 315556 303541 315620
rect 303475 315555 303541 315556
rect 303478 204373 303538 315555
rect 477355 315348 477421 315349
rect 477355 315284 477356 315348
rect 477420 315284 477421 315348
rect 477355 315283 477421 315284
rect 313868 295954 314868 295986
rect 313868 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 314868 295954
rect 313868 295634 314868 295718
rect 313868 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 314868 295634
rect 313868 295366 314868 295398
rect 333868 295954 334868 295986
rect 333868 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 334868 295954
rect 333868 295634 334868 295718
rect 333868 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 334868 295634
rect 333868 295366 334868 295398
rect 353868 295954 354868 295986
rect 353868 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 354868 295954
rect 353868 295634 354868 295718
rect 353868 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 354868 295634
rect 353868 295366 354868 295398
rect 373868 295954 374868 295986
rect 373868 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 374868 295954
rect 373868 295634 374868 295718
rect 373868 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 374868 295634
rect 373868 295366 374868 295398
rect 393868 295954 394868 295986
rect 393868 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 394868 295954
rect 393868 295634 394868 295718
rect 393868 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 394868 295634
rect 393868 295366 394868 295398
rect 413868 295954 414868 295986
rect 413868 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 414868 295954
rect 413868 295634 414868 295718
rect 413868 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 414868 295634
rect 413868 295366 414868 295398
rect 433868 295954 434868 295986
rect 433868 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 434868 295954
rect 433868 295634 434868 295718
rect 433868 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 434868 295634
rect 433868 295366 434868 295398
rect 453868 295954 454868 295986
rect 453868 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 454868 295954
rect 453868 295634 454868 295718
rect 453868 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 454868 295634
rect 453868 295366 454868 295398
rect 473868 295954 474868 295986
rect 473868 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 474868 295954
rect 473868 295634 474868 295718
rect 473868 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 474868 295634
rect 473868 295366 474868 295398
rect 303868 291454 304868 291486
rect 303868 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 304868 291454
rect 303868 291134 304868 291218
rect 303868 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 304868 291134
rect 303868 290866 304868 290898
rect 323868 291454 324868 291486
rect 323868 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 324868 291454
rect 323868 291134 324868 291218
rect 323868 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 324868 291134
rect 323868 290866 324868 290898
rect 343868 291454 344868 291486
rect 343868 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 344868 291454
rect 343868 291134 344868 291218
rect 343868 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 344868 291134
rect 343868 290866 344868 290898
rect 363868 291454 364868 291486
rect 363868 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 364868 291454
rect 363868 291134 364868 291218
rect 363868 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 364868 291134
rect 363868 290866 364868 290898
rect 383868 291454 384868 291486
rect 383868 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 384868 291454
rect 383868 291134 384868 291218
rect 383868 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 384868 291134
rect 383868 290866 384868 290898
rect 403868 291454 404868 291486
rect 403868 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 404868 291454
rect 403868 291134 404868 291218
rect 403868 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 404868 291134
rect 403868 290866 404868 290898
rect 423868 291454 424868 291486
rect 423868 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 424868 291454
rect 423868 291134 424868 291218
rect 423868 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 424868 291134
rect 423868 290866 424868 290898
rect 443868 291454 444868 291486
rect 443868 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 444868 291454
rect 443868 291134 444868 291218
rect 443868 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 444868 291134
rect 443868 290866 444868 290898
rect 463868 291454 464868 291486
rect 463868 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 464868 291454
rect 463868 291134 464868 291218
rect 463868 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 464868 291134
rect 463868 290866 464868 290898
rect 477358 280170 477418 315283
rect 477542 282930 477602 331195
rect 478094 329765 478154 456859
rect 478091 329764 478157 329765
rect 478091 329700 478092 329764
rect 478156 329700 478157 329764
rect 478091 329699 478157 329700
rect 477542 282870 477970 282930
rect 477358 280110 477786 280170
rect 477539 275364 477605 275365
rect 477539 275300 477540 275364
rect 477604 275300 477605 275364
rect 477539 275299 477605 275300
rect 313868 259954 314868 259986
rect 313868 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 314868 259954
rect 313868 259634 314868 259718
rect 313868 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 314868 259634
rect 313868 259366 314868 259398
rect 333868 259954 334868 259986
rect 333868 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 334868 259954
rect 333868 259634 334868 259718
rect 333868 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 334868 259634
rect 333868 259366 334868 259398
rect 353868 259954 354868 259986
rect 353868 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 354868 259954
rect 353868 259634 354868 259718
rect 353868 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 354868 259634
rect 353868 259366 354868 259398
rect 373868 259954 374868 259986
rect 373868 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 374868 259954
rect 373868 259634 374868 259718
rect 373868 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 374868 259634
rect 373868 259366 374868 259398
rect 393868 259954 394868 259986
rect 393868 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 394868 259954
rect 393868 259634 394868 259718
rect 393868 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 394868 259634
rect 393868 259366 394868 259398
rect 413868 259954 414868 259986
rect 413868 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 414868 259954
rect 413868 259634 414868 259718
rect 413868 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 414868 259634
rect 413868 259366 414868 259398
rect 433868 259954 434868 259986
rect 433868 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 434868 259954
rect 433868 259634 434868 259718
rect 433868 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 434868 259634
rect 433868 259366 434868 259398
rect 453868 259954 454868 259986
rect 453868 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 454868 259954
rect 453868 259634 454868 259718
rect 453868 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 454868 259634
rect 453868 259366 454868 259398
rect 473868 259954 474868 259986
rect 473868 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 474868 259954
rect 473868 259634 474868 259718
rect 473868 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 474868 259634
rect 473868 259366 474868 259398
rect 303868 255454 304868 255486
rect 303868 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 304868 255454
rect 303868 255134 304868 255218
rect 303868 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 304868 255134
rect 303868 254866 304868 254898
rect 323868 255454 324868 255486
rect 323868 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 324868 255454
rect 323868 255134 324868 255218
rect 323868 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 324868 255134
rect 323868 254866 324868 254898
rect 343868 255454 344868 255486
rect 343868 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 344868 255454
rect 343868 255134 344868 255218
rect 343868 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 344868 255134
rect 343868 254866 344868 254898
rect 363868 255454 364868 255486
rect 363868 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 364868 255454
rect 363868 255134 364868 255218
rect 363868 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 364868 255134
rect 363868 254866 364868 254898
rect 383868 255454 384868 255486
rect 383868 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 384868 255454
rect 383868 255134 384868 255218
rect 383868 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 384868 255134
rect 383868 254866 384868 254898
rect 403868 255454 404868 255486
rect 403868 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 404868 255454
rect 403868 255134 404868 255218
rect 403868 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 404868 255134
rect 403868 254866 404868 254898
rect 423868 255454 424868 255486
rect 423868 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 424868 255454
rect 423868 255134 424868 255218
rect 423868 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 424868 255134
rect 423868 254866 424868 254898
rect 443868 255454 444868 255486
rect 443868 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 444868 255454
rect 443868 255134 444868 255218
rect 443868 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 444868 255134
rect 443868 254866 444868 254898
rect 463868 255454 464868 255486
rect 463868 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 464868 255454
rect 463868 255134 464868 255218
rect 463868 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 464868 255134
rect 463868 254866 464868 254898
rect 313868 223954 314868 223986
rect 313868 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 314868 223954
rect 313868 223634 314868 223718
rect 313868 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 314868 223634
rect 313868 223366 314868 223398
rect 333868 223954 334868 223986
rect 333868 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 334868 223954
rect 333868 223634 334868 223718
rect 333868 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 334868 223634
rect 333868 223366 334868 223398
rect 353868 223954 354868 223986
rect 353868 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 354868 223954
rect 353868 223634 354868 223718
rect 353868 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 354868 223634
rect 353868 223366 354868 223398
rect 373868 223954 374868 223986
rect 373868 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 374868 223954
rect 373868 223634 374868 223718
rect 373868 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 374868 223634
rect 373868 223366 374868 223398
rect 393868 223954 394868 223986
rect 393868 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 394868 223954
rect 393868 223634 394868 223718
rect 393868 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 394868 223634
rect 393868 223366 394868 223398
rect 413868 223954 414868 223986
rect 413868 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 414868 223954
rect 413868 223634 414868 223718
rect 413868 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 414868 223634
rect 413868 223366 414868 223398
rect 433868 223954 434868 223986
rect 433868 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 434868 223954
rect 433868 223634 434868 223718
rect 433868 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 434868 223634
rect 433868 223366 434868 223398
rect 453868 223954 454868 223986
rect 453868 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 454868 223954
rect 453868 223634 454868 223718
rect 453868 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 454868 223634
rect 453868 223366 454868 223398
rect 473868 223954 474868 223986
rect 473868 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 474868 223954
rect 473868 223634 474868 223718
rect 473868 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 474868 223634
rect 473868 223366 474868 223398
rect 303868 219454 304868 219486
rect 303868 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 304868 219454
rect 303868 219134 304868 219218
rect 303868 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 304868 219134
rect 303868 218866 304868 218898
rect 323868 219454 324868 219486
rect 323868 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 324868 219454
rect 323868 219134 324868 219218
rect 323868 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 324868 219134
rect 323868 218866 324868 218898
rect 343868 219454 344868 219486
rect 343868 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 344868 219454
rect 343868 219134 344868 219218
rect 343868 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 344868 219134
rect 343868 218866 344868 218898
rect 363868 219454 364868 219486
rect 363868 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 364868 219454
rect 363868 219134 364868 219218
rect 363868 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 364868 219134
rect 363868 218866 364868 218898
rect 383868 219454 384868 219486
rect 383868 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 384868 219454
rect 383868 219134 384868 219218
rect 383868 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 384868 219134
rect 383868 218866 384868 218898
rect 403868 219454 404868 219486
rect 403868 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 404868 219454
rect 403868 219134 404868 219218
rect 403868 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 404868 219134
rect 403868 218866 404868 218898
rect 423868 219454 424868 219486
rect 423868 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 424868 219454
rect 423868 219134 424868 219218
rect 423868 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 424868 219134
rect 423868 218866 424868 218898
rect 443868 219454 444868 219486
rect 443868 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 444868 219454
rect 443868 219134 444868 219218
rect 443868 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 444868 219134
rect 443868 218866 444868 218898
rect 463868 219454 464868 219486
rect 463868 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 464868 219454
rect 463868 219134 464868 219218
rect 463868 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 464868 219134
rect 463868 218866 464868 218898
rect 477355 205732 477421 205733
rect 477355 205668 477356 205732
rect 477420 205668 477421 205732
rect 477355 205667 477421 205668
rect 303475 204372 303541 204373
rect 303475 204370 303476 204372
rect 303294 204310 303476 204370
rect 302739 204236 302805 204237
rect 302739 204172 302740 204236
rect 302804 204172 302805 204236
rect 302739 204171 302805 204172
rect 303294 77893 303354 204310
rect 303475 204308 303476 204310
rect 303540 204308 303541 204372
rect 303475 204307 303541 204308
rect 303475 204236 303541 204237
rect 303475 204172 303476 204236
rect 303540 204172 303541 204236
rect 303475 204171 303541 204172
rect 303291 77892 303357 77893
rect 303291 77828 303292 77892
rect 303356 77828 303357 77892
rect 303291 77827 303357 77828
rect 303478 75173 303538 204171
rect 303868 183454 304868 183486
rect 303868 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 304868 183454
rect 303868 183134 304868 183218
rect 303868 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 304868 183134
rect 303868 182866 304868 182898
rect 323868 183454 324868 183486
rect 323868 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 324868 183454
rect 323868 183134 324868 183218
rect 323868 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 324868 183134
rect 323868 182866 324868 182898
rect 343868 183454 344868 183486
rect 343868 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 344868 183454
rect 343868 183134 344868 183218
rect 343868 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 344868 183134
rect 343868 182866 344868 182898
rect 363868 183454 364868 183486
rect 363868 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 364868 183454
rect 363868 183134 364868 183218
rect 363868 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 364868 183134
rect 363868 182866 364868 182898
rect 383868 183454 384868 183486
rect 383868 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 384868 183454
rect 383868 183134 384868 183218
rect 383868 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 384868 183134
rect 383868 182866 384868 182898
rect 403868 183454 404868 183486
rect 403868 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 404868 183454
rect 403868 183134 404868 183218
rect 403868 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 404868 183134
rect 403868 182866 404868 182898
rect 423868 183454 424868 183486
rect 423868 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 424868 183454
rect 423868 183134 424868 183218
rect 423868 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 424868 183134
rect 423868 182866 424868 182898
rect 443868 183454 444868 183486
rect 443868 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 444868 183454
rect 443868 183134 444868 183218
rect 443868 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 444868 183134
rect 443868 182866 444868 182898
rect 463868 183454 464868 183486
rect 463868 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 464868 183454
rect 463868 183134 464868 183218
rect 463868 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 464868 183134
rect 463868 182866 464868 182898
rect 313868 151954 314868 151986
rect 313868 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 314868 151954
rect 313868 151634 314868 151718
rect 313868 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 314868 151634
rect 313868 151366 314868 151398
rect 333868 151954 334868 151986
rect 333868 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 334868 151954
rect 333868 151634 334868 151718
rect 333868 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 334868 151634
rect 333868 151366 334868 151398
rect 353868 151954 354868 151986
rect 353868 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 354868 151954
rect 353868 151634 354868 151718
rect 353868 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 354868 151634
rect 353868 151366 354868 151398
rect 373868 151954 374868 151986
rect 373868 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 374868 151954
rect 373868 151634 374868 151718
rect 373868 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 374868 151634
rect 373868 151366 374868 151398
rect 393868 151954 394868 151986
rect 393868 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 394868 151954
rect 393868 151634 394868 151718
rect 393868 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 394868 151634
rect 393868 151366 394868 151398
rect 413868 151954 414868 151986
rect 413868 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 414868 151954
rect 413868 151634 414868 151718
rect 413868 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 414868 151634
rect 413868 151366 414868 151398
rect 433868 151954 434868 151986
rect 433868 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 434868 151954
rect 433868 151634 434868 151718
rect 433868 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 434868 151634
rect 433868 151366 434868 151398
rect 453868 151954 454868 151986
rect 453868 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 454868 151954
rect 453868 151634 454868 151718
rect 453868 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 454868 151634
rect 453868 151366 454868 151398
rect 473868 151954 474868 151986
rect 473868 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 474868 151954
rect 473868 151634 474868 151718
rect 473868 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 474868 151634
rect 473868 151366 474868 151398
rect 477358 149970 477418 205667
rect 477542 151330 477602 275299
rect 477726 275090 477786 280110
rect 477910 275365 477970 282870
rect 477907 275364 477973 275365
rect 477907 275300 477908 275364
rect 477972 275300 477973 275364
rect 477907 275299 477973 275300
rect 477726 275030 477970 275090
rect 477910 270510 477970 275030
rect 477726 270450 477970 270510
rect 477726 202877 477786 270450
rect 477723 202876 477789 202877
rect 477723 202812 477724 202876
rect 477788 202812 477789 202876
rect 477723 202811 477789 202812
rect 477726 151830 477786 202811
rect 477726 151770 478154 151830
rect 477542 151270 477970 151330
rect 477539 149972 477605 149973
rect 477539 149970 477540 149972
rect 477358 149910 477540 149970
rect 477539 149908 477540 149910
rect 477604 149908 477605 149972
rect 477539 149907 477605 149908
rect 303868 147454 304868 147486
rect 303868 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 304868 147454
rect 303868 147134 304868 147218
rect 303868 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 304868 147134
rect 303868 146866 304868 146898
rect 323868 147454 324868 147486
rect 323868 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 324868 147454
rect 323868 147134 324868 147218
rect 323868 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 324868 147134
rect 323868 146866 324868 146898
rect 343868 147454 344868 147486
rect 343868 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 344868 147454
rect 343868 147134 344868 147218
rect 343868 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 344868 147134
rect 343868 146866 344868 146898
rect 363868 147454 364868 147486
rect 363868 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 364868 147454
rect 363868 147134 364868 147218
rect 363868 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 364868 147134
rect 363868 146866 364868 146898
rect 383868 147454 384868 147486
rect 383868 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 384868 147454
rect 383868 147134 384868 147218
rect 383868 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 384868 147134
rect 383868 146866 384868 146898
rect 403868 147454 404868 147486
rect 403868 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 404868 147454
rect 403868 147134 404868 147218
rect 403868 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 404868 147134
rect 403868 146866 404868 146898
rect 423868 147454 424868 147486
rect 423868 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 424868 147454
rect 423868 147134 424868 147218
rect 423868 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 424868 147134
rect 423868 146866 424868 146898
rect 443868 147454 444868 147486
rect 443868 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 444868 147454
rect 443868 147134 444868 147218
rect 443868 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 444868 147134
rect 443868 146866 444868 146898
rect 463868 147454 464868 147486
rect 463868 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 464868 147454
rect 477910 147250 477970 151270
rect 463868 147134 464868 147218
rect 463868 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 464868 147134
rect 463868 146866 464868 146898
rect 477542 147190 477970 147250
rect 313868 115954 314868 115986
rect 313868 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 314868 115954
rect 313868 115634 314868 115718
rect 313868 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 314868 115634
rect 313868 115366 314868 115398
rect 333868 115954 334868 115986
rect 333868 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 334868 115954
rect 333868 115634 334868 115718
rect 333868 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 334868 115634
rect 333868 115366 334868 115398
rect 353868 115954 354868 115986
rect 353868 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 354868 115954
rect 353868 115634 354868 115718
rect 353868 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 354868 115634
rect 353868 115366 354868 115398
rect 373868 115954 374868 115986
rect 373868 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 374868 115954
rect 373868 115634 374868 115718
rect 373868 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 374868 115634
rect 373868 115366 374868 115398
rect 393868 115954 394868 115986
rect 393868 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 394868 115954
rect 393868 115634 394868 115718
rect 393868 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 394868 115634
rect 393868 115366 394868 115398
rect 413868 115954 414868 115986
rect 413868 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 414868 115954
rect 413868 115634 414868 115718
rect 413868 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 414868 115634
rect 413868 115366 414868 115398
rect 433868 115954 434868 115986
rect 433868 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 434868 115954
rect 433868 115634 434868 115718
rect 433868 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 434868 115634
rect 433868 115366 434868 115398
rect 453868 115954 454868 115986
rect 453868 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 454868 115954
rect 453868 115634 454868 115718
rect 453868 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 454868 115634
rect 453868 115366 454868 115398
rect 473868 115954 474868 115986
rect 473868 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 474868 115954
rect 473868 115634 474868 115718
rect 473868 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 474868 115634
rect 473868 115366 474868 115398
rect 303868 111454 304868 111486
rect 303868 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 304868 111454
rect 303868 111134 304868 111218
rect 303868 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 304868 111134
rect 303868 110866 304868 110898
rect 323868 111454 324868 111486
rect 323868 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 324868 111454
rect 323868 111134 324868 111218
rect 323868 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 324868 111134
rect 323868 110866 324868 110898
rect 343868 111454 344868 111486
rect 343868 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 344868 111454
rect 343868 111134 344868 111218
rect 343868 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 344868 111134
rect 343868 110866 344868 110898
rect 363868 111454 364868 111486
rect 363868 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 364868 111454
rect 363868 111134 364868 111218
rect 363868 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 364868 111134
rect 363868 110866 364868 110898
rect 383868 111454 384868 111486
rect 383868 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 384868 111454
rect 383868 111134 384868 111218
rect 383868 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 384868 111134
rect 383868 110866 384868 110898
rect 403868 111454 404868 111486
rect 403868 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 404868 111454
rect 403868 111134 404868 111218
rect 403868 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 404868 111134
rect 403868 110866 404868 110898
rect 423868 111454 424868 111486
rect 423868 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 424868 111454
rect 423868 111134 424868 111218
rect 423868 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 424868 111134
rect 423868 110866 424868 110898
rect 443868 111454 444868 111486
rect 443868 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 444868 111454
rect 443868 111134 444868 111218
rect 443868 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 444868 111134
rect 443868 110866 444868 110898
rect 463868 111454 464868 111486
rect 463868 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 464868 111454
rect 463868 111134 464868 111218
rect 463868 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 464868 111134
rect 463868 110866 464868 110898
rect 477542 84210 477602 147190
rect 478094 142170 478154 151770
rect 477726 142110 478154 142170
rect 477726 93870 477786 142110
rect 477726 93810 477970 93870
rect 477542 84150 477786 84210
rect 477539 81972 477605 81973
rect 477539 81970 477540 81972
rect 476622 81910 477540 81970
rect 303475 75172 303541 75173
rect 303475 75108 303476 75172
rect 303540 75108 303541 75172
rect 303475 75107 303541 75108
rect 299979 64836 300045 64837
rect 299979 64772 299980 64836
rect 300044 64772 300045 64836
rect 299979 64771 300045 64772
rect 298875 57220 298941 57221
rect 298875 57156 298876 57220
rect 298940 57156 298941 57220
rect 298875 57155 298941 57156
rect 213868 43954 214868 43986
rect 213868 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 214868 43954
rect 213868 43634 214868 43718
rect 213868 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 214868 43634
rect 213868 43366 214868 43398
rect 233868 43954 234868 43986
rect 233868 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 234868 43954
rect 233868 43634 234868 43718
rect 233868 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 234868 43634
rect 233868 43366 234868 43398
rect 253868 43954 254868 43986
rect 253868 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 254868 43954
rect 253868 43634 254868 43718
rect 253868 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 254868 43634
rect 253868 43366 254868 43398
rect 273868 43954 274868 43986
rect 273868 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 274868 43954
rect 273868 43634 274868 43718
rect 273868 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 274868 43634
rect 273868 43366 274868 43398
rect 293868 43954 294868 43986
rect 293868 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 294868 43954
rect 293868 43634 294868 43718
rect 293868 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 294868 43634
rect 293868 43366 294868 43398
rect 313868 43954 314868 43986
rect 313868 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 314868 43954
rect 313868 43634 314868 43718
rect 313868 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 314868 43634
rect 313868 43366 314868 43398
rect 333868 43954 334868 43986
rect 333868 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 334868 43954
rect 333868 43634 334868 43718
rect 333868 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 334868 43634
rect 333868 43366 334868 43398
rect 353868 43954 354868 43986
rect 353868 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 354868 43954
rect 353868 43634 354868 43718
rect 353868 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 354868 43634
rect 353868 43366 354868 43398
rect 373868 43954 374868 43986
rect 373868 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 374868 43954
rect 373868 43634 374868 43718
rect 373868 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 374868 43634
rect 373868 43366 374868 43398
rect 393868 43954 394868 43986
rect 393868 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 394868 43954
rect 393868 43634 394868 43718
rect 393868 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 394868 43634
rect 393868 43366 394868 43398
rect 402294 43954 402914 76000
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 203868 39454 204868 39486
rect 203868 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 204868 39454
rect 203868 39134 204868 39218
rect 203868 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 204868 39134
rect 203868 38866 204868 38898
rect 223868 39454 224868 39486
rect 223868 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 224868 39454
rect 223868 39134 224868 39218
rect 223868 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 224868 39134
rect 223868 38866 224868 38898
rect 243868 39454 244868 39486
rect 243868 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 244868 39454
rect 243868 39134 244868 39218
rect 243868 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 244868 39134
rect 243868 38866 244868 38898
rect 263868 39454 264868 39486
rect 263868 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 264868 39454
rect 263868 39134 264868 39218
rect 263868 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 264868 39134
rect 263868 38866 264868 38898
rect 283868 39454 284868 39486
rect 283868 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 284868 39454
rect 283868 39134 284868 39218
rect 283868 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 284868 39134
rect 283868 38866 284868 38898
rect 303868 39454 304868 39486
rect 303868 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 304868 39454
rect 303868 39134 304868 39218
rect 303868 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 304868 39134
rect 303868 38866 304868 38898
rect 323868 39454 324868 39486
rect 323868 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 324868 39454
rect 323868 39134 324868 39218
rect 323868 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 324868 39134
rect 323868 38866 324868 38898
rect 343868 39454 344868 39486
rect 343868 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 344868 39454
rect 343868 39134 344868 39218
rect 343868 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 344868 39134
rect 343868 38866 344868 38898
rect 363868 39454 364868 39486
rect 363868 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 364868 39454
rect 363868 39134 364868 39218
rect 363868 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 364868 39134
rect 363868 38866 364868 38898
rect 383868 39454 384868 39486
rect 383868 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 384868 39454
rect 383868 39134 384868 39218
rect 383868 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 384868 39134
rect 383868 38866 384868 38898
rect 199331 21860 199397 21861
rect 199331 21796 199332 21860
rect 199396 21796 199397 21860
rect 199331 21795 199397 21796
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 22000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 217794 3454 218414 22000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 22000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 22000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 22000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 22000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 253794 3454 254414 22000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 22000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 22000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 22000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 22000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 289794 3454 290414 22000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 22000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 22000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 22000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 22000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 325794 3454 326414 22000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 22000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 22000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 22000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 22000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 361794 3454 362414 22000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 22000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 22000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 22000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 22000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 397794 3454 398414 22000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 48454 407414 76000
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 52954 411914 76000
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 57454 416414 76000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 61954 420914 76000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 76000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 70954 429914 76000
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 75454 434414 76000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 43954 438914 76000
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 48454 443414 76000
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 52954 447914 76000
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 57454 452414 76000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 76000
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 66454 461414 76000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 70954 465914 76000
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 75454 470414 76000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 43954 474914 76000
rect 476622 73133 476682 81910
rect 477539 81908 477540 81910
rect 477604 81908 477605 81972
rect 477539 81907 477605 81908
rect 477726 78165 477786 84150
rect 477910 81973 477970 93810
rect 477907 81972 477973 81973
rect 477907 81908 477908 81972
rect 477972 81908 477973 81972
rect 477907 81907 477973 81908
rect 477723 78164 477789 78165
rect 477723 78100 477724 78164
rect 477788 78100 477789 78164
rect 477723 78099 477789 78100
rect 478830 78029 478890 458219
rect 478827 78028 478893 78029
rect 478827 77964 478828 78028
rect 478892 77964 478893 78028
rect 478827 77963 478893 77964
rect 480302 77349 480362 585787
rect 481587 585172 481653 585173
rect 481587 585108 481588 585172
rect 481652 585108 481653 585172
rect 481587 585107 481653 585108
rect 481590 77893 481650 585107
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 481587 77892 481653 77893
rect 481587 77828 481588 77892
rect 481652 77828 481653 77892
rect 481587 77827 481653 77828
rect 480299 77348 480365 77349
rect 480299 77284 480300 77348
rect 480364 77284 480365 77348
rect 480299 77283 480365 77284
rect 476619 73132 476685 73133
rect 476619 73068 476620 73132
rect 476684 73068 476685 73132
rect 476619 73067 476685 73068
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 48454 479414 76000
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 580763 418300 580829 418301
rect 580763 418236 580764 418300
rect 580828 418236 580829 418300
rect 580763 418235 580829 418236
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 580766 78437 580826 418235
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 580763 78436 580829 78437
rect 580763 78372 580764 78436
rect 580828 78372 580829 78436
rect 580763 78371 580829 78372
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 33930 691718 34166 691954
rect 34250 691718 34486 691954
rect 34570 691718 34806 691954
rect 33930 691398 34166 691634
rect 34250 691398 34486 691634
rect 34570 691398 34806 691634
rect 53930 691718 54166 691954
rect 54250 691718 54486 691954
rect 54570 691718 54806 691954
rect 53930 691398 54166 691634
rect 54250 691398 54486 691634
rect 54570 691398 54806 691634
rect 73930 691718 74166 691954
rect 74250 691718 74486 691954
rect 74570 691718 74806 691954
rect 73930 691398 74166 691634
rect 74250 691398 74486 691634
rect 74570 691398 74806 691634
rect 93930 691718 94166 691954
rect 94250 691718 94486 691954
rect 94570 691718 94806 691954
rect 93930 691398 94166 691634
rect 94250 691398 94486 691634
rect 94570 691398 94806 691634
rect 113930 691718 114166 691954
rect 114250 691718 114486 691954
rect 114570 691718 114806 691954
rect 113930 691398 114166 691634
rect 114250 691398 114486 691634
rect 114570 691398 114806 691634
rect 133930 691718 134166 691954
rect 134250 691718 134486 691954
rect 134570 691718 134806 691954
rect 133930 691398 134166 691634
rect 134250 691398 134486 691634
rect 134570 691398 134806 691634
rect 153930 691718 154166 691954
rect 154250 691718 154486 691954
rect 154570 691718 154806 691954
rect 153930 691398 154166 691634
rect 154250 691398 154486 691634
rect 154570 691398 154806 691634
rect 173930 691718 174166 691954
rect 174250 691718 174486 691954
rect 174570 691718 174806 691954
rect 173930 691398 174166 691634
rect 174250 691398 174486 691634
rect 174570 691398 174806 691634
rect 193930 691718 194166 691954
rect 194250 691718 194486 691954
rect 194570 691718 194806 691954
rect 193930 691398 194166 691634
rect 194250 691398 194486 691634
rect 194570 691398 194806 691634
rect 23930 687218 24166 687454
rect 24250 687218 24486 687454
rect 24570 687218 24806 687454
rect 23930 686898 24166 687134
rect 24250 686898 24486 687134
rect 24570 686898 24806 687134
rect 43930 687218 44166 687454
rect 44250 687218 44486 687454
rect 44570 687218 44806 687454
rect 43930 686898 44166 687134
rect 44250 686898 44486 687134
rect 44570 686898 44806 687134
rect 63930 687218 64166 687454
rect 64250 687218 64486 687454
rect 64570 687218 64806 687454
rect 63930 686898 64166 687134
rect 64250 686898 64486 687134
rect 64570 686898 64806 687134
rect 83930 687218 84166 687454
rect 84250 687218 84486 687454
rect 84570 687218 84806 687454
rect 83930 686898 84166 687134
rect 84250 686898 84486 687134
rect 84570 686898 84806 687134
rect 103930 687218 104166 687454
rect 104250 687218 104486 687454
rect 104570 687218 104806 687454
rect 103930 686898 104166 687134
rect 104250 686898 104486 687134
rect 104570 686898 104806 687134
rect 123930 687218 124166 687454
rect 124250 687218 124486 687454
rect 124570 687218 124806 687454
rect 123930 686898 124166 687134
rect 124250 686898 124486 687134
rect 124570 686898 124806 687134
rect 143930 687218 144166 687454
rect 144250 687218 144486 687454
rect 144570 687218 144806 687454
rect 143930 686898 144166 687134
rect 144250 686898 144486 687134
rect 144570 686898 144806 687134
rect 163930 687218 164166 687454
rect 164250 687218 164486 687454
rect 164570 687218 164806 687454
rect 163930 686898 164166 687134
rect 164250 686898 164486 687134
rect 164570 686898 164806 687134
rect 183930 687218 184166 687454
rect 184250 687218 184486 687454
rect 184570 687218 184806 687454
rect 183930 686898 184166 687134
rect 184250 686898 184486 687134
rect 184570 686898 184806 687134
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 33930 655718 34166 655954
rect 34250 655718 34486 655954
rect 34570 655718 34806 655954
rect 33930 655398 34166 655634
rect 34250 655398 34486 655634
rect 34570 655398 34806 655634
rect 53930 655718 54166 655954
rect 54250 655718 54486 655954
rect 54570 655718 54806 655954
rect 53930 655398 54166 655634
rect 54250 655398 54486 655634
rect 54570 655398 54806 655634
rect 73930 655718 74166 655954
rect 74250 655718 74486 655954
rect 74570 655718 74806 655954
rect 73930 655398 74166 655634
rect 74250 655398 74486 655634
rect 74570 655398 74806 655634
rect 93930 655718 94166 655954
rect 94250 655718 94486 655954
rect 94570 655718 94806 655954
rect 93930 655398 94166 655634
rect 94250 655398 94486 655634
rect 94570 655398 94806 655634
rect 113930 655718 114166 655954
rect 114250 655718 114486 655954
rect 114570 655718 114806 655954
rect 113930 655398 114166 655634
rect 114250 655398 114486 655634
rect 114570 655398 114806 655634
rect 133930 655718 134166 655954
rect 134250 655718 134486 655954
rect 134570 655718 134806 655954
rect 133930 655398 134166 655634
rect 134250 655398 134486 655634
rect 134570 655398 134806 655634
rect 153930 655718 154166 655954
rect 154250 655718 154486 655954
rect 154570 655718 154806 655954
rect 153930 655398 154166 655634
rect 154250 655398 154486 655634
rect 154570 655398 154806 655634
rect 173930 655718 174166 655954
rect 174250 655718 174486 655954
rect 174570 655718 174806 655954
rect 173930 655398 174166 655634
rect 174250 655398 174486 655634
rect 174570 655398 174806 655634
rect 193930 655718 194166 655954
rect 194250 655718 194486 655954
rect 194570 655718 194806 655954
rect 193930 655398 194166 655634
rect 194250 655398 194486 655634
rect 194570 655398 194806 655634
rect 23930 651218 24166 651454
rect 24250 651218 24486 651454
rect 24570 651218 24806 651454
rect 23930 650898 24166 651134
rect 24250 650898 24486 651134
rect 24570 650898 24806 651134
rect 43930 651218 44166 651454
rect 44250 651218 44486 651454
rect 44570 651218 44806 651454
rect 43930 650898 44166 651134
rect 44250 650898 44486 651134
rect 44570 650898 44806 651134
rect 63930 651218 64166 651454
rect 64250 651218 64486 651454
rect 64570 651218 64806 651454
rect 63930 650898 64166 651134
rect 64250 650898 64486 651134
rect 64570 650898 64806 651134
rect 83930 651218 84166 651454
rect 84250 651218 84486 651454
rect 84570 651218 84806 651454
rect 83930 650898 84166 651134
rect 84250 650898 84486 651134
rect 84570 650898 84806 651134
rect 103930 651218 104166 651454
rect 104250 651218 104486 651454
rect 104570 651218 104806 651454
rect 103930 650898 104166 651134
rect 104250 650898 104486 651134
rect 104570 650898 104806 651134
rect 123930 651218 124166 651454
rect 124250 651218 124486 651454
rect 124570 651218 124806 651454
rect 123930 650898 124166 651134
rect 124250 650898 124486 651134
rect 124570 650898 124806 651134
rect 143930 651218 144166 651454
rect 144250 651218 144486 651454
rect 144570 651218 144806 651454
rect 143930 650898 144166 651134
rect 144250 650898 144486 651134
rect 144570 650898 144806 651134
rect 163930 651218 164166 651454
rect 164250 651218 164486 651454
rect 164570 651218 164806 651454
rect 163930 650898 164166 651134
rect 164250 650898 164486 651134
rect 164570 650898 164806 651134
rect 183930 651218 184166 651454
rect 184250 651218 184486 651454
rect 184570 651218 184806 651454
rect 183930 650898 184166 651134
rect 184250 650898 184486 651134
rect 184570 650898 184806 651134
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 33930 619718 34166 619954
rect 34250 619718 34486 619954
rect 34570 619718 34806 619954
rect 33930 619398 34166 619634
rect 34250 619398 34486 619634
rect 34570 619398 34806 619634
rect 53930 619718 54166 619954
rect 54250 619718 54486 619954
rect 54570 619718 54806 619954
rect 53930 619398 54166 619634
rect 54250 619398 54486 619634
rect 54570 619398 54806 619634
rect 73930 619718 74166 619954
rect 74250 619718 74486 619954
rect 74570 619718 74806 619954
rect 73930 619398 74166 619634
rect 74250 619398 74486 619634
rect 74570 619398 74806 619634
rect 93930 619718 94166 619954
rect 94250 619718 94486 619954
rect 94570 619718 94806 619954
rect 93930 619398 94166 619634
rect 94250 619398 94486 619634
rect 94570 619398 94806 619634
rect 113930 619718 114166 619954
rect 114250 619718 114486 619954
rect 114570 619718 114806 619954
rect 113930 619398 114166 619634
rect 114250 619398 114486 619634
rect 114570 619398 114806 619634
rect 133930 619718 134166 619954
rect 134250 619718 134486 619954
rect 134570 619718 134806 619954
rect 133930 619398 134166 619634
rect 134250 619398 134486 619634
rect 134570 619398 134806 619634
rect 153930 619718 154166 619954
rect 154250 619718 154486 619954
rect 154570 619718 154806 619954
rect 153930 619398 154166 619634
rect 154250 619398 154486 619634
rect 154570 619398 154806 619634
rect 173930 619718 174166 619954
rect 174250 619718 174486 619954
rect 174570 619718 174806 619954
rect 173930 619398 174166 619634
rect 174250 619398 174486 619634
rect 174570 619398 174806 619634
rect 193930 619718 194166 619954
rect 194250 619718 194486 619954
rect 194570 619718 194806 619954
rect 193930 619398 194166 619634
rect 194250 619398 194486 619634
rect 194570 619398 194806 619634
rect 23930 615218 24166 615454
rect 24250 615218 24486 615454
rect 24570 615218 24806 615454
rect 23930 614898 24166 615134
rect 24250 614898 24486 615134
rect 24570 614898 24806 615134
rect 43930 615218 44166 615454
rect 44250 615218 44486 615454
rect 44570 615218 44806 615454
rect 43930 614898 44166 615134
rect 44250 614898 44486 615134
rect 44570 614898 44806 615134
rect 63930 615218 64166 615454
rect 64250 615218 64486 615454
rect 64570 615218 64806 615454
rect 63930 614898 64166 615134
rect 64250 614898 64486 615134
rect 64570 614898 64806 615134
rect 83930 615218 84166 615454
rect 84250 615218 84486 615454
rect 84570 615218 84806 615454
rect 83930 614898 84166 615134
rect 84250 614898 84486 615134
rect 84570 614898 84806 615134
rect 103930 615218 104166 615454
rect 104250 615218 104486 615454
rect 104570 615218 104806 615454
rect 103930 614898 104166 615134
rect 104250 614898 104486 615134
rect 104570 614898 104806 615134
rect 123930 615218 124166 615454
rect 124250 615218 124486 615454
rect 124570 615218 124806 615454
rect 123930 614898 124166 615134
rect 124250 614898 124486 615134
rect 124570 614898 124806 615134
rect 143930 615218 144166 615454
rect 144250 615218 144486 615454
rect 144570 615218 144806 615454
rect 143930 614898 144166 615134
rect 144250 614898 144486 615134
rect 144570 614898 144806 615134
rect 163930 615218 164166 615454
rect 164250 615218 164486 615454
rect 164570 615218 164806 615454
rect 163930 614898 164166 615134
rect 164250 614898 164486 615134
rect 164570 614898 164806 615134
rect 183930 615218 184166 615454
rect 184250 615218 184486 615454
rect 184570 615218 184806 615454
rect 183930 614898 184166 615134
rect 184250 614898 184486 615134
rect 184570 614898 184806 615134
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 33930 547718 34166 547954
rect 34250 547718 34486 547954
rect 34570 547718 34806 547954
rect 33930 547398 34166 547634
rect 34250 547398 34486 547634
rect 34570 547398 34806 547634
rect 53930 547718 54166 547954
rect 54250 547718 54486 547954
rect 54570 547718 54806 547954
rect 53930 547398 54166 547634
rect 54250 547398 54486 547634
rect 54570 547398 54806 547634
rect 73930 547718 74166 547954
rect 74250 547718 74486 547954
rect 74570 547718 74806 547954
rect 73930 547398 74166 547634
rect 74250 547398 74486 547634
rect 74570 547398 74806 547634
rect 93930 547718 94166 547954
rect 94250 547718 94486 547954
rect 94570 547718 94806 547954
rect 93930 547398 94166 547634
rect 94250 547398 94486 547634
rect 94570 547398 94806 547634
rect 113930 547718 114166 547954
rect 114250 547718 114486 547954
rect 114570 547718 114806 547954
rect 113930 547398 114166 547634
rect 114250 547398 114486 547634
rect 114570 547398 114806 547634
rect 133930 547718 134166 547954
rect 134250 547718 134486 547954
rect 134570 547718 134806 547954
rect 133930 547398 134166 547634
rect 134250 547398 134486 547634
rect 134570 547398 134806 547634
rect 153930 547718 154166 547954
rect 154250 547718 154486 547954
rect 154570 547718 154806 547954
rect 153930 547398 154166 547634
rect 154250 547398 154486 547634
rect 154570 547398 154806 547634
rect 173930 547718 174166 547954
rect 174250 547718 174486 547954
rect 174570 547718 174806 547954
rect 173930 547398 174166 547634
rect 174250 547398 174486 547634
rect 174570 547398 174806 547634
rect 193930 547718 194166 547954
rect 194250 547718 194486 547954
rect 194570 547718 194806 547954
rect 193930 547398 194166 547634
rect 194250 547398 194486 547634
rect 194570 547398 194806 547634
rect 23930 543218 24166 543454
rect 24250 543218 24486 543454
rect 24570 543218 24806 543454
rect 23930 542898 24166 543134
rect 24250 542898 24486 543134
rect 24570 542898 24806 543134
rect 43930 543218 44166 543454
rect 44250 543218 44486 543454
rect 44570 543218 44806 543454
rect 43930 542898 44166 543134
rect 44250 542898 44486 543134
rect 44570 542898 44806 543134
rect 63930 543218 64166 543454
rect 64250 543218 64486 543454
rect 64570 543218 64806 543454
rect 63930 542898 64166 543134
rect 64250 542898 64486 543134
rect 64570 542898 64806 543134
rect 83930 543218 84166 543454
rect 84250 543218 84486 543454
rect 84570 543218 84806 543454
rect 83930 542898 84166 543134
rect 84250 542898 84486 543134
rect 84570 542898 84806 543134
rect 103930 543218 104166 543454
rect 104250 543218 104486 543454
rect 104570 543218 104806 543454
rect 103930 542898 104166 543134
rect 104250 542898 104486 543134
rect 104570 542898 104806 543134
rect 123930 543218 124166 543454
rect 124250 543218 124486 543454
rect 124570 543218 124806 543454
rect 123930 542898 124166 543134
rect 124250 542898 124486 543134
rect 124570 542898 124806 543134
rect 143930 543218 144166 543454
rect 144250 543218 144486 543454
rect 144570 543218 144806 543454
rect 143930 542898 144166 543134
rect 144250 542898 144486 543134
rect 144570 542898 144806 543134
rect 163930 543218 164166 543454
rect 164250 543218 164486 543454
rect 164570 543218 164806 543454
rect 163930 542898 164166 543134
rect 164250 542898 164486 543134
rect 164570 542898 164806 543134
rect 183930 543218 184166 543454
rect 184250 543218 184486 543454
rect 184570 543218 184806 543454
rect 183930 542898 184166 543134
rect 184250 542898 184486 543134
rect 184570 542898 184806 543134
rect 33930 511718 34166 511954
rect 34250 511718 34486 511954
rect 34570 511718 34806 511954
rect 33930 511398 34166 511634
rect 34250 511398 34486 511634
rect 34570 511398 34806 511634
rect 53930 511718 54166 511954
rect 54250 511718 54486 511954
rect 54570 511718 54806 511954
rect 53930 511398 54166 511634
rect 54250 511398 54486 511634
rect 54570 511398 54806 511634
rect 73930 511718 74166 511954
rect 74250 511718 74486 511954
rect 74570 511718 74806 511954
rect 73930 511398 74166 511634
rect 74250 511398 74486 511634
rect 74570 511398 74806 511634
rect 93930 511718 94166 511954
rect 94250 511718 94486 511954
rect 94570 511718 94806 511954
rect 93930 511398 94166 511634
rect 94250 511398 94486 511634
rect 94570 511398 94806 511634
rect 113930 511718 114166 511954
rect 114250 511718 114486 511954
rect 114570 511718 114806 511954
rect 113930 511398 114166 511634
rect 114250 511398 114486 511634
rect 114570 511398 114806 511634
rect 133930 511718 134166 511954
rect 134250 511718 134486 511954
rect 134570 511718 134806 511954
rect 133930 511398 134166 511634
rect 134250 511398 134486 511634
rect 134570 511398 134806 511634
rect 153930 511718 154166 511954
rect 154250 511718 154486 511954
rect 154570 511718 154806 511954
rect 153930 511398 154166 511634
rect 154250 511398 154486 511634
rect 154570 511398 154806 511634
rect 173930 511718 174166 511954
rect 174250 511718 174486 511954
rect 174570 511718 174806 511954
rect 173930 511398 174166 511634
rect 174250 511398 174486 511634
rect 174570 511398 174806 511634
rect 193930 511718 194166 511954
rect 194250 511718 194486 511954
rect 194570 511718 194806 511954
rect 193930 511398 194166 511634
rect 194250 511398 194486 511634
rect 194570 511398 194806 511634
rect 23930 507218 24166 507454
rect 24250 507218 24486 507454
rect 24570 507218 24806 507454
rect 23930 506898 24166 507134
rect 24250 506898 24486 507134
rect 24570 506898 24806 507134
rect 43930 507218 44166 507454
rect 44250 507218 44486 507454
rect 44570 507218 44806 507454
rect 43930 506898 44166 507134
rect 44250 506898 44486 507134
rect 44570 506898 44806 507134
rect 63930 507218 64166 507454
rect 64250 507218 64486 507454
rect 64570 507218 64806 507454
rect 63930 506898 64166 507134
rect 64250 506898 64486 507134
rect 64570 506898 64806 507134
rect 83930 507218 84166 507454
rect 84250 507218 84486 507454
rect 84570 507218 84806 507454
rect 83930 506898 84166 507134
rect 84250 506898 84486 507134
rect 84570 506898 84806 507134
rect 103930 507218 104166 507454
rect 104250 507218 104486 507454
rect 104570 507218 104806 507454
rect 103930 506898 104166 507134
rect 104250 506898 104486 507134
rect 104570 506898 104806 507134
rect 123930 507218 124166 507454
rect 124250 507218 124486 507454
rect 124570 507218 124806 507454
rect 123930 506898 124166 507134
rect 124250 506898 124486 507134
rect 124570 506898 124806 507134
rect 143930 507218 144166 507454
rect 144250 507218 144486 507454
rect 144570 507218 144806 507454
rect 143930 506898 144166 507134
rect 144250 506898 144486 507134
rect 144570 506898 144806 507134
rect 163930 507218 164166 507454
rect 164250 507218 164486 507454
rect 164570 507218 164806 507454
rect 163930 506898 164166 507134
rect 164250 506898 164486 507134
rect 164570 506898 164806 507134
rect 183930 507218 184166 507454
rect 184250 507218 184486 507454
rect 184570 507218 184806 507454
rect 183930 506898 184166 507134
rect 184250 506898 184486 507134
rect 184570 506898 184806 507134
rect 33930 475718 34166 475954
rect 34250 475718 34486 475954
rect 34570 475718 34806 475954
rect 33930 475398 34166 475634
rect 34250 475398 34486 475634
rect 34570 475398 34806 475634
rect 53930 475718 54166 475954
rect 54250 475718 54486 475954
rect 54570 475718 54806 475954
rect 53930 475398 54166 475634
rect 54250 475398 54486 475634
rect 54570 475398 54806 475634
rect 73930 475718 74166 475954
rect 74250 475718 74486 475954
rect 74570 475718 74806 475954
rect 73930 475398 74166 475634
rect 74250 475398 74486 475634
rect 74570 475398 74806 475634
rect 93930 475718 94166 475954
rect 94250 475718 94486 475954
rect 94570 475718 94806 475954
rect 93930 475398 94166 475634
rect 94250 475398 94486 475634
rect 94570 475398 94806 475634
rect 113930 475718 114166 475954
rect 114250 475718 114486 475954
rect 114570 475718 114806 475954
rect 113930 475398 114166 475634
rect 114250 475398 114486 475634
rect 114570 475398 114806 475634
rect 133930 475718 134166 475954
rect 134250 475718 134486 475954
rect 134570 475718 134806 475954
rect 133930 475398 134166 475634
rect 134250 475398 134486 475634
rect 134570 475398 134806 475634
rect 153930 475718 154166 475954
rect 154250 475718 154486 475954
rect 154570 475718 154806 475954
rect 153930 475398 154166 475634
rect 154250 475398 154486 475634
rect 154570 475398 154806 475634
rect 173930 475718 174166 475954
rect 174250 475718 174486 475954
rect 174570 475718 174806 475954
rect 173930 475398 174166 475634
rect 174250 475398 174486 475634
rect 174570 475398 174806 475634
rect 193930 475718 194166 475954
rect 194250 475718 194486 475954
rect 194570 475718 194806 475954
rect 193930 475398 194166 475634
rect 194250 475398 194486 475634
rect 194570 475398 194806 475634
rect 23930 471218 24166 471454
rect 24250 471218 24486 471454
rect 24570 471218 24806 471454
rect 23930 470898 24166 471134
rect 24250 470898 24486 471134
rect 24570 470898 24806 471134
rect 43930 471218 44166 471454
rect 44250 471218 44486 471454
rect 44570 471218 44806 471454
rect 43930 470898 44166 471134
rect 44250 470898 44486 471134
rect 44570 470898 44806 471134
rect 63930 471218 64166 471454
rect 64250 471218 64486 471454
rect 64570 471218 64806 471454
rect 63930 470898 64166 471134
rect 64250 470898 64486 471134
rect 64570 470898 64806 471134
rect 83930 471218 84166 471454
rect 84250 471218 84486 471454
rect 84570 471218 84806 471454
rect 83930 470898 84166 471134
rect 84250 470898 84486 471134
rect 84570 470898 84806 471134
rect 103930 471218 104166 471454
rect 104250 471218 104486 471454
rect 104570 471218 104806 471454
rect 103930 470898 104166 471134
rect 104250 470898 104486 471134
rect 104570 470898 104806 471134
rect 123930 471218 124166 471454
rect 124250 471218 124486 471454
rect 124570 471218 124806 471454
rect 123930 470898 124166 471134
rect 124250 470898 124486 471134
rect 124570 470898 124806 471134
rect 143930 471218 144166 471454
rect 144250 471218 144486 471454
rect 144570 471218 144806 471454
rect 143930 470898 144166 471134
rect 144250 470898 144486 471134
rect 144570 470898 144806 471134
rect 163930 471218 164166 471454
rect 164250 471218 164486 471454
rect 164570 471218 164806 471454
rect 163930 470898 164166 471134
rect 164250 470898 164486 471134
rect 164570 470898 164806 471134
rect 183930 471218 184166 471454
rect 184250 471218 184486 471454
rect 184570 471218 184806 471454
rect 183930 470898 184166 471134
rect 184250 470898 184486 471134
rect 184570 470898 184806 471134
rect 33930 439718 34166 439954
rect 34250 439718 34486 439954
rect 34570 439718 34806 439954
rect 33930 439398 34166 439634
rect 34250 439398 34486 439634
rect 34570 439398 34806 439634
rect 53930 439718 54166 439954
rect 54250 439718 54486 439954
rect 54570 439718 54806 439954
rect 53930 439398 54166 439634
rect 54250 439398 54486 439634
rect 54570 439398 54806 439634
rect 73930 439718 74166 439954
rect 74250 439718 74486 439954
rect 74570 439718 74806 439954
rect 73930 439398 74166 439634
rect 74250 439398 74486 439634
rect 74570 439398 74806 439634
rect 93930 439718 94166 439954
rect 94250 439718 94486 439954
rect 94570 439718 94806 439954
rect 93930 439398 94166 439634
rect 94250 439398 94486 439634
rect 94570 439398 94806 439634
rect 113930 439718 114166 439954
rect 114250 439718 114486 439954
rect 114570 439718 114806 439954
rect 113930 439398 114166 439634
rect 114250 439398 114486 439634
rect 114570 439398 114806 439634
rect 133930 439718 134166 439954
rect 134250 439718 134486 439954
rect 134570 439718 134806 439954
rect 133930 439398 134166 439634
rect 134250 439398 134486 439634
rect 134570 439398 134806 439634
rect 153930 439718 154166 439954
rect 154250 439718 154486 439954
rect 154570 439718 154806 439954
rect 153930 439398 154166 439634
rect 154250 439398 154486 439634
rect 154570 439398 154806 439634
rect 173930 439718 174166 439954
rect 174250 439718 174486 439954
rect 174570 439718 174806 439954
rect 173930 439398 174166 439634
rect 174250 439398 174486 439634
rect 174570 439398 174806 439634
rect 193930 439718 194166 439954
rect 194250 439718 194486 439954
rect 194570 439718 194806 439954
rect 193930 439398 194166 439634
rect 194250 439398 194486 439634
rect 194570 439398 194806 439634
rect 23930 435218 24166 435454
rect 24250 435218 24486 435454
rect 24570 435218 24806 435454
rect 23930 434898 24166 435134
rect 24250 434898 24486 435134
rect 24570 434898 24806 435134
rect 43930 435218 44166 435454
rect 44250 435218 44486 435454
rect 44570 435218 44806 435454
rect 43930 434898 44166 435134
rect 44250 434898 44486 435134
rect 44570 434898 44806 435134
rect 63930 435218 64166 435454
rect 64250 435218 64486 435454
rect 64570 435218 64806 435454
rect 63930 434898 64166 435134
rect 64250 434898 64486 435134
rect 64570 434898 64806 435134
rect 83930 435218 84166 435454
rect 84250 435218 84486 435454
rect 84570 435218 84806 435454
rect 83930 434898 84166 435134
rect 84250 434898 84486 435134
rect 84570 434898 84806 435134
rect 103930 435218 104166 435454
rect 104250 435218 104486 435454
rect 104570 435218 104806 435454
rect 103930 434898 104166 435134
rect 104250 434898 104486 435134
rect 104570 434898 104806 435134
rect 123930 435218 124166 435454
rect 124250 435218 124486 435454
rect 124570 435218 124806 435454
rect 123930 434898 124166 435134
rect 124250 434898 124486 435134
rect 124570 434898 124806 435134
rect 143930 435218 144166 435454
rect 144250 435218 144486 435454
rect 144570 435218 144806 435454
rect 143930 434898 144166 435134
rect 144250 434898 144486 435134
rect 144570 434898 144806 435134
rect 163930 435218 164166 435454
rect 164250 435218 164486 435454
rect 164570 435218 164806 435454
rect 163930 434898 164166 435134
rect 164250 434898 164486 435134
rect 164570 434898 164806 435134
rect 183930 435218 184166 435454
rect 184250 435218 184486 435454
rect 184570 435218 184806 435454
rect 183930 434898 184166 435134
rect 184250 434898 184486 435134
rect 184570 434898 184806 435134
rect 33930 403718 34166 403954
rect 34250 403718 34486 403954
rect 34570 403718 34806 403954
rect 33930 403398 34166 403634
rect 34250 403398 34486 403634
rect 34570 403398 34806 403634
rect 53930 403718 54166 403954
rect 54250 403718 54486 403954
rect 54570 403718 54806 403954
rect 53930 403398 54166 403634
rect 54250 403398 54486 403634
rect 54570 403398 54806 403634
rect 73930 403718 74166 403954
rect 74250 403718 74486 403954
rect 74570 403718 74806 403954
rect 73930 403398 74166 403634
rect 74250 403398 74486 403634
rect 74570 403398 74806 403634
rect 93930 403718 94166 403954
rect 94250 403718 94486 403954
rect 94570 403718 94806 403954
rect 93930 403398 94166 403634
rect 94250 403398 94486 403634
rect 94570 403398 94806 403634
rect 113930 403718 114166 403954
rect 114250 403718 114486 403954
rect 114570 403718 114806 403954
rect 113930 403398 114166 403634
rect 114250 403398 114486 403634
rect 114570 403398 114806 403634
rect 133930 403718 134166 403954
rect 134250 403718 134486 403954
rect 134570 403718 134806 403954
rect 133930 403398 134166 403634
rect 134250 403398 134486 403634
rect 134570 403398 134806 403634
rect 153930 403718 154166 403954
rect 154250 403718 154486 403954
rect 154570 403718 154806 403954
rect 153930 403398 154166 403634
rect 154250 403398 154486 403634
rect 154570 403398 154806 403634
rect 173930 403718 174166 403954
rect 174250 403718 174486 403954
rect 174570 403718 174806 403954
rect 173930 403398 174166 403634
rect 174250 403398 174486 403634
rect 174570 403398 174806 403634
rect 193930 403718 194166 403954
rect 194250 403718 194486 403954
rect 194570 403718 194806 403954
rect 193930 403398 194166 403634
rect 194250 403398 194486 403634
rect 194570 403398 194806 403634
rect 23930 399218 24166 399454
rect 24250 399218 24486 399454
rect 24570 399218 24806 399454
rect 23930 398898 24166 399134
rect 24250 398898 24486 399134
rect 24570 398898 24806 399134
rect 43930 399218 44166 399454
rect 44250 399218 44486 399454
rect 44570 399218 44806 399454
rect 43930 398898 44166 399134
rect 44250 398898 44486 399134
rect 44570 398898 44806 399134
rect 63930 399218 64166 399454
rect 64250 399218 64486 399454
rect 64570 399218 64806 399454
rect 63930 398898 64166 399134
rect 64250 398898 64486 399134
rect 64570 398898 64806 399134
rect 83930 399218 84166 399454
rect 84250 399218 84486 399454
rect 84570 399218 84806 399454
rect 83930 398898 84166 399134
rect 84250 398898 84486 399134
rect 84570 398898 84806 399134
rect 103930 399218 104166 399454
rect 104250 399218 104486 399454
rect 104570 399218 104806 399454
rect 103930 398898 104166 399134
rect 104250 398898 104486 399134
rect 104570 398898 104806 399134
rect 123930 399218 124166 399454
rect 124250 399218 124486 399454
rect 124570 399218 124806 399454
rect 123930 398898 124166 399134
rect 124250 398898 124486 399134
rect 124570 398898 124806 399134
rect 143930 399218 144166 399454
rect 144250 399218 144486 399454
rect 144570 399218 144806 399454
rect 143930 398898 144166 399134
rect 144250 398898 144486 399134
rect 144570 398898 144806 399134
rect 163930 399218 164166 399454
rect 164250 399218 164486 399454
rect 164570 399218 164806 399454
rect 163930 398898 164166 399134
rect 164250 398898 164486 399134
rect 164570 398898 164806 399134
rect 183930 399218 184166 399454
rect 184250 399218 184486 399454
rect 184570 399218 184806 399454
rect 183930 398898 184166 399134
rect 184250 398898 184486 399134
rect 184570 398898 184806 399134
rect 33930 367718 34166 367954
rect 34250 367718 34486 367954
rect 34570 367718 34806 367954
rect 33930 367398 34166 367634
rect 34250 367398 34486 367634
rect 34570 367398 34806 367634
rect 53930 367718 54166 367954
rect 54250 367718 54486 367954
rect 54570 367718 54806 367954
rect 53930 367398 54166 367634
rect 54250 367398 54486 367634
rect 54570 367398 54806 367634
rect 73930 367718 74166 367954
rect 74250 367718 74486 367954
rect 74570 367718 74806 367954
rect 73930 367398 74166 367634
rect 74250 367398 74486 367634
rect 74570 367398 74806 367634
rect 93930 367718 94166 367954
rect 94250 367718 94486 367954
rect 94570 367718 94806 367954
rect 93930 367398 94166 367634
rect 94250 367398 94486 367634
rect 94570 367398 94806 367634
rect 113930 367718 114166 367954
rect 114250 367718 114486 367954
rect 114570 367718 114806 367954
rect 113930 367398 114166 367634
rect 114250 367398 114486 367634
rect 114570 367398 114806 367634
rect 133930 367718 134166 367954
rect 134250 367718 134486 367954
rect 134570 367718 134806 367954
rect 133930 367398 134166 367634
rect 134250 367398 134486 367634
rect 134570 367398 134806 367634
rect 153930 367718 154166 367954
rect 154250 367718 154486 367954
rect 154570 367718 154806 367954
rect 153930 367398 154166 367634
rect 154250 367398 154486 367634
rect 154570 367398 154806 367634
rect 173930 367718 174166 367954
rect 174250 367718 174486 367954
rect 174570 367718 174806 367954
rect 173930 367398 174166 367634
rect 174250 367398 174486 367634
rect 174570 367398 174806 367634
rect 193930 367718 194166 367954
rect 194250 367718 194486 367954
rect 194570 367718 194806 367954
rect 193930 367398 194166 367634
rect 194250 367398 194486 367634
rect 194570 367398 194806 367634
rect 23930 363218 24166 363454
rect 24250 363218 24486 363454
rect 24570 363218 24806 363454
rect 23930 362898 24166 363134
rect 24250 362898 24486 363134
rect 24570 362898 24806 363134
rect 43930 363218 44166 363454
rect 44250 363218 44486 363454
rect 44570 363218 44806 363454
rect 43930 362898 44166 363134
rect 44250 362898 44486 363134
rect 44570 362898 44806 363134
rect 63930 363218 64166 363454
rect 64250 363218 64486 363454
rect 64570 363218 64806 363454
rect 63930 362898 64166 363134
rect 64250 362898 64486 363134
rect 64570 362898 64806 363134
rect 83930 363218 84166 363454
rect 84250 363218 84486 363454
rect 84570 363218 84806 363454
rect 83930 362898 84166 363134
rect 84250 362898 84486 363134
rect 84570 362898 84806 363134
rect 103930 363218 104166 363454
rect 104250 363218 104486 363454
rect 104570 363218 104806 363454
rect 103930 362898 104166 363134
rect 104250 362898 104486 363134
rect 104570 362898 104806 363134
rect 123930 363218 124166 363454
rect 124250 363218 124486 363454
rect 124570 363218 124806 363454
rect 123930 362898 124166 363134
rect 124250 362898 124486 363134
rect 124570 362898 124806 363134
rect 143930 363218 144166 363454
rect 144250 363218 144486 363454
rect 144570 363218 144806 363454
rect 143930 362898 144166 363134
rect 144250 362898 144486 363134
rect 144570 362898 144806 363134
rect 163930 363218 164166 363454
rect 164250 363218 164486 363454
rect 164570 363218 164806 363454
rect 163930 362898 164166 363134
rect 164250 362898 164486 363134
rect 164570 362898 164806 363134
rect 183930 363218 184166 363454
rect 184250 363218 184486 363454
rect 184570 363218 184806 363454
rect 183930 362898 184166 363134
rect 184250 362898 184486 363134
rect 184570 362898 184806 363134
rect 33930 295718 34166 295954
rect 34250 295718 34486 295954
rect 34570 295718 34806 295954
rect 33930 295398 34166 295634
rect 34250 295398 34486 295634
rect 34570 295398 34806 295634
rect 53930 295718 54166 295954
rect 54250 295718 54486 295954
rect 54570 295718 54806 295954
rect 53930 295398 54166 295634
rect 54250 295398 54486 295634
rect 54570 295398 54806 295634
rect 73930 295718 74166 295954
rect 74250 295718 74486 295954
rect 74570 295718 74806 295954
rect 73930 295398 74166 295634
rect 74250 295398 74486 295634
rect 74570 295398 74806 295634
rect 93930 295718 94166 295954
rect 94250 295718 94486 295954
rect 94570 295718 94806 295954
rect 93930 295398 94166 295634
rect 94250 295398 94486 295634
rect 94570 295398 94806 295634
rect 113930 295718 114166 295954
rect 114250 295718 114486 295954
rect 114570 295718 114806 295954
rect 113930 295398 114166 295634
rect 114250 295398 114486 295634
rect 114570 295398 114806 295634
rect 133930 295718 134166 295954
rect 134250 295718 134486 295954
rect 134570 295718 134806 295954
rect 133930 295398 134166 295634
rect 134250 295398 134486 295634
rect 134570 295398 134806 295634
rect 153930 295718 154166 295954
rect 154250 295718 154486 295954
rect 154570 295718 154806 295954
rect 153930 295398 154166 295634
rect 154250 295398 154486 295634
rect 154570 295398 154806 295634
rect 173930 295718 174166 295954
rect 174250 295718 174486 295954
rect 174570 295718 174806 295954
rect 173930 295398 174166 295634
rect 174250 295398 174486 295634
rect 174570 295398 174806 295634
rect 193930 295718 194166 295954
rect 194250 295718 194486 295954
rect 194570 295718 194806 295954
rect 193930 295398 194166 295634
rect 194250 295398 194486 295634
rect 194570 295398 194806 295634
rect 23930 291218 24166 291454
rect 24250 291218 24486 291454
rect 24570 291218 24806 291454
rect 23930 290898 24166 291134
rect 24250 290898 24486 291134
rect 24570 290898 24806 291134
rect 43930 291218 44166 291454
rect 44250 291218 44486 291454
rect 44570 291218 44806 291454
rect 43930 290898 44166 291134
rect 44250 290898 44486 291134
rect 44570 290898 44806 291134
rect 63930 291218 64166 291454
rect 64250 291218 64486 291454
rect 64570 291218 64806 291454
rect 63930 290898 64166 291134
rect 64250 290898 64486 291134
rect 64570 290898 64806 291134
rect 83930 291218 84166 291454
rect 84250 291218 84486 291454
rect 84570 291218 84806 291454
rect 83930 290898 84166 291134
rect 84250 290898 84486 291134
rect 84570 290898 84806 291134
rect 103930 291218 104166 291454
rect 104250 291218 104486 291454
rect 104570 291218 104806 291454
rect 103930 290898 104166 291134
rect 104250 290898 104486 291134
rect 104570 290898 104806 291134
rect 123930 291218 124166 291454
rect 124250 291218 124486 291454
rect 124570 291218 124806 291454
rect 123930 290898 124166 291134
rect 124250 290898 124486 291134
rect 124570 290898 124806 291134
rect 143930 291218 144166 291454
rect 144250 291218 144486 291454
rect 144570 291218 144806 291454
rect 143930 290898 144166 291134
rect 144250 290898 144486 291134
rect 144570 290898 144806 291134
rect 163930 291218 164166 291454
rect 164250 291218 164486 291454
rect 164570 291218 164806 291454
rect 163930 290898 164166 291134
rect 164250 290898 164486 291134
rect 164570 290898 164806 291134
rect 183930 291218 184166 291454
rect 184250 291218 184486 291454
rect 184570 291218 184806 291454
rect 183930 290898 184166 291134
rect 184250 290898 184486 291134
rect 184570 290898 184806 291134
rect 33930 259718 34166 259954
rect 34250 259718 34486 259954
rect 34570 259718 34806 259954
rect 33930 259398 34166 259634
rect 34250 259398 34486 259634
rect 34570 259398 34806 259634
rect 53930 259718 54166 259954
rect 54250 259718 54486 259954
rect 54570 259718 54806 259954
rect 53930 259398 54166 259634
rect 54250 259398 54486 259634
rect 54570 259398 54806 259634
rect 73930 259718 74166 259954
rect 74250 259718 74486 259954
rect 74570 259718 74806 259954
rect 73930 259398 74166 259634
rect 74250 259398 74486 259634
rect 74570 259398 74806 259634
rect 93930 259718 94166 259954
rect 94250 259718 94486 259954
rect 94570 259718 94806 259954
rect 93930 259398 94166 259634
rect 94250 259398 94486 259634
rect 94570 259398 94806 259634
rect 113930 259718 114166 259954
rect 114250 259718 114486 259954
rect 114570 259718 114806 259954
rect 113930 259398 114166 259634
rect 114250 259398 114486 259634
rect 114570 259398 114806 259634
rect 133930 259718 134166 259954
rect 134250 259718 134486 259954
rect 134570 259718 134806 259954
rect 133930 259398 134166 259634
rect 134250 259398 134486 259634
rect 134570 259398 134806 259634
rect 153930 259718 154166 259954
rect 154250 259718 154486 259954
rect 154570 259718 154806 259954
rect 153930 259398 154166 259634
rect 154250 259398 154486 259634
rect 154570 259398 154806 259634
rect 173930 259718 174166 259954
rect 174250 259718 174486 259954
rect 174570 259718 174806 259954
rect 173930 259398 174166 259634
rect 174250 259398 174486 259634
rect 174570 259398 174806 259634
rect 193930 259718 194166 259954
rect 194250 259718 194486 259954
rect 194570 259718 194806 259954
rect 193930 259398 194166 259634
rect 194250 259398 194486 259634
rect 194570 259398 194806 259634
rect 23930 255218 24166 255454
rect 24250 255218 24486 255454
rect 24570 255218 24806 255454
rect 23930 254898 24166 255134
rect 24250 254898 24486 255134
rect 24570 254898 24806 255134
rect 43930 255218 44166 255454
rect 44250 255218 44486 255454
rect 44570 255218 44806 255454
rect 43930 254898 44166 255134
rect 44250 254898 44486 255134
rect 44570 254898 44806 255134
rect 63930 255218 64166 255454
rect 64250 255218 64486 255454
rect 64570 255218 64806 255454
rect 63930 254898 64166 255134
rect 64250 254898 64486 255134
rect 64570 254898 64806 255134
rect 83930 255218 84166 255454
rect 84250 255218 84486 255454
rect 84570 255218 84806 255454
rect 83930 254898 84166 255134
rect 84250 254898 84486 255134
rect 84570 254898 84806 255134
rect 103930 255218 104166 255454
rect 104250 255218 104486 255454
rect 104570 255218 104806 255454
rect 103930 254898 104166 255134
rect 104250 254898 104486 255134
rect 104570 254898 104806 255134
rect 123930 255218 124166 255454
rect 124250 255218 124486 255454
rect 124570 255218 124806 255454
rect 123930 254898 124166 255134
rect 124250 254898 124486 255134
rect 124570 254898 124806 255134
rect 143930 255218 144166 255454
rect 144250 255218 144486 255454
rect 144570 255218 144806 255454
rect 143930 254898 144166 255134
rect 144250 254898 144486 255134
rect 144570 254898 144806 255134
rect 163930 255218 164166 255454
rect 164250 255218 164486 255454
rect 164570 255218 164806 255454
rect 163930 254898 164166 255134
rect 164250 254898 164486 255134
rect 164570 254898 164806 255134
rect 183930 255218 184166 255454
rect 184250 255218 184486 255454
rect 184570 255218 184806 255454
rect 183930 254898 184166 255134
rect 184250 254898 184486 255134
rect 184570 254898 184806 255134
rect 33930 223718 34166 223954
rect 34250 223718 34486 223954
rect 34570 223718 34806 223954
rect 33930 223398 34166 223634
rect 34250 223398 34486 223634
rect 34570 223398 34806 223634
rect 53930 223718 54166 223954
rect 54250 223718 54486 223954
rect 54570 223718 54806 223954
rect 53930 223398 54166 223634
rect 54250 223398 54486 223634
rect 54570 223398 54806 223634
rect 73930 223718 74166 223954
rect 74250 223718 74486 223954
rect 74570 223718 74806 223954
rect 73930 223398 74166 223634
rect 74250 223398 74486 223634
rect 74570 223398 74806 223634
rect 93930 223718 94166 223954
rect 94250 223718 94486 223954
rect 94570 223718 94806 223954
rect 93930 223398 94166 223634
rect 94250 223398 94486 223634
rect 94570 223398 94806 223634
rect 113930 223718 114166 223954
rect 114250 223718 114486 223954
rect 114570 223718 114806 223954
rect 113930 223398 114166 223634
rect 114250 223398 114486 223634
rect 114570 223398 114806 223634
rect 133930 223718 134166 223954
rect 134250 223718 134486 223954
rect 134570 223718 134806 223954
rect 133930 223398 134166 223634
rect 134250 223398 134486 223634
rect 134570 223398 134806 223634
rect 153930 223718 154166 223954
rect 154250 223718 154486 223954
rect 154570 223718 154806 223954
rect 153930 223398 154166 223634
rect 154250 223398 154486 223634
rect 154570 223398 154806 223634
rect 173930 223718 174166 223954
rect 174250 223718 174486 223954
rect 174570 223718 174806 223954
rect 173930 223398 174166 223634
rect 174250 223398 174486 223634
rect 174570 223398 174806 223634
rect 193930 223718 194166 223954
rect 194250 223718 194486 223954
rect 194570 223718 194806 223954
rect 193930 223398 194166 223634
rect 194250 223398 194486 223634
rect 194570 223398 194806 223634
rect 23930 219218 24166 219454
rect 24250 219218 24486 219454
rect 24570 219218 24806 219454
rect 23930 218898 24166 219134
rect 24250 218898 24486 219134
rect 24570 218898 24806 219134
rect 43930 219218 44166 219454
rect 44250 219218 44486 219454
rect 44570 219218 44806 219454
rect 43930 218898 44166 219134
rect 44250 218898 44486 219134
rect 44570 218898 44806 219134
rect 63930 219218 64166 219454
rect 64250 219218 64486 219454
rect 64570 219218 64806 219454
rect 63930 218898 64166 219134
rect 64250 218898 64486 219134
rect 64570 218898 64806 219134
rect 83930 219218 84166 219454
rect 84250 219218 84486 219454
rect 84570 219218 84806 219454
rect 83930 218898 84166 219134
rect 84250 218898 84486 219134
rect 84570 218898 84806 219134
rect 103930 219218 104166 219454
rect 104250 219218 104486 219454
rect 104570 219218 104806 219454
rect 103930 218898 104166 219134
rect 104250 218898 104486 219134
rect 104570 218898 104806 219134
rect 123930 219218 124166 219454
rect 124250 219218 124486 219454
rect 124570 219218 124806 219454
rect 123930 218898 124166 219134
rect 124250 218898 124486 219134
rect 124570 218898 124806 219134
rect 143930 219218 144166 219454
rect 144250 219218 144486 219454
rect 144570 219218 144806 219454
rect 143930 218898 144166 219134
rect 144250 218898 144486 219134
rect 144570 218898 144806 219134
rect 163930 219218 164166 219454
rect 164250 219218 164486 219454
rect 164570 219218 164806 219454
rect 163930 218898 164166 219134
rect 164250 218898 164486 219134
rect 164570 218898 164806 219134
rect 183930 219218 184166 219454
rect 184250 219218 184486 219454
rect 184570 219218 184806 219454
rect 183930 218898 184166 219134
rect 184250 218898 184486 219134
rect 184570 218898 184806 219134
rect 23930 183218 24166 183454
rect 24250 183218 24486 183454
rect 24570 183218 24806 183454
rect 23930 182898 24166 183134
rect 24250 182898 24486 183134
rect 24570 182898 24806 183134
rect 43930 183218 44166 183454
rect 44250 183218 44486 183454
rect 44570 183218 44806 183454
rect 43930 182898 44166 183134
rect 44250 182898 44486 183134
rect 44570 182898 44806 183134
rect 63930 183218 64166 183454
rect 64250 183218 64486 183454
rect 64570 183218 64806 183454
rect 63930 182898 64166 183134
rect 64250 182898 64486 183134
rect 64570 182898 64806 183134
rect 83930 183218 84166 183454
rect 84250 183218 84486 183454
rect 84570 183218 84806 183454
rect 83930 182898 84166 183134
rect 84250 182898 84486 183134
rect 84570 182898 84806 183134
rect 103930 183218 104166 183454
rect 104250 183218 104486 183454
rect 104570 183218 104806 183454
rect 103930 182898 104166 183134
rect 104250 182898 104486 183134
rect 104570 182898 104806 183134
rect 123930 183218 124166 183454
rect 124250 183218 124486 183454
rect 124570 183218 124806 183454
rect 123930 182898 124166 183134
rect 124250 182898 124486 183134
rect 124570 182898 124806 183134
rect 143930 183218 144166 183454
rect 144250 183218 144486 183454
rect 144570 183218 144806 183454
rect 143930 182898 144166 183134
rect 144250 182898 144486 183134
rect 144570 182898 144806 183134
rect 163930 183218 164166 183454
rect 164250 183218 164486 183454
rect 164570 183218 164806 183454
rect 163930 182898 164166 183134
rect 164250 182898 164486 183134
rect 164570 182898 164806 183134
rect 183930 183218 184166 183454
rect 184250 183218 184486 183454
rect 184570 183218 184806 183454
rect 183930 182898 184166 183134
rect 184250 182898 184486 183134
rect 184570 182898 184806 183134
rect 33930 151718 34166 151954
rect 34250 151718 34486 151954
rect 34570 151718 34806 151954
rect 33930 151398 34166 151634
rect 34250 151398 34486 151634
rect 34570 151398 34806 151634
rect 53930 151718 54166 151954
rect 54250 151718 54486 151954
rect 54570 151718 54806 151954
rect 53930 151398 54166 151634
rect 54250 151398 54486 151634
rect 54570 151398 54806 151634
rect 73930 151718 74166 151954
rect 74250 151718 74486 151954
rect 74570 151718 74806 151954
rect 73930 151398 74166 151634
rect 74250 151398 74486 151634
rect 74570 151398 74806 151634
rect 93930 151718 94166 151954
rect 94250 151718 94486 151954
rect 94570 151718 94806 151954
rect 93930 151398 94166 151634
rect 94250 151398 94486 151634
rect 94570 151398 94806 151634
rect 113930 151718 114166 151954
rect 114250 151718 114486 151954
rect 114570 151718 114806 151954
rect 113930 151398 114166 151634
rect 114250 151398 114486 151634
rect 114570 151398 114806 151634
rect 133930 151718 134166 151954
rect 134250 151718 134486 151954
rect 134570 151718 134806 151954
rect 133930 151398 134166 151634
rect 134250 151398 134486 151634
rect 134570 151398 134806 151634
rect 153930 151718 154166 151954
rect 154250 151718 154486 151954
rect 154570 151718 154806 151954
rect 153930 151398 154166 151634
rect 154250 151398 154486 151634
rect 154570 151398 154806 151634
rect 173930 151718 174166 151954
rect 174250 151718 174486 151954
rect 174570 151718 174806 151954
rect 173930 151398 174166 151634
rect 174250 151398 174486 151634
rect 174570 151398 174806 151634
rect 193930 151718 194166 151954
rect 194250 151718 194486 151954
rect 194570 151718 194806 151954
rect 193930 151398 194166 151634
rect 194250 151398 194486 151634
rect 194570 151398 194806 151634
rect 23930 147218 24166 147454
rect 24250 147218 24486 147454
rect 24570 147218 24806 147454
rect 23930 146898 24166 147134
rect 24250 146898 24486 147134
rect 24570 146898 24806 147134
rect 43930 147218 44166 147454
rect 44250 147218 44486 147454
rect 44570 147218 44806 147454
rect 43930 146898 44166 147134
rect 44250 146898 44486 147134
rect 44570 146898 44806 147134
rect 63930 147218 64166 147454
rect 64250 147218 64486 147454
rect 64570 147218 64806 147454
rect 63930 146898 64166 147134
rect 64250 146898 64486 147134
rect 64570 146898 64806 147134
rect 83930 147218 84166 147454
rect 84250 147218 84486 147454
rect 84570 147218 84806 147454
rect 83930 146898 84166 147134
rect 84250 146898 84486 147134
rect 84570 146898 84806 147134
rect 103930 147218 104166 147454
rect 104250 147218 104486 147454
rect 104570 147218 104806 147454
rect 103930 146898 104166 147134
rect 104250 146898 104486 147134
rect 104570 146898 104806 147134
rect 123930 147218 124166 147454
rect 124250 147218 124486 147454
rect 124570 147218 124806 147454
rect 123930 146898 124166 147134
rect 124250 146898 124486 147134
rect 124570 146898 124806 147134
rect 143930 147218 144166 147454
rect 144250 147218 144486 147454
rect 144570 147218 144806 147454
rect 143930 146898 144166 147134
rect 144250 146898 144486 147134
rect 144570 146898 144806 147134
rect 163930 147218 164166 147454
rect 164250 147218 164486 147454
rect 164570 147218 164806 147454
rect 163930 146898 164166 147134
rect 164250 146898 164486 147134
rect 164570 146898 164806 147134
rect 183930 147218 184166 147454
rect 184250 147218 184486 147454
rect 184570 147218 184806 147454
rect 183930 146898 184166 147134
rect 184250 146898 184486 147134
rect 184570 146898 184806 147134
rect 33930 115718 34166 115954
rect 34250 115718 34486 115954
rect 34570 115718 34806 115954
rect 33930 115398 34166 115634
rect 34250 115398 34486 115634
rect 34570 115398 34806 115634
rect 53930 115718 54166 115954
rect 54250 115718 54486 115954
rect 54570 115718 54806 115954
rect 53930 115398 54166 115634
rect 54250 115398 54486 115634
rect 54570 115398 54806 115634
rect 73930 115718 74166 115954
rect 74250 115718 74486 115954
rect 74570 115718 74806 115954
rect 73930 115398 74166 115634
rect 74250 115398 74486 115634
rect 74570 115398 74806 115634
rect 93930 115718 94166 115954
rect 94250 115718 94486 115954
rect 94570 115718 94806 115954
rect 93930 115398 94166 115634
rect 94250 115398 94486 115634
rect 94570 115398 94806 115634
rect 113930 115718 114166 115954
rect 114250 115718 114486 115954
rect 114570 115718 114806 115954
rect 113930 115398 114166 115634
rect 114250 115398 114486 115634
rect 114570 115398 114806 115634
rect 133930 115718 134166 115954
rect 134250 115718 134486 115954
rect 134570 115718 134806 115954
rect 133930 115398 134166 115634
rect 134250 115398 134486 115634
rect 134570 115398 134806 115634
rect 153930 115718 154166 115954
rect 154250 115718 154486 115954
rect 154570 115718 154806 115954
rect 153930 115398 154166 115634
rect 154250 115398 154486 115634
rect 154570 115398 154806 115634
rect 173930 115718 174166 115954
rect 174250 115718 174486 115954
rect 174570 115718 174806 115954
rect 173930 115398 174166 115634
rect 174250 115398 174486 115634
rect 174570 115398 174806 115634
rect 193930 115718 194166 115954
rect 194250 115718 194486 115954
rect 194570 115718 194806 115954
rect 193930 115398 194166 115634
rect 194250 115398 194486 115634
rect 194570 115398 194806 115634
rect 23930 111218 24166 111454
rect 24250 111218 24486 111454
rect 24570 111218 24806 111454
rect 23930 110898 24166 111134
rect 24250 110898 24486 111134
rect 24570 110898 24806 111134
rect 43930 111218 44166 111454
rect 44250 111218 44486 111454
rect 44570 111218 44806 111454
rect 43930 110898 44166 111134
rect 44250 110898 44486 111134
rect 44570 110898 44806 111134
rect 63930 111218 64166 111454
rect 64250 111218 64486 111454
rect 64570 111218 64806 111454
rect 63930 110898 64166 111134
rect 64250 110898 64486 111134
rect 64570 110898 64806 111134
rect 83930 111218 84166 111454
rect 84250 111218 84486 111454
rect 84570 111218 84806 111454
rect 83930 110898 84166 111134
rect 84250 110898 84486 111134
rect 84570 110898 84806 111134
rect 103930 111218 104166 111454
rect 104250 111218 104486 111454
rect 104570 111218 104806 111454
rect 103930 110898 104166 111134
rect 104250 110898 104486 111134
rect 104570 110898 104806 111134
rect 123930 111218 124166 111454
rect 124250 111218 124486 111454
rect 124570 111218 124806 111454
rect 123930 110898 124166 111134
rect 124250 110898 124486 111134
rect 124570 110898 124806 111134
rect 143930 111218 144166 111454
rect 144250 111218 144486 111454
rect 144570 111218 144806 111454
rect 143930 110898 144166 111134
rect 144250 110898 144486 111134
rect 144570 110898 144806 111134
rect 163930 111218 164166 111454
rect 164250 111218 164486 111454
rect 164570 111218 164806 111454
rect 163930 110898 164166 111134
rect 164250 110898 164486 111134
rect 164570 110898 164806 111134
rect 183930 111218 184166 111454
rect 184250 111218 184486 111454
rect 184570 111218 184806 111454
rect 183930 110898 184166 111134
rect 184250 110898 184486 111134
rect 184570 110898 184806 111134
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 79610 43718 79846 43954
rect 79610 43398 79846 43634
rect 64250 39218 64486 39454
rect 64250 38898 64486 39134
rect 94970 39218 95206 39454
rect 94970 38898 95206 39134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 313930 691718 314166 691954
rect 314250 691718 314486 691954
rect 314570 691718 314806 691954
rect 313930 691398 314166 691634
rect 314250 691398 314486 691634
rect 314570 691398 314806 691634
rect 333930 691718 334166 691954
rect 334250 691718 334486 691954
rect 334570 691718 334806 691954
rect 333930 691398 334166 691634
rect 334250 691398 334486 691634
rect 334570 691398 334806 691634
rect 353930 691718 354166 691954
rect 354250 691718 354486 691954
rect 354570 691718 354806 691954
rect 353930 691398 354166 691634
rect 354250 691398 354486 691634
rect 354570 691398 354806 691634
rect 373930 691718 374166 691954
rect 374250 691718 374486 691954
rect 374570 691718 374806 691954
rect 373930 691398 374166 691634
rect 374250 691398 374486 691634
rect 374570 691398 374806 691634
rect 393930 691718 394166 691954
rect 394250 691718 394486 691954
rect 394570 691718 394806 691954
rect 393930 691398 394166 691634
rect 394250 691398 394486 691634
rect 394570 691398 394806 691634
rect 413930 691718 414166 691954
rect 414250 691718 414486 691954
rect 414570 691718 414806 691954
rect 413930 691398 414166 691634
rect 414250 691398 414486 691634
rect 414570 691398 414806 691634
rect 433930 691718 434166 691954
rect 434250 691718 434486 691954
rect 434570 691718 434806 691954
rect 433930 691398 434166 691634
rect 434250 691398 434486 691634
rect 434570 691398 434806 691634
rect 453930 691718 454166 691954
rect 454250 691718 454486 691954
rect 454570 691718 454806 691954
rect 453930 691398 454166 691634
rect 454250 691398 454486 691634
rect 454570 691398 454806 691634
rect 473930 691718 474166 691954
rect 474250 691718 474486 691954
rect 474570 691718 474806 691954
rect 473930 691398 474166 691634
rect 474250 691398 474486 691634
rect 474570 691398 474806 691634
rect 303930 687218 304166 687454
rect 304250 687218 304486 687454
rect 304570 687218 304806 687454
rect 303930 686898 304166 687134
rect 304250 686898 304486 687134
rect 304570 686898 304806 687134
rect 323930 687218 324166 687454
rect 324250 687218 324486 687454
rect 324570 687218 324806 687454
rect 323930 686898 324166 687134
rect 324250 686898 324486 687134
rect 324570 686898 324806 687134
rect 343930 687218 344166 687454
rect 344250 687218 344486 687454
rect 344570 687218 344806 687454
rect 343930 686898 344166 687134
rect 344250 686898 344486 687134
rect 344570 686898 344806 687134
rect 363930 687218 364166 687454
rect 364250 687218 364486 687454
rect 364570 687218 364806 687454
rect 363930 686898 364166 687134
rect 364250 686898 364486 687134
rect 364570 686898 364806 687134
rect 383930 687218 384166 687454
rect 384250 687218 384486 687454
rect 384570 687218 384806 687454
rect 383930 686898 384166 687134
rect 384250 686898 384486 687134
rect 384570 686898 384806 687134
rect 403930 687218 404166 687454
rect 404250 687218 404486 687454
rect 404570 687218 404806 687454
rect 403930 686898 404166 687134
rect 404250 686898 404486 687134
rect 404570 686898 404806 687134
rect 423930 687218 424166 687454
rect 424250 687218 424486 687454
rect 424570 687218 424806 687454
rect 423930 686898 424166 687134
rect 424250 686898 424486 687134
rect 424570 686898 424806 687134
rect 443930 687218 444166 687454
rect 444250 687218 444486 687454
rect 444570 687218 444806 687454
rect 443930 686898 444166 687134
rect 444250 686898 444486 687134
rect 444570 686898 444806 687134
rect 463930 687218 464166 687454
rect 464250 687218 464486 687454
rect 464570 687218 464806 687454
rect 463930 686898 464166 687134
rect 464250 686898 464486 687134
rect 464570 686898 464806 687134
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 313930 655718 314166 655954
rect 314250 655718 314486 655954
rect 314570 655718 314806 655954
rect 313930 655398 314166 655634
rect 314250 655398 314486 655634
rect 314570 655398 314806 655634
rect 333930 655718 334166 655954
rect 334250 655718 334486 655954
rect 334570 655718 334806 655954
rect 333930 655398 334166 655634
rect 334250 655398 334486 655634
rect 334570 655398 334806 655634
rect 353930 655718 354166 655954
rect 354250 655718 354486 655954
rect 354570 655718 354806 655954
rect 353930 655398 354166 655634
rect 354250 655398 354486 655634
rect 354570 655398 354806 655634
rect 373930 655718 374166 655954
rect 374250 655718 374486 655954
rect 374570 655718 374806 655954
rect 373930 655398 374166 655634
rect 374250 655398 374486 655634
rect 374570 655398 374806 655634
rect 393930 655718 394166 655954
rect 394250 655718 394486 655954
rect 394570 655718 394806 655954
rect 393930 655398 394166 655634
rect 394250 655398 394486 655634
rect 394570 655398 394806 655634
rect 413930 655718 414166 655954
rect 414250 655718 414486 655954
rect 414570 655718 414806 655954
rect 413930 655398 414166 655634
rect 414250 655398 414486 655634
rect 414570 655398 414806 655634
rect 433930 655718 434166 655954
rect 434250 655718 434486 655954
rect 434570 655718 434806 655954
rect 433930 655398 434166 655634
rect 434250 655398 434486 655634
rect 434570 655398 434806 655634
rect 453930 655718 454166 655954
rect 454250 655718 454486 655954
rect 454570 655718 454806 655954
rect 453930 655398 454166 655634
rect 454250 655398 454486 655634
rect 454570 655398 454806 655634
rect 473930 655718 474166 655954
rect 474250 655718 474486 655954
rect 474570 655718 474806 655954
rect 473930 655398 474166 655634
rect 474250 655398 474486 655634
rect 474570 655398 474806 655634
rect 303930 651218 304166 651454
rect 304250 651218 304486 651454
rect 304570 651218 304806 651454
rect 303930 650898 304166 651134
rect 304250 650898 304486 651134
rect 304570 650898 304806 651134
rect 323930 651218 324166 651454
rect 324250 651218 324486 651454
rect 324570 651218 324806 651454
rect 323930 650898 324166 651134
rect 324250 650898 324486 651134
rect 324570 650898 324806 651134
rect 343930 651218 344166 651454
rect 344250 651218 344486 651454
rect 344570 651218 344806 651454
rect 343930 650898 344166 651134
rect 344250 650898 344486 651134
rect 344570 650898 344806 651134
rect 363930 651218 364166 651454
rect 364250 651218 364486 651454
rect 364570 651218 364806 651454
rect 363930 650898 364166 651134
rect 364250 650898 364486 651134
rect 364570 650898 364806 651134
rect 383930 651218 384166 651454
rect 384250 651218 384486 651454
rect 384570 651218 384806 651454
rect 383930 650898 384166 651134
rect 384250 650898 384486 651134
rect 384570 650898 384806 651134
rect 403930 651218 404166 651454
rect 404250 651218 404486 651454
rect 404570 651218 404806 651454
rect 403930 650898 404166 651134
rect 404250 650898 404486 651134
rect 404570 650898 404806 651134
rect 423930 651218 424166 651454
rect 424250 651218 424486 651454
rect 424570 651218 424806 651454
rect 423930 650898 424166 651134
rect 424250 650898 424486 651134
rect 424570 650898 424806 651134
rect 443930 651218 444166 651454
rect 444250 651218 444486 651454
rect 444570 651218 444806 651454
rect 443930 650898 444166 651134
rect 444250 650898 444486 651134
rect 444570 650898 444806 651134
rect 463930 651218 464166 651454
rect 464250 651218 464486 651454
rect 464570 651218 464806 651454
rect 463930 650898 464166 651134
rect 464250 650898 464486 651134
rect 464570 650898 464806 651134
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 313930 619718 314166 619954
rect 314250 619718 314486 619954
rect 314570 619718 314806 619954
rect 313930 619398 314166 619634
rect 314250 619398 314486 619634
rect 314570 619398 314806 619634
rect 333930 619718 334166 619954
rect 334250 619718 334486 619954
rect 334570 619718 334806 619954
rect 333930 619398 334166 619634
rect 334250 619398 334486 619634
rect 334570 619398 334806 619634
rect 353930 619718 354166 619954
rect 354250 619718 354486 619954
rect 354570 619718 354806 619954
rect 353930 619398 354166 619634
rect 354250 619398 354486 619634
rect 354570 619398 354806 619634
rect 373930 619718 374166 619954
rect 374250 619718 374486 619954
rect 374570 619718 374806 619954
rect 373930 619398 374166 619634
rect 374250 619398 374486 619634
rect 374570 619398 374806 619634
rect 393930 619718 394166 619954
rect 394250 619718 394486 619954
rect 394570 619718 394806 619954
rect 393930 619398 394166 619634
rect 394250 619398 394486 619634
rect 394570 619398 394806 619634
rect 413930 619718 414166 619954
rect 414250 619718 414486 619954
rect 414570 619718 414806 619954
rect 413930 619398 414166 619634
rect 414250 619398 414486 619634
rect 414570 619398 414806 619634
rect 433930 619718 434166 619954
rect 434250 619718 434486 619954
rect 434570 619718 434806 619954
rect 433930 619398 434166 619634
rect 434250 619398 434486 619634
rect 434570 619398 434806 619634
rect 453930 619718 454166 619954
rect 454250 619718 454486 619954
rect 454570 619718 454806 619954
rect 453930 619398 454166 619634
rect 454250 619398 454486 619634
rect 454570 619398 454806 619634
rect 473930 619718 474166 619954
rect 474250 619718 474486 619954
rect 474570 619718 474806 619954
rect 473930 619398 474166 619634
rect 474250 619398 474486 619634
rect 474570 619398 474806 619634
rect 303930 615218 304166 615454
rect 304250 615218 304486 615454
rect 304570 615218 304806 615454
rect 303930 614898 304166 615134
rect 304250 614898 304486 615134
rect 304570 614898 304806 615134
rect 323930 615218 324166 615454
rect 324250 615218 324486 615454
rect 324570 615218 324806 615454
rect 323930 614898 324166 615134
rect 324250 614898 324486 615134
rect 324570 614898 324806 615134
rect 343930 615218 344166 615454
rect 344250 615218 344486 615454
rect 344570 615218 344806 615454
rect 343930 614898 344166 615134
rect 344250 614898 344486 615134
rect 344570 614898 344806 615134
rect 363930 615218 364166 615454
rect 364250 615218 364486 615454
rect 364570 615218 364806 615454
rect 363930 614898 364166 615134
rect 364250 614898 364486 615134
rect 364570 614898 364806 615134
rect 383930 615218 384166 615454
rect 384250 615218 384486 615454
rect 384570 615218 384806 615454
rect 383930 614898 384166 615134
rect 384250 614898 384486 615134
rect 384570 614898 384806 615134
rect 403930 615218 404166 615454
rect 404250 615218 404486 615454
rect 404570 615218 404806 615454
rect 403930 614898 404166 615134
rect 404250 614898 404486 615134
rect 404570 614898 404806 615134
rect 423930 615218 424166 615454
rect 424250 615218 424486 615454
rect 424570 615218 424806 615454
rect 423930 614898 424166 615134
rect 424250 614898 424486 615134
rect 424570 614898 424806 615134
rect 443930 615218 444166 615454
rect 444250 615218 444486 615454
rect 444570 615218 444806 615454
rect 443930 614898 444166 615134
rect 444250 614898 444486 615134
rect 444570 614898 444806 615134
rect 463930 615218 464166 615454
rect 464250 615218 464486 615454
rect 464570 615218 464806 615454
rect 463930 614898 464166 615134
rect 464250 614898 464486 615134
rect 464570 614898 464806 615134
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 313930 547718 314166 547954
rect 314250 547718 314486 547954
rect 314570 547718 314806 547954
rect 313930 547398 314166 547634
rect 314250 547398 314486 547634
rect 314570 547398 314806 547634
rect 333930 547718 334166 547954
rect 334250 547718 334486 547954
rect 334570 547718 334806 547954
rect 333930 547398 334166 547634
rect 334250 547398 334486 547634
rect 334570 547398 334806 547634
rect 353930 547718 354166 547954
rect 354250 547718 354486 547954
rect 354570 547718 354806 547954
rect 353930 547398 354166 547634
rect 354250 547398 354486 547634
rect 354570 547398 354806 547634
rect 373930 547718 374166 547954
rect 374250 547718 374486 547954
rect 374570 547718 374806 547954
rect 373930 547398 374166 547634
rect 374250 547398 374486 547634
rect 374570 547398 374806 547634
rect 393930 547718 394166 547954
rect 394250 547718 394486 547954
rect 394570 547718 394806 547954
rect 393930 547398 394166 547634
rect 394250 547398 394486 547634
rect 394570 547398 394806 547634
rect 413930 547718 414166 547954
rect 414250 547718 414486 547954
rect 414570 547718 414806 547954
rect 413930 547398 414166 547634
rect 414250 547398 414486 547634
rect 414570 547398 414806 547634
rect 433930 547718 434166 547954
rect 434250 547718 434486 547954
rect 434570 547718 434806 547954
rect 433930 547398 434166 547634
rect 434250 547398 434486 547634
rect 434570 547398 434806 547634
rect 453930 547718 454166 547954
rect 454250 547718 454486 547954
rect 454570 547718 454806 547954
rect 453930 547398 454166 547634
rect 454250 547398 454486 547634
rect 454570 547398 454806 547634
rect 473930 547718 474166 547954
rect 474250 547718 474486 547954
rect 474570 547718 474806 547954
rect 473930 547398 474166 547634
rect 474250 547398 474486 547634
rect 474570 547398 474806 547634
rect 303930 543218 304166 543454
rect 304250 543218 304486 543454
rect 304570 543218 304806 543454
rect 303930 542898 304166 543134
rect 304250 542898 304486 543134
rect 304570 542898 304806 543134
rect 323930 543218 324166 543454
rect 324250 543218 324486 543454
rect 324570 543218 324806 543454
rect 323930 542898 324166 543134
rect 324250 542898 324486 543134
rect 324570 542898 324806 543134
rect 343930 543218 344166 543454
rect 344250 543218 344486 543454
rect 344570 543218 344806 543454
rect 343930 542898 344166 543134
rect 344250 542898 344486 543134
rect 344570 542898 344806 543134
rect 363930 543218 364166 543454
rect 364250 543218 364486 543454
rect 364570 543218 364806 543454
rect 363930 542898 364166 543134
rect 364250 542898 364486 543134
rect 364570 542898 364806 543134
rect 383930 543218 384166 543454
rect 384250 543218 384486 543454
rect 384570 543218 384806 543454
rect 383930 542898 384166 543134
rect 384250 542898 384486 543134
rect 384570 542898 384806 543134
rect 403930 543218 404166 543454
rect 404250 543218 404486 543454
rect 404570 543218 404806 543454
rect 403930 542898 404166 543134
rect 404250 542898 404486 543134
rect 404570 542898 404806 543134
rect 423930 543218 424166 543454
rect 424250 543218 424486 543454
rect 424570 543218 424806 543454
rect 423930 542898 424166 543134
rect 424250 542898 424486 543134
rect 424570 542898 424806 543134
rect 443930 543218 444166 543454
rect 444250 543218 444486 543454
rect 444570 543218 444806 543454
rect 443930 542898 444166 543134
rect 444250 542898 444486 543134
rect 444570 542898 444806 543134
rect 463930 543218 464166 543454
rect 464250 543218 464486 543454
rect 464570 543218 464806 543454
rect 463930 542898 464166 543134
rect 464250 542898 464486 543134
rect 464570 542898 464806 543134
rect 313930 511718 314166 511954
rect 314250 511718 314486 511954
rect 314570 511718 314806 511954
rect 313930 511398 314166 511634
rect 314250 511398 314486 511634
rect 314570 511398 314806 511634
rect 333930 511718 334166 511954
rect 334250 511718 334486 511954
rect 334570 511718 334806 511954
rect 333930 511398 334166 511634
rect 334250 511398 334486 511634
rect 334570 511398 334806 511634
rect 353930 511718 354166 511954
rect 354250 511718 354486 511954
rect 354570 511718 354806 511954
rect 353930 511398 354166 511634
rect 354250 511398 354486 511634
rect 354570 511398 354806 511634
rect 373930 511718 374166 511954
rect 374250 511718 374486 511954
rect 374570 511718 374806 511954
rect 373930 511398 374166 511634
rect 374250 511398 374486 511634
rect 374570 511398 374806 511634
rect 393930 511718 394166 511954
rect 394250 511718 394486 511954
rect 394570 511718 394806 511954
rect 393930 511398 394166 511634
rect 394250 511398 394486 511634
rect 394570 511398 394806 511634
rect 413930 511718 414166 511954
rect 414250 511718 414486 511954
rect 414570 511718 414806 511954
rect 413930 511398 414166 511634
rect 414250 511398 414486 511634
rect 414570 511398 414806 511634
rect 433930 511718 434166 511954
rect 434250 511718 434486 511954
rect 434570 511718 434806 511954
rect 433930 511398 434166 511634
rect 434250 511398 434486 511634
rect 434570 511398 434806 511634
rect 453930 511718 454166 511954
rect 454250 511718 454486 511954
rect 454570 511718 454806 511954
rect 453930 511398 454166 511634
rect 454250 511398 454486 511634
rect 454570 511398 454806 511634
rect 473930 511718 474166 511954
rect 474250 511718 474486 511954
rect 474570 511718 474806 511954
rect 473930 511398 474166 511634
rect 474250 511398 474486 511634
rect 474570 511398 474806 511634
rect 303930 507218 304166 507454
rect 304250 507218 304486 507454
rect 304570 507218 304806 507454
rect 303930 506898 304166 507134
rect 304250 506898 304486 507134
rect 304570 506898 304806 507134
rect 323930 507218 324166 507454
rect 324250 507218 324486 507454
rect 324570 507218 324806 507454
rect 323930 506898 324166 507134
rect 324250 506898 324486 507134
rect 324570 506898 324806 507134
rect 343930 507218 344166 507454
rect 344250 507218 344486 507454
rect 344570 507218 344806 507454
rect 343930 506898 344166 507134
rect 344250 506898 344486 507134
rect 344570 506898 344806 507134
rect 363930 507218 364166 507454
rect 364250 507218 364486 507454
rect 364570 507218 364806 507454
rect 363930 506898 364166 507134
rect 364250 506898 364486 507134
rect 364570 506898 364806 507134
rect 383930 507218 384166 507454
rect 384250 507218 384486 507454
rect 384570 507218 384806 507454
rect 383930 506898 384166 507134
rect 384250 506898 384486 507134
rect 384570 506898 384806 507134
rect 403930 507218 404166 507454
rect 404250 507218 404486 507454
rect 404570 507218 404806 507454
rect 403930 506898 404166 507134
rect 404250 506898 404486 507134
rect 404570 506898 404806 507134
rect 423930 507218 424166 507454
rect 424250 507218 424486 507454
rect 424570 507218 424806 507454
rect 423930 506898 424166 507134
rect 424250 506898 424486 507134
rect 424570 506898 424806 507134
rect 443930 507218 444166 507454
rect 444250 507218 444486 507454
rect 444570 507218 444806 507454
rect 443930 506898 444166 507134
rect 444250 506898 444486 507134
rect 444570 506898 444806 507134
rect 463930 507218 464166 507454
rect 464250 507218 464486 507454
rect 464570 507218 464806 507454
rect 463930 506898 464166 507134
rect 464250 506898 464486 507134
rect 464570 506898 464806 507134
rect 313930 475718 314166 475954
rect 314250 475718 314486 475954
rect 314570 475718 314806 475954
rect 313930 475398 314166 475634
rect 314250 475398 314486 475634
rect 314570 475398 314806 475634
rect 333930 475718 334166 475954
rect 334250 475718 334486 475954
rect 334570 475718 334806 475954
rect 333930 475398 334166 475634
rect 334250 475398 334486 475634
rect 334570 475398 334806 475634
rect 353930 475718 354166 475954
rect 354250 475718 354486 475954
rect 354570 475718 354806 475954
rect 353930 475398 354166 475634
rect 354250 475398 354486 475634
rect 354570 475398 354806 475634
rect 373930 475718 374166 475954
rect 374250 475718 374486 475954
rect 374570 475718 374806 475954
rect 373930 475398 374166 475634
rect 374250 475398 374486 475634
rect 374570 475398 374806 475634
rect 393930 475718 394166 475954
rect 394250 475718 394486 475954
rect 394570 475718 394806 475954
rect 393930 475398 394166 475634
rect 394250 475398 394486 475634
rect 394570 475398 394806 475634
rect 413930 475718 414166 475954
rect 414250 475718 414486 475954
rect 414570 475718 414806 475954
rect 413930 475398 414166 475634
rect 414250 475398 414486 475634
rect 414570 475398 414806 475634
rect 433930 475718 434166 475954
rect 434250 475718 434486 475954
rect 434570 475718 434806 475954
rect 433930 475398 434166 475634
rect 434250 475398 434486 475634
rect 434570 475398 434806 475634
rect 453930 475718 454166 475954
rect 454250 475718 454486 475954
rect 454570 475718 454806 475954
rect 453930 475398 454166 475634
rect 454250 475398 454486 475634
rect 454570 475398 454806 475634
rect 473930 475718 474166 475954
rect 474250 475718 474486 475954
rect 474570 475718 474806 475954
rect 473930 475398 474166 475634
rect 474250 475398 474486 475634
rect 474570 475398 474806 475634
rect 303930 471218 304166 471454
rect 304250 471218 304486 471454
rect 304570 471218 304806 471454
rect 303930 470898 304166 471134
rect 304250 470898 304486 471134
rect 304570 470898 304806 471134
rect 323930 471218 324166 471454
rect 324250 471218 324486 471454
rect 324570 471218 324806 471454
rect 323930 470898 324166 471134
rect 324250 470898 324486 471134
rect 324570 470898 324806 471134
rect 343930 471218 344166 471454
rect 344250 471218 344486 471454
rect 344570 471218 344806 471454
rect 343930 470898 344166 471134
rect 344250 470898 344486 471134
rect 344570 470898 344806 471134
rect 363930 471218 364166 471454
rect 364250 471218 364486 471454
rect 364570 471218 364806 471454
rect 363930 470898 364166 471134
rect 364250 470898 364486 471134
rect 364570 470898 364806 471134
rect 383930 471218 384166 471454
rect 384250 471218 384486 471454
rect 384570 471218 384806 471454
rect 383930 470898 384166 471134
rect 384250 470898 384486 471134
rect 384570 470898 384806 471134
rect 403930 471218 404166 471454
rect 404250 471218 404486 471454
rect 404570 471218 404806 471454
rect 403930 470898 404166 471134
rect 404250 470898 404486 471134
rect 404570 470898 404806 471134
rect 423930 471218 424166 471454
rect 424250 471218 424486 471454
rect 424570 471218 424806 471454
rect 423930 470898 424166 471134
rect 424250 470898 424486 471134
rect 424570 470898 424806 471134
rect 443930 471218 444166 471454
rect 444250 471218 444486 471454
rect 444570 471218 444806 471454
rect 443930 470898 444166 471134
rect 444250 470898 444486 471134
rect 444570 470898 444806 471134
rect 463930 471218 464166 471454
rect 464250 471218 464486 471454
rect 464570 471218 464806 471454
rect 463930 470898 464166 471134
rect 464250 470898 464486 471134
rect 464570 470898 464806 471134
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 313930 439718 314166 439954
rect 314250 439718 314486 439954
rect 314570 439718 314806 439954
rect 313930 439398 314166 439634
rect 314250 439398 314486 439634
rect 314570 439398 314806 439634
rect 333930 439718 334166 439954
rect 334250 439718 334486 439954
rect 334570 439718 334806 439954
rect 333930 439398 334166 439634
rect 334250 439398 334486 439634
rect 334570 439398 334806 439634
rect 353930 439718 354166 439954
rect 354250 439718 354486 439954
rect 354570 439718 354806 439954
rect 353930 439398 354166 439634
rect 354250 439398 354486 439634
rect 354570 439398 354806 439634
rect 373930 439718 374166 439954
rect 374250 439718 374486 439954
rect 374570 439718 374806 439954
rect 373930 439398 374166 439634
rect 374250 439398 374486 439634
rect 374570 439398 374806 439634
rect 393930 439718 394166 439954
rect 394250 439718 394486 439954
rect 394570 439718 394806 439954
rect 393930 439398 394166 439634
rect 394250 439398 394486 439634
rect 394570 439398 394806 439634
rect 413930 439718 414166 439954
rect 414250 439718 414486 439954
rect 414570 439718 414806 439954
rect 413930 439398 414166 439634
rect 414250 439398 414486 439634
rect 414570 439398 414806 439634
rect 433930 439718 434166 439954
rect 434250 439718 434486 439954
rect 434570 439718 434806 439954
rect 433930 439398 434166 439634
rect 434250 439398 434486 439634
rect 434570 439398 434806 439634
rect 453930 439718 454166 439954
rect 454250 439718 454486 439954
rect 454570 439718 454806 439954
rect 453930 439398 454166 439634
rect 454250 439398 454486 439634
rect 454570 439398 454806 439634
rect 473930 439718 474166 439954
rect 474250 439718 474486 439954
rect 474570 439718 474806 439954
rect 473930 439398 474166 439634
rect 474250 439398 474486 439634
rect 474570 439398 474806 439634
rect 303930 435218 304166 435454
rect 304250 435218 304486 435454
rect 304570 435218 304806 435454
rect 303930 434898 304166 435134
rect 304250 434898 304486 435134
rect 304570 434898 304806 435134
rect 323930 435218 324166 435454
rect 324250 435218 324486 435454
rect 324570 435218 324806 435454
rect 323930 434898 324166 435134
rect 324250 434898 324486 435134
rect 324570 434898 324806 435134
rect 343930 435218 344166 435454
rect 344250 435218 344486 435454
rect 344570 435218 344806 435454
rect 343930 434898 344166 435134
rect 344250 434898 344486 435134
rect 344570 434898 344806 435134
rect 363930 435218 364166 435454
rect 364250 435218 364486 435454
rect 364570 435218 364806 435454
rect 363930 434898 364166 435134
rect 364250 434898 364486 435134
rect 364570 434898 364806 435134
rect 383930 435218 384166 435454
rect 384250 435218 384486 435454
rect 384570 435218 384806 435454
rect 383930 434898 384166 435134
rect 384250 434898 384486 435134
rect 384570 434898 384806 435134
rect 403930 435218 404166 435454
rect 404250 435218 404486 435454
rect 404570 435218 404806 435454
rect 403930 434898 404166 435134
rect 404250 434898 404486 435134
rect 404570 434898 404806 435134
rect 423930 435218 424166 435454
rect 424250 435218 424486 435454
rect 424570 435218 424806 435454
rect 423930 434898 424166 435134
rect 424250 434898 424486 435134
rect 424570 434898 424806 435134
rect 443930 435218 444166 435454
rect 444250 435218 444486 435454
rect 444570 435218 444806 435454
rect 443930 434898 444166 435134
rect 444250 434898 444486 435134
rect 444570 434898 444806 435134
rect 463930 435218 464166 435454
rect 464250 435218 464486 435454
rect 464570 435218 464806 435454
rect 463930 434898 464166 435134
rect 464250 434898 464486 435134
rect 464570 434898 464806 435134
rect 313930 403718 314166 403954
rect 314250 403718 314486 403954
rect 314570 403718 314806 403954
rect 313930 403398 314166 403634
rect 314250 403398 314486 403634
rect 314570 403398 314806 403634
rect 333930 403718 334166 403954
rect 334250 403718 334486 403954
rect 334570 403718 334806 403954
rect 333930 403398 334166 403634
rect 334250 403398 334486 403634
rect 334570 403398 334806 403634
rect 353930 403718 354166 403954
rect 354250 403718 354486 403954
rect 354570 403718 354806 403954
rect 353930 403398 354166 403634
rect 354250 403398 354486 403634
rect 354570 403398 354806 403634
rect 373930 403718 374166 403954
rect 374250 403718 374486 403954
rect 374570 403718 374806 403954
rect 373930 403398 374166 403634
rect 374250 403398 374486 403634
rect 374570 403398 374806 403634
rect 393930 403718 394166 403954
rect 394250 403718 394486 403954
rect 394570 403718 394806 403954
rect 393930 403398 394166 403634
rect 394250 403398 394486 403634
rect 394570 403398 394806 403634
rect 413930 403718 414166 403954
rect 414250 403718 414486 403954
rect 414570 403718 414806 403954
rect 413930 403398 414166 403634
rect 414250 403398 414486 403634
rect 414570 403398 414806 403634
rect 433930 403718 434166 403954
rect 434250 403718 434486 403954
rect 434570 403718 434806 403954
rect 433930 403398 434166 403634
rect 434250 403398 434486 403634
rect 434570 403398 434806 403634
rect 453930 403718 454166 403954
rect 454250 403718 454486 403954
rect 454570 403718 454806 403954
rect 453930 403398 454166 403634
rect 454250 403398 454486 403634
rect 454570 403398 454806 403634
rect 473930 403718 474166 403954
rect 474250 403718 474486 403954
rect 474570 403718 474806 403954
rect 473930 403398 474166 403634
rect 474250 403398 474486 403634
rect 474570 403398 474806 403634
rect 303930 399218 304166 399454
rect 304250 399218 304486 399454
rect 304570 399218 304806 399454
rect 303930 398898 304166 399134
rect 304250 398898 304486 399134
rect 304570 398898 304806 399134
rect 323930 399218 324166 399454
rect 324250 399218 324486 399454
rect 324570 399218 324806 399454
rect 323930 398898 324166 399134
rect 324250 398898 324486 399134
rect 324570 398898 324806 399134
rect 343930 399218 344166 399454
rect 344250 399218 344486 399454
rect 344570 399218 344806 399454
rect 343930 398898 344166 399134
rect 344250 398898 344486 399134
rect 344570 398898 344806 399134
rect 363930 399218 364166 399454
rect 364250 399218 364486 399454
rect 364570 399218 364806 399454
rect 363930 398898 364166 399134
rect 364250 398898 364486 399134
rect 364570 398898 364806 399134
rect 383930 399218 384166 399454
rect 384250 399218 384486 399454
rect 384570 399218 384806 399454
rect 383930 398898 384166 399134
rect 384250 398898 384486 399134
rect 384570 398898 384806 399134
rect 403930 399218 404166 399454
rect 404250 399218 404486 399454
rect 404570 399218 404806 399454
rect 403930 398898 404166 399134
rect 404250 398898 404486 399134
rect 404570 398898 404806 399134
rect 423930 399218 424166 399454
rect 424250 399218 424486 399454
rect 424570 399218 424806 399454
rect 423930 398898 424166 399134
rect 424250 398898 424486 399134
rect 424570 398898 424806 399134
rect 443930 399218 444166 399454
rect 444250 399218 444486 399454
rect 444570 399218 444806 399454
rect 443930 398898 444166 399134
rect 444250 398898 444486 399134
rect 444570 398898 444806 399134
rect 463930 399218 464166 399454
rect 464250 399218 464486 399454
rect 464570 399218 464806 399454
rect 463930 398898 464166 399134
rect 464250 398898 464486 399134
rect 464570 398898 464806 399134
rect 313930 367718 314166 367954
rect 314250 367718 314486 367954
rect 314570 367718 314806 367954
rect 313930 367398 314166 367634
rect 314250 367398 314486 367634
rect 314570 367398 314806 367634
rect 333930 367718 334166 367954
rect 334250 367718 334486 367954
rect 334570 367718 334806 367954
rect 333930 367398 334166 367634
rect 334250 367398 334486 367634
rect 334570 367398 334806 367634
rect 353930 367718 354166 367954
rect 354250 367718 354486 367954
rect 354570 367718 354806 367954
rect 353930 367398 354166 367634
rect 354250 367398 354486 367634
rect 354570 367398 354806 367634
rect 373930 367718 374166 367954
rect 374250 367718 374486 367954
rect 374570 367718 374806 367954
rect 373930 367398 374166 367634
rect 374250 367398 374486 367634
rect 374570 367398 374806 367634
rect 393930 367718 394166 367954
rect 394250 367718 394486 367954
rect 394570 367718 394806 367954
rect 393930 367398 394166 367634
rect 394250 367398 394486 367634
rect 394570 367398 394806 367634
rect 413930 367718 414166 367954
rect 414250 367718 414486 367954
rect 414570 367718 414806 367954
rect 413930 367398 414166 367634
rect 414250 367398 414486 367634
rect 414570 367398 414806 367634
rect 433930 367718 434166 367954
rect 434250 367718 434486 367954
rect 434570 367718 434806 367954
rect 433930 367398 434166 367634
rect 434250 367398 434486 367634
rect 434570 367398 434806 367634
rect 453930 367718 454166 367954
rect 454250 367718 454486 367954
rect 454570 367718 454806 367954
rect 453930 367398 454166 367634
rect 454250 367398 454486 367634
rect 454570 367398 454806 367634
rect 473930 367718 474166 367954
rect 474250 367718 474486 367954
rect 474570 367718 474806 367954
rect 473930 367398 474166 367634
rect 474250 367398 474486 367634
rect 474570 367398 474806 367634
rect 303930 363218 304166 363454
rect 304250 363218 304486 363454
rect 304570 363218 304806 363454
rect 303930 362898 304166 363134
rect 304250 362898 304486 363134
rect 304570 362898 304806 363134
rect 323930 363218 324166 363454
rect 324250 363218 324486 363454
rect 324570 363218 324806 363454
rect 323930 362898 324166 363134
rect 324250 362898 324486 363134
rect 324570 362898 324806 363134
rect 343930 363218 344166 363454
rect 344250 363218 344486 363454
rect 344570 363218 344806 363454
rect 343930 362898 344166 363134
rect 344250 362898 344486 363134
rect 344570 362898 344806 363134
rect 363930 363218 364166 363454
rect 364250 363218 364486 363454
rect 364570 363218 364806 363454
rect 363930 362898 364166 363134
rect 364250 362898 364486 363134
rect 364570 362898 364806 363134
rect 383930 363218 384166 363454
rect 384250 363218 384486 363454
rect 384570 363218 384806 363454
rect 383930 362898 384166 363134
rect 384250 362898 384486 363134
rect 384570 362898 384806 363134
rect 403930 363218 404166 363454
rect 404250 363218 404486 363454
rect 404570 363218 404806 363454
rect 403930 362898 404166 363134
rect 404250 362898 404486 363134
rect 404570 362898 404806 363134
rect 423930 363218 424166 363454
rect 424250 363218 424486 363454
rect 424570 363218 424806 363454
rect 423930 362898 424166 363134
rect 424250 362898 424486 363134
rect 424570 362898 424806 363134
rect 443930 363218 444166 363454
rect 444250 363218 444486 363454
rect 444570 363218 444806 363454
rect 443930 362898 444166 363134
rect 444250 362898 444486 363134
rect 444570 362898 444806 363134
rect 463930 363218 464166 363454
rect 464250 363218 464486 363454
rect 464570 363218 464806 363454
rect 463930 362898 464166 363134
rect 464250 362898 464486 363134
rect 464570 362898 464806 363134
rect 313930 295718 314166 295954
rect 314250 295718 314486 295954
rect 314570 295718 314806 295954
rect 313930 295398 314166 295634
rect 314250 295398 314486 295634
rect 314570 295398 314806 295634
rect 333930 295718 334166 295954
rect 334250 295718 334486 295954
rect 334570 295718 334806 295954
rect 333930 295398 334166 295634
rect 334250 295398 334486 295634
rect 334570 295398 334806 295634
rect 353930 295718 354166 295954
rect 354250 295718 354486 295954
rect 354570 295718 354806 295954
rect 353930 295398 354166 295634
rect 354250 295398 354486 295634
rect 354570 295398 354806 295634
rect 373930 295718 374166 295954
rect 374250 295718 374486 295954
rect 374570 295718 374806 295954
rect 373930 295398 374166 295634
rect 374250 295398 374486 295634
rect 374570 295398 374806 295634
rect 393930 295718 394166 295954
rect 394250 295718 394486 295954
rect 394570 295718 394806 295954
rect 393930 295398 394166 295634
rect 394250 295398 394486 295634
rect 394570 295398 394806 295634
rect 413930 295718 414166 295954
rect 414250 295718 414486 295954
rect 414570 295718 414806 295954
rect 413930 295398 414166 295634
rect 414250 295398 414486 295634
rect 414570 295398 414806 295634
rect 433930 295718 434166 295954
rect 434250 295718 434486 295954
rect 434570 295718 434806 295954
rect 433930 295398 434166 295634
rect 434250 295398 434486 295634
rect 434570 295398 434806 295634
rect 453930 295718 454166 295954
rect 454250 295718 454486 295954
rect 454570 295718 454806 295954
rect 453930 295398 454166 295634
rect 454250 295398 454486 295634
rect 454570 295398 454806 295634
rect 473930 295718 474166 295954
rect 474250 295718 474486 295954
rect 474570 295718 474806 295954
rect 473930 295398 474166 295634
rect 474250 295398 474486 295634
rect 474570 295398 474806 295634
rect 303930 291218 304166 291454
rect 304250 291218 304486 291454
rect 304570 291218 304806 291454
rect 303930 290898 304166 291134
rect 304250 290898 304486 291134
rect 304570 290898 304806 291134
rect 323930 291218 324166 291454
rect 324250 291218 324486 291454
rect 324570 291218 324806 291454
rect 323930 290898 324166 291134
rect 324250 290898 324486 291134
rect 324570 290898 324806 291134
rect 343930 291218 344166 291454
rect 344250 291218 344486 291454
rect 344570 291218 344806 291454
rect 343930 290898 344166 291134
rect 344250 290898 344486 291134
rect 344570 290898 344806 291134
rect 363930 291218 364166 291454
rect 364250 291218 364486 291454
rect 364570 291218 364806 291454
rect 363930 290898 364166 291134
rect 364250 290898 364486 291134
rect 364570 290898 364806 291134
rect 383930 291218 384166 291454
rect 384250 291218 384486 291454
rect 384570 291218 384806 291454
rect 383930 290898 384166 291134
rect 384250 290898 384486 291134
rect 384570 290898 384806 291134
rect 403930 291218 404166 291454
rect 404250 291218 404486 291454
rect 404570 291218 404806 291454
rect 403930 290898 404166 291134
rect 404250 290898 404486 291134
rect 404570 290898 404806 291134
rect 423930 291218 424166 291454
rect 424250 291218 424486 291454
rect 424570 291218 424806 291454
rect 423930 290898 424166 291134
rect 424250 290898 424486 291134
rect 424570 290898 424806 291134
rect 443930 291218 444166 291454
rect 444250 291218 444486 291454
rect 444570 291218 444806 291454
rect 443930 290898 444166 291134
rect 444250 290898 444486 291134
rect 444570 290898 444806 291134
rect 463930 291218 464166 291454
rect 464250 291218 464486 291454
rect 464570 291218 464806 291454
rect 463930 290898 464166 291134
rect 464250 290898 464486 291134
rect 464570 290898 464806 291134
rect 313930 259718 314166 259954
rect 314250 259718 314486 259954
rect 314570 259718 314806 259954
rect 313930 259398 314166 259634
rect 314250 259398 314486 259634
rect 314570 259398 314806 259634
rect 333930 259718 334166 259954
rect 334250 259718 334486 259954
rect 334570 259718 334806 259954
rect 333930 259398 334166 259634
rect 334250 259398 334486 259634
rect 334570 259398 334806 259634
rect 353930 259718 354166 259954
rect 354250 259718 354486 259954
rect 354570 259718 354806 259954
rect 353930 259398 354166 259634
rect 354250 259398 354486 259634
rect 354570 259398 354806 259634
rect 373930 259718 374166 259954
rect 374250 259718 374486 259954
rect 374570 259718 374806 259954
rect 373930 259398 374166 259634
rect 374250 259398 374486 259634
rect 374570 259398 374806 259634
rect 393930 259718 394166 259954
rect 394250 259718 394486 259954
rect 394570 259718 394806 259954
rect 393930 259398 394166 259634
rect 394250 259398 394486 259634
rect 394570 259398 394806 259634
rect 413930 259718 414166 259954
rect 414250 259718 414486 259954
rect 414570 259718 414806 259954
rect 413930 259398 414166 259634
rect 414250 259398 414486 259634
rect 414570 259398 414806 259634
rect 433930 259718 434166 259954
rect 434250 259718 434486 259954
rect 434570 259718 434806 259954
rect 433930 259398 434166 259634
rect 434250 259398 434486 259634
rect 434570 259398 434806 259634
rect 453930 259718 454166 259954
rect 454250 259718 454486 259954
rect 454570 259718 454806 259954
rect 453930 259398 454166 259634
rect 454250 259398 454486 259634
rect 454570 259398 454806 259634
rect 473930 259718 474166 259954
rect 474250 259718 474486 259954
rect 474570 259718 474806 259954
rect 473930 259398 474166 259634
rect 474250 259398 474486 259634
rect 474570 259398 474806 259634
rect 303930 255218 304166 255454
rect 304250 255218 304486 255454
rect 304570 255218 304806 255454
rect 303930 254898 304166 255134
rect 304250 254898 304486 255134
rect 304570 254898 304806 255134
rect 323930 255218 324166 255454
rect 324250 255218 324486 255454
rect 324570 255218 324806 255454
rect 323930 254898 324166 255134
rect 324250 254898 324486 255134
rect 324570 254898 324806 255134
rect 343930 255218 344166 255454
rect 344250 255218 344486 255454
rect 344570 255218 344806 255454
rect 343930 254898 344166 255134
rect 344250 254898 344486 255134
rect 344570 254898 344806 255134
rect 363930 255218 364166 255454
rect 364250 255218 364486 255454
rect 364570 255218 364806 255454
rect 363930 254898 364166 255134
rect 364250 254898 364486 255134
rect 364570 254898 364806 255134
rect 383930 255218 384166 255454
rect 384250 255218 384486 255454
rect 384570 255218 384806 255454
rect 383930 254898 384166 255134
rect 384250 254898 384486 255134
rect 384570 254898 384806 255134
rect 403930 255218 404166 255454
rect 404250 255218 404486 255454
rect 404570 255218 404806 255454
rect 403930 254898 404166 255134
rect 404250 254898 404486 255134
rect 404570 254898 404806 255134
rect 423930 255218 424166 255454
rect 424250 255218 424486 255454
rect 424570 255218 424806 255454
rect 423930 254898 424166 255134
rect 424250 254898 424486 255134
rect 424570 254898 424806 255134
rect 443930 255218 444166 255454
rect 444250 255218 444486 255454
rect 444570 255218 444806 255454
rect 443930 254898 444166 255134
rect 444250 254898 444486 255134
rect 444570 254898 444806 255134
rect 463930 255218 464166 255454
rect 464250 255218 464486 255454
rect 464570 255218 464806 255454
rect 463930 254898 464166 255134
rect 464250 254898 464486 255134
rect 464570 254898 464806 255134
rect 313930 223718 314166 223954
rect 314250 223718 314486 223954
rect 314570 223718 314806 223954
rect 313930 223398 314166 223634
rect 314250 223398 314486 223634
rect 314570 223398 314806 223634
rect 333930 223718 334166 223954
rect 334250 223718 334486 223954
rect 334570 223718 334806 223954
rect 333930 223398 334166 223634
rect 334250 223398 334486 223634
rect 334570 223398 334806 223634
rect 353930 223718 354166 223954
rect 354250 223718 354486 223954
rect 354570 223718 354806 223954
rect 353930 223398 354166 223634
rect 354250 223398 354486 223634
rect 354570 223398 354806 223634
rect 373930 223718 374166 223954
rect 374250 223718 374486 223954
rect 374570 223718 374806 223954
rect 373930 223398 374166 223634
rect 374250 223398 374486 223634
rect 374570 223398 374806 223634
rect 393930 223718 394166 223954
rect 394250 223718 394486 223954
rect 394570 223718 394806 223954
rect 393930 223398 394166 223634
rect 394250 223398 394486 223634
rect 394570 223398 394806 223634
rect 413930 223718 414166 223954
rect 414250 223718 414486 223954
rect 414570 223718 414806 223954
rect 413930 223398 414166 223634
rect 414250 223398 414486 223634
rect 414570 223398 414806 223634
rect 433930 223718 434166 223954
rect 434250 223718 434486 223954
rect 434570 223718 434806 223954
rect 433930 223398 434166 223634
rect 434250 223398 434486 223634
rect 434570 223398 434806 223634
rect 453930 223718 454166 223954
rect 454250 223718 454486 223954
rect 454570 223718 454806 223954
rect 453930 223398 454166 223634
rect 454250 223398 454486 223634
rect 454570 223398 454806 223634
rect 473930 223718 474166 223954
rect 474250 223718 474486 223954
rect 474570 223718 474806 223954
rect 473930 223398 474166 223634
rect 474250 223398 474486 223634
rect 474570 223398 474806 223634
rect 303930 219218 304166 219454
rect 304250 219218 304486 219454
rect 304570 219218 304806 219454
rect 303930 218898 304166 219134
rect 304250 218898 304486 219134
rect 304570 218898 304806 219134
rect 323930 219218 324166 219454
rect 324250 219218 324486 219454
rect 324570 219218 324806 219454
rect 323930 218898 324166 219134
rect 324250 218898 324486 219134
rect 324570 218898 324806 219134
rect 343930 219218 344166 219454
rect 344250 219218 344486 219454
rect 344570 219218 344806 219454
rect 343930 218898 344166 219134
rect 344250 218898 344486 219134
rect 344570 218898 344806 219134
rect 363930 219218 364166 219454
rect 364250 219218 364486 219454
rect 364570 219218 364806 219454
rect 363930 218898 364166 219134
rect 364250 218898 364486 219134
rect 364570 218898 364806 219134
rect 383930 219218 384166 219454
rect 384250 219218 384486 219454
rect 384570 219218 384806 219454
rect 383930 218898 384166 219134
rect 384250 218898 384486 219134
rect 384570 218898 384806 219134
rect 403930 219218 404166 219454
rect 404250 219218 404486 219454
rect 404570 219218 404806 219454
rect 403930 218898 404166 219134
rect 404250 218898 404486 219134
rect 404570 218898 404806 219134
rect 423930 219218 424166 219454
rect 424250 219218 424486 219454
rect 424570 219218 424806 219454
rect 423930 218898 424166 219134
rect 424250 218898 424486 219134
rect 424570 218898 424806 219134
rect 443930 219218 444166 219454
rect 444250 219218 444486 219454
rect 444570 219218 444806 219454
rect 443930 218898 444166 219134
rect 444250 218898 444486 219134
rect 444570 218898 444806 219134
rect 463930 219218 464166 219454
rect 464250 219218 464486 219454
rect 464570 219218 464806 219454
rect 463930 218898 464166 219134
rect 464250 218898 464486 219134
rect 464570 218898 464806 219134
rect 303930 183218 304166 183454
rect 304250 183218 304486 183454
rect 304570 183218 304806 183454
rect 303930 182898 304166 183134
rect 304250 182898 304486 183134
rect 304570 182898 304806 183134
rect 323930 183218 324166 183454
rect 324250 183218 324486 183454
rect 324570 183218 324806 183454
rect 323930 182898 324166 183134
rect 324250 182898 324486 183134
rect 324570 182898 324806 183134
rect 343930 183218 344166 183454
rect 344250 183218 344486 183454
rect 344570 183218 344806 183454
rect 343930 182898 344166 183134
rect 344250 182898 344486 183134
rect 344570 182898 344806 183134
rect 363930 183218 364166 183454
rect 364250 183218 364486 183454
rect 364570 183218 364806 183454
rect 363930 182898 364166 183134
rect 364250 182898 364486 183134
rect 364570 182898 364806 183134
rect 383930 183218 384166 183454
rect 384250 183218 384486 183454
rect 384570 183218 384806 183454
rect 383930 182898 384166 183134
rect 384250 182898 384486 183134
rect 384570 182898 384806 183134
rect 403930 183218 404166 183454
rect 404250 183218 404486 183454
rect 404570 183218 404806 183454
rect 403930 182898 404166 183134
rect 404250 182898 404486 183134
rect 404570 182898 404806 183134
rect 423930 183218 424166 183454
rect 424250 183218 424486 183454
rect 424570 183218 424806 183454
rect 423930 182898 424166 183134
rect 424250 182898 424486 183134
rect 424570 182898 424806 183134
rect 443930 183218 444166 183454
rect 444250 183218 444486 183454
rect 444570 183218 444806 183454
rect 443930 182898 444166 183134
rect 444250 182898 444486 183134
rect 444570 182898 444806 183134
rect 463930 183218 464166 183454
rect 464250 183218 464486 183454
rect 464570 183218 464806 183454
rect 463930 182898 464166 183134
rect 464250 182898 464486 183134
rect 464570 182898 464806 183134
rect 313930 151718 314166 151954
rect 314250 151718 314486 151954
rect 314570 151718 314806 151954
rect 313930 151398 314166 151634
rect 314250 151398 314486 151634
rect 314570 151398 314806 151634
rect 333930 151718 334166 151954
rect 334250 151718 334486 151954
rect 334570 151718 334806 151954
rect 333930 151398 334166 151634
rect 334250 151398 334486 151634
rect 334570 151398 334806 151634
rect 353930 151718 354166 151954
rect 354250 151718 354486 151954
rect 354570 151718 354806 151954
rect 353930 151398 354166 151634
rect 354250 151398 354486 151634
rect 354570 151398 354806 151634
rect 373930 151718 374166 151954
rect 374250 151718 374486 151954
rect 374570 151718 374806 151954
rect 373930 151398 374166 151634
rect 374250 151398 374486 151634
rect 374570 151398 374806 151634
rect 393930 151718 394166 151954
rect 394250 151718 394486 151954
rect 394570 151718 394806 151954
rect 393930 151398 394166 151634
rect 394250 151398 394486 151634
rect 394570 151398 394806 151634
rect 413930 151718 414166 151954
rect 414250 151718 414486 151954
rect 414570 151718 414806 151954
rect 413930 151398 414166 151634
rect 414250 151398 414486 151634
rect 414570 151398 414806 151634
rect 433930 151718 434166 151954
rect 434250 151718 434486 151954
rect 434570 151718 434806 151954
rect 433930 151398 434166 151634
rect 434250 151398 434486 151634
rect 434570 151398 434806 151634
rect 453930 151718 454166 151954
rect 454250 151718 454486 151954
rect 454570 151718 454806 151954
rect 453930 151398 454166 151634
rect 454250 151398 454486 151634
rect 454570 151398 454806 151634
rect 473930 151718 474166 151954
rect 474250 151718 474486 151954
rect 474570 151718 474806 151954
rect 473930 151398 474166 151634
rect 474250 151398 474486 151634
rect 474570 151398 474806 151634
rect 303930 147218 304166 147454
rect 304250 147218 304486 147454
rect 304570 147218 304806 147454
rect 303930 146898 304166 147134
rect 304250 146898 304486 147134
rect 304570 146898 304806 147134
rect 323930 147218 324166 147454
rect 324250 147218 324486 147454
rect 324570 147218 324806 147454
rect 323930 146898 324166 147134
rect 324250 146898 324486 147134
rect 324570 146898 324806 147134
rect 343930 147218 344166 147454
rect 344250 147218 344486 147454
rect 344570 147218 344806 147454
rect 343930 146898 344166 147134
rect 344250 146898 344486 147134
rect 344570 146898 344806 147134
rect 363930 147218 364166 147454
rect 364250 147218 364486 147454
rect 364570 147218 364806 147454
rect 363930 146898 364166 147134
rect 364250 146898 364486 147134
rect 364570 146898 364806 147134
rect 383930 147218 384166 147454
rect 384250 147218 384486 147454
rect 384570 147218 384806 147454
rect 383930 146898 384166 147134
rect 384250 146898 384486 147134
rect 384570 146898 384806 147134
rect 403930 147218 404166 147454
rect 404250 147218 404486 147454
rect 404570 147218 404806 147454
rect 403930 146898 404166 147134
rect 404250 146898 404486 147134
rect 404570 146898 404806 147134
rect 423930 147218 424166 147454
rect 424250 147218 424486 147454
rect 424570 147218 424806 147454
rect 423930 146898 424166 147134
rect 424250 146898 424486 147134
rect 424570 146898 424806 147134
rect 443930 147218 444166 147454
rect 444250 147218 444486 147454
rect 444570 147218 444806 147454
rect 443930 146898 444166 147134
rect 444250 146898 444486 147134
rect 444570 146898 444806 147134
rect 463930 147218 464166 147454
rect 464250 147218 464486 147454
rect 464570 147218 464806 147454
rect 463930 146898 464166 147134
rect 464250 146898 464486 147134
rect 464570 146898 464806 147134
rect 313930 115718 314166 115954
rect 314250 115718 314486 115954
rect 314570 115718 314806 115954
rect 313930 115398 314166 115634
rect 314250 115398 314486 115634
rect 314570 115398 314806 115634
rect 333930 115718 334166 115954
rect 334250 115718 334486 115954
rect 334570 115718 334806 115954
rect 333930 115398 334166 115634
rect 334250 115398 334486 115634
rect 334570 115398 334806 115634
rect 353930 115718 354166 115954
rect 354250 115718 354486 115954
rect 354570 115718 354806 115954
rect 353930 115398 354166 115634
rect 354250 115398 354486 115634
rect 354570 115398 354806 115634
rect 373930 115718 374166 115954
rect 374250 115718 374486 115954
rect 374570 115718 374806 115954
rect 373930 115398 374166 115634
rect 374250 115398 374486 115634
rect 374570 115398 374806 115634
rect 393930 115718 394166 115954
rect 394250 115718 394486 115954
rect 394570 115718 394806 115954
rect 393930 115398 394166 115634
rect 394250 115398 394486 115634
rect 394570 115398 394806 115634
rect 413930 115718 414166 115954
rect 414250 115718 414486 115954
rect 414570 115718 414806 115954
rect 413930 115398 414166 115634
rect 414250 115398 414486 115634
rect 414570 115398 414806 115634
rect 433930 115718 434166 115954
rect 434250 115718 434486 115954
rect 434570 115718 434806 115954
rect 433930 115398 434166 115634
rect 434250 115398 434486 115634
rect 434570 115398 434806 115634
rect 453930 115718 454166 115954
rect 454250 115718 454486 115954
rect 454570 115718 454806 115954
rect 453930 115398 454166 115634
rect 454250 115398 454486 115634
rect 454570 115398 454806 115634
rect 473930 115718 474166 115954
rect 474250 115718 474486 115954
rect 474570 115718 474806 115954
rect 473930 115398 474166 115634
rect 474250 115398 474486 115634
rect 474570 115398 474806 115634
rect 303930 111218 304166 111454
rect 304250 111218 304486 111454
rect 304570 111218 304806 111454
rect 303930 110898 304166 111134
rect 304250 110898 304486 111134
rect 304570 110898 304806 111134
rect 323930 111218 324166 111454
rect 324250 111218 324486 111454
rect 324570 111218 324806 111454
rect 323930 110898 324166 111134
rect 324250 110898 324486 111134
rect 324570 110898 324806 111134
rect 343930 111218 344166 111454
rect 344250 111218 344486 111454
rect 344570 111218 344806 111454
rect 343930 110898 344166 111134
rect 344250 110898 344486 111134
rect 344570 110898 344806 111134
rect 363930 111218 364166 111454
rect 364250 111218 364486 111454
rect 364570 111218 364806 111454
rect 363930 110898 364166 111134
rect 364250 110898 364486 111134
rect 364570 110898 364806 111134
rect 383930 111218 384166 111454
rect 384250 111218 384486 111454
rect 384570 111218 384806 111454
rect 383930 110898 384166 111134
rect 384250 110898 384486 111134
rect 384570 110898 384806 111134
rect 403930 111218 404166 111454
rect 404250 111218 404486 111454
rect 404570 111218 404806 111454
rect 403930 110898 404166 111134
rect 404250 110898 404486 111134
rect 404570 110898 404806 111134
rect 423930 111218 424166 111454
rect 424250 111218 424486 111454
rect 424570 111218 424806 111454
rect 423930 110898 424166 111134
rect 424250 110898 424486 111134
rect 424570 110898 424806 111134
rect 443930 111218 444166 111454
rect 444250 111218 444486 111454
rect 444570 111218 444806 111454
rect 443930 110898 444166 111134
rect 444250 110898 444486 111134
rect 444570 110898 444806 111134
rect 463930 111218 464166 111454
rect 464250 111218 464486 111454
rect 464570 111218 464806 111454
rect 463930 110898 464166 111134
rect 464250 110898 464486 111134
rect 464570 110898 464806 111134
rect 213930 43718 214166 43954
rect 214250 43718 214486 43954
rect 214570 43718 214806 43954
rect 213930 43398 214166 43634
rect 214250 43398 214486 43634
rect 214570 43398 214806 43634
rect 233930 43718 234166 43954
rect 234250 43718 234486 43954
rect 234570 43718 234806 43954
rect 233930 43398 234166 43634
rect 234250 43398 234486 43634
rect 234570 43398 234806 43634
rect 253930 43718 254166 43954
rect 254250 43718 254486 43954
rect 254570 43718 254806 43954
rect 253930 43398 254166 43634
rect 254250 43398 254486 43634
rect 254570 43398 254806 43634
rect 273930 43718 274166 43954
rect 274250 43718 274486 43954
rect 274570 43718 274806 43954
rect 273930 43398 274166 43634
rect 274250 43398 274486 43634
rect 274570 43398 274806 43634
rect 293930 43718 294166 43954
rect 294250 43718 294486 43954
rect 294570 43718 294806 43954
rect 293930 43398 294166 43634
rect 294250 43398 294486 43634
rect 294570 43398 294806 43634
rect 313930 43718 314166 43954
rect 314250 43718 314486 43954
rect 314570 43718 314806 43954
rect 313930 43398 314166 43634
rect 314250 43398 314486 43634
rect 314570 43398 314806 43634
rect 333930 43718 334166 43954
rect 334250 43718 334486 43954
rect 334570 43718 334806 43954
rect 333930 43398 334166 43634
rect 334250 43398 334486 43634
rect 334570 43398 334806 43634
rect 353930 43718 354166 43954
rect 354250 43718 354486 43954
rect 354570 43718 354806 43954
rect 353930 43398 354166 43634
rect 354250 43398 354486 43634
rect 354570 43398 354806 43634
rect 373930 43718 374166 43954
rect 374250 43718 374486 43954
rect 374570 43718 374806 43954
rect 373930 43398 374166 43634
rect 374250 43398 374486 43634
rect 374570 43398 374806 43634
rect 393930 43718 394166 43954
rect 394250 43718 394486 43954
rect 394570 43718 394806 43954
rect 393930 43398 394166 43634
rect 394250 43398 394486 43634
rect 394570 43398 394806 43634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 203930 39218 204166 39454
rect 204250 39218 204486 39454
rect 204570 39218 204806 39454
rect 203930 38898 204166 39134
rect 204250 38898 204486 39134
rect 204570 38898 204806 39134
rect 223930 39218 224166 39454
rect 224250 39218 224486 39454
rect 224570 39218 224806 39454
rect 223930 38898 224166 39134
rect 224250 38898 224486 39134
rect 224570 38898 224806 39134
rect 243930 39218 244166 39454
rect 244250 39218 244486 39454
rect 244570 39218 244806 39454
rect 243930 38898 244166 39134
rect 244250 38898 244486 39134
rect 244570 38898 244806 39134
rect 263930 39218 264166 39454
rect 264250 39218 264486 39454
rect 264570 39218 264806 39454
rect 263930 38898 264166 39134
rect 264250 38898 264486 39134
rect 264570 38898 264806 39134
rect 283930 39218 284166 39454
rect 284250 39218 284486 39454
rect 284570 39218 284806 39454
rect 283930 38898 284166 39134
rect 284250 38898 284486 39134
rect 284570 38898 284806 39134
rect 303930 39218 304166 39454
rect 304250 39218 304486 39454
rect 304570 39218 304806 39454
rect 303930 38898 304166 39134
rect 304250 38898 304486 39134
rect 304570 38898 304806 39134
rect 323930 39218 324166 39454
rect 324250 39218 324486 39454
rect 324570 39218 324806 39454
rect 323930 38898 324166 39134
rect 324250 38898 324486 39134
rect 324570 38898 324806 39134
rect 343930 39218 344166 39454
rect 344250 39218 344486 39454
rect 344570 39218 344806 39454
rect 343930 38898 344166 39134
rect 344250 38898 344486 39134
rect 344570 38898 344806 39134
rect 363930 39218 364166 39454
rect 364250 39218 364486 39454
rect 364570 39218 364806 39454
rect 363930 38898 364166 39134
rect 364250 38898 364486 39134
rect 364570 38898 364806 39134
rect 383930 39218 384166 39454
rect 384250 39218 384486 39454
rect 384570 39218 384806 39454
rect 383930 38898 384166 39134
rect 384250 38898 384486 39134
rect 384570 38898 384806 39134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 79610 43954
rect 79846 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 79610 43634
rect 79846 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 64250 39454
rect 64486 39218 94970 39454
rect 95206 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 64250 39134
rect 64486 38898 94970 39134
rect 95206 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use controller_core  controller_core_mod
timestamp 0
transform 1 0 200000 0 1 24000
box -800 -800 198812 30800
use driver_core  driver_core_0
timestamp 0
transform 1 0 20000 0 1 78000
box 1066 -800 178886 107760
use driver_core  driver_core_1
timestamp 0
transform 1 0 20000 0 1 206000
box 1066 -800 178886 107760
use driver_core  driver_core_2
timestamp 0
transform 1 0 20000 0 1 334000
box 1066 -800 178886 107760
use driver_core  driver_core_3
timestamp 0
transform 1 0 20000 0 1 462000
box 1066 -800 178886 107760
use driver_core  driver_core_4
timestamp 0
transform 1 0 20000 0 1 588000
box 1066 -800 178886 107760
use driver_core  driver_core_5
timestamp 0
transform 1 0 300000 0 1 588000
box 1066 -800 178886 107760
use driver_core  driver_core_6
timestamp 0
transform 1 0 300000 0 1 462000
box 1066 -800 178886 107760
use driver_core  driver_core_7
timestamp 0
transform 1 0 300000 0 1 334000
box 1066 -800 178886 107760
use driver_core  driver_core_8
timestamp 0
transform 1 0 300000 0 1 206000
box 1066 -800 178886 107760
use driver_core  driver_core_9
timestamp 0
transform 1 0 300000 0 1 78000
box 1066 -800 178886 107760
use spi_controller  spi_controller_mod
timestamp 0
transform 1 0 60000 0 1 24000
box 0 0 40000 37584
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 56000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 56000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 56000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 56000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 56000 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 56000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 56000 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 56000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 56000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 56000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 56000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 56000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 56000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 56000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 56000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 56000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 56000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 56000 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 56000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 700000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 700000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 700000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 700000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 700000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 56000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 56000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 700000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 700000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 700000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 700000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 700000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
