magic
tech sky130B
magscale 1 2
timestamp 1662518344
<< metal1 >>
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 72970 700992 72976 701004
rect 8168 700964 72976 700992
rect 8168 700952 8174 700964
rect 72970 700952 72976 700964
rect 73028 700952 73034 701004
rect 397454 700952 397460 701004
rect 397512 700992 397518 701004
rect 418154 700992 418160 701004
rect 397512 700964 418160 700992
rect 397512 700952 397518 700964
rect 418154 700952 418160 700964
rect 418212 700992 418218 701004
rect 462314 700992 462320 701004
rect 418212 700964 462320 700992
rect 418212 700952 418218 700964
rect 462314 700952 462320 700964
rect 462372 700952 462378 701004
rect 20622 700340 20628 700392
rect 20680 700380 20686 700392
rect 89162 700380 89168 700392
rect 20680 700352 89168 700380
rect 20680 700340 20686 700352
rect 89162 700340 89168 700352
rect 89220 700340 89226 700392
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 198734 700380 198740 700392
rect 137888 700352 198740 700380
rect 137888 700340 137894 700352
rect 198734 700340 198740 700352
rect 198792 700340 198798 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 199378 700312 199384 700324
rect 73028 700284 199384 700312
rect 73028 700272 73034 700284
rect 199378 700272 199384 700284
rect 199436 700272 199442 700324
rect 198734 699796 198740 699848
rect 198792 699836 198798 699848
rect 200022 699836 200028 699848
rect 198792 699808 200028 699836
rect 198792 699796 198798 699808
rect 200022 699796 200028 699808
rect 200080 699836 200086 699848
rect 202782 699836 202788 699848
rect 200080 699808 202788 699836
rect 200080 699796 200086 699808
rect 202782 699796 202788 699808
rect 202840 699796 202846 699848
rect 20714 699660 20720 699712
rect 20772 699700 20778 699712
rect 24302 699700 24308 699712
rect 20772 699672 24308 699700
rect 20772 699660 20778 699672
rect 24302 699660 24308 699672
rect 24360 699660 24366 699712
rect 527174 697552 527180 697604
rect 527232 697592 527238 697604
rect 527818 697592 527824 697604
rect 527232 697564 527824 697592
rect 527232 697552 527238 697564
rect 527818 697552 527824 697564
rect 527876 697592 527882 697604
rect 580166 697592 580172 697604
rect 527876 697564 580172 697592
rect 527876 697552 527882 697564
rect 580166 697552 580172 697564
rect 580224 697552 580230 697604
rect 300854 667156 300860 667208
rect 300912 667196 300918 667208
rect 412634 667196 412640 667208
rect 300912 667168 412640 667196
rect 300912 667156 300918 667168
rect 412634 667156 412640 667168
rect 412692 667156 412698 667208
rect 304534 586508 304540 586560
rect 304592 586548 304598 586560
rect 477494 586548 477500 586560
rect 304592 586520 477500 586548
rect 304592 586508 304598 586520
rect 477494 586508 477500 586520
rect 477552 586508 477558 586560
rect 22002 586440 22008 586492
rect 22060 586480 22066 586492
rect 153194 586480 153200 586492
rect 22060 586452 153200 586480
rect 22060 586440 22066 586452
rect 153194 586440 153200 586452
rect 153252 586440 153258 586492
rect 348418 586440 348424 586492
rect 348476 586480 348482 586492
rect 350902 586480 350908 586492
rect 348476 586452 350908 586480
rect 348476 586440 348482 586452
rect 350902 586440 350908 586452
rect 350960 586440 350966 586492
rect 68646 586372 68652 586424
rect 68704 586412 68710 586424
rect 71038 586412 71044 586424
rect 68704 586384 71044 586412
rect 68704 586372 68710 586384
rect 71038 586372 71044 586384
rect 71096 586372 71102 586424
rect 300762 586100 300768 586152
rect 300820 586140 300826 586152
rect 309686 586140 309692 586152
rect 300820 586112 309692 586140
rect 300820 586100 300826 586112
rect 309686 586100 309692 586112
rect 309744 586100 309750 586152
rect 410150 586100 410156 586152
rect 410208 586140 410214 586152
rect 418798 586140 418804 586152
rect 410208 586112 418804 586140
rect 410208 586100 410214 586112
rect 418798 586100 418804 586112
rect 418856 586100 418862 586152
rect 20346 586032 20352 586084
rect 20404 586072 20410 586084
rect 29362 586072 29368 586084
rect 20404 586044 29368 586072
rect 20404 586032 20410 586044
rect 29362 586032 29368 586044
rect 29420 586032 29426 586084
rect 130470 586032 130476 586084
rect 130528 586072 130534 586084
rect 139486 586072 139492 586084
rect 130528 586044 139492 586072
rect 130528 586032 130534 586044
rect 139486 586032 139492 586044
rect 139544 586032 139550 586084
rect 300578 586032 300584 586084
rect 300636 586072 300642 586084
rect 312262 586072 312268 586084
rect 300636 586044 312268 586072
rect 300636 586032 300642 586044
rect 312262 586032 312268 586044
rect 312320 586032 312326 586084
rect 407574 586032 407580 586084
rect 407632 586072 407638 586084
rect 419534 586072 419540 586084
rect 407632 586044 419540 586072
rect 407632 586032 407638 586044
rect 419534 586032 419540 586044
rect 419592 586032 419598 586084
rect 21358 585964 21364 586016
rect 21416 586004 21422 586016
rect 31938 586004 31944 586016
rect 21416 585976 31944 586004
rect 21416 585964 21422 585976
rect 31938 585964 31944 585976
rect 31996 585964 32002 586016
rect 127894 585964 127900 586016
rect 127952 586004 127958 586016
rect 138658 586004 138664 586016
rect 127952 585976 138664 586004
rect 127952 585964 127958 585976
rect 138658 585964 138664 585976
rect 138716 585964 138722 586016
rect 301222 585964 301228 586016
rect 301280 586004 301286 586016
rect 314838 586004 314844 586016
rect 301280 585976 314844 586004
rect 301280 585964 301286 585976
rect 314838 585964 314844 585976
rect 314896 585964 314902 586016
rect 404998 585964 405004 586016
rect 405056 586004 405062 586016
rect 405056 585976 415256 586004
rect 405056 585964 405062 585976
rect 19242 585896 19248 585948
rect 19300 585936 19306 585948
rect 34514 585936 34520 585948
rect 19300 585908 34520 585936
rect 19300 585896 19306 585908
rect 34514 585896 34520 585908
rect 34572 585896 34578 585948
rect 125318 585896 125324 585948
rect 125376 585936 125382 585948
rect 139394 585936 139400 585948
rect 125376 585908 139400 585936
rect 125376 585896 125382 585908
rect 139394 585896 139400 585908
rect 139452 585896 139458 585948
rect 299382 585896 299388 585948
rect 299440 585936 299446 585948
rect 317414 585936 317420 585948
rect 299440 585908 317420 585936
rect 299440 585896 299446 585908
rect 317414 585896 317420 585908
rect 317472 585896 317478 585948
rect 402422 585896 402428 585948
rect 402480 585936 402486 585948
rect 415118 585936 415124 585948
rect 402480 585908 415124 585936
rect 402480 585896 402486 585908
rect 415118 585896 415124 585908
rect 415176 585896 415182 585948
rect 415228 585936 415256 585976
rect 415302 585964 415308 586016
rect 415360 586004 415366 586016
rect 419626 586004 419632 586016
rect 415360 585976 419632 586004
rect 415360 585964 415366 585976
rect 419626 585964 419632 585976
rect 419684 585964 419690 586016
rect 418430 585936 418436 585948
rect 415228 585908 418436 585936
rect 418430 585896 418436 585908
rect 418488 585896 418494 585948
rect 17862 585828 17868 585880
rect 17920 585868 17926 585880
rect 37274 585868 37280 585880
rect 17920 585840 37280 585868
rect 17920 585828 17926 585840
rect 37274 585828 37280 585840
rect 37332 585828 37338 585880
rect 122742 585828 122748 585880
rect 122800 585868 122806 585880
rect 138566 585868 138572 585880
rect 122800 585840 138572 585868
rect 122800 585828 122806 585840
rect 138566 585828 138572 585840
rect 138624 585828 138630 585880
rect 299106 585828 299112 585880
rect 299164 585868 299170 585880
rect 319990 585868 319996 585880
rect 299164 585840 319996 585868
rect 299164 585828 299170 585840
rect 319990 585828 319996 585840
rect 320048 585828 320054 585880
rect 399846 585828 399852 585880
rect 399904 585868 399910 585880
rect 418338 585868 418344 585880
rect 399904 585840 418344 585868
rect 399904 585828 399910 585840
rect 418338 585828 418344 585840
rect 418396 585828 418402 585880
rect 19150 585760 19156 585812
rect 19208 585800 19214 585812
rect 39666 585800 39672 585812
rect 19208 585772 39672 585800
rect 19208 585760 19214 585772
rect 39666 585760 39672 585772
rect 39724 585760 39730 585812
rect 119982 585760 119988 585812
rect 120040 585800 120046 585812
rect 139854 585800 139860 585812
rect 120040 585772 139860 585800
rect 120040 585760 120046 585772
rect 139854 585760 139860 585772
rect 139912 585760 139918 585812
rect 301406 585760 301412 585812
rect 301464 585800 301470 585812
rect 332870 585800 332876 585812
rect 301464 585772 332876 585800
rect 301464 585760 301470 585772
rect 332870 585760 332876 585772
rect 332928 585760 332934 585812
rect 397270 585760 397276 585812
rect 397328 585800 397334 585812
rect 419810 585800 419816 585812
rect 397328 585772 419816 585800
rect 397328 585760 397334 585772
rect 419810 585760 419816 585772
rect 419868 585760 419874 585812
rect 415118 585692 415124 585744
rect 415176 585732 415182 585744
rect 419718 585732 419724 585744
rect 415176 585704 419724 585732
rect 415176 585692 415182 585704
rect 419718 585692 419724 585704
rect 419776 585692 419782 585744
rect 20530 585148 20536 585200
rect 20588 585188 20594 585200
rect 26786 585188 26792 585200
rect 20588 585160 26792 585188
rect 20588 585148 20594 585160
rect 26786 585148 26792 585160
rect 26844 585148 26850 585200
rect 135622 585148 135628 585200
rect 135680 585188 135686 585200
rect 138382 585188 138388 585200
rect 135680 585160 138388 585188
rect 135680 585148 135686 585160
rect 138382 585148 138388 585160
rect 138440 585148 138446 585200
rect 300394 585148 300400 585200
rect 300452 585188 300458 585200
rect 307110 585188 307116 585200
rect 300452 585160 307116 585188
rect 300452 585148 300458 585160
rect 307110 585148 307116 585160
rect 307168 585148 307174 585200
rect 299290 583380 299296 583432
rect 299348 583420 299354 583432
rect 322566 583420 322572 583432
rect 299348 583392 322572 583420
rect 299348 583380 299354 583392
rect 322566 583380 322572 583392
rect 322624 583380 322630 583432
rect 394694 583380 394700 583432
rect 394752 583420 394758 583432
rect 420914 583420 420920 583432
rect 394752 583392 420920 583420
rect 394752 583380 394758 583392
rect 420914 583380 420920 583392
rect 420972 583380 420978 583432
rect 17770 583312 17776 583364
rect 17828 583352 17834 583364
rect 42242 583352 42248 583364
rect 17828 583324 42248 583352
rect 17828 583312 17834 583324
rect 42242 583312 42248 583324
rect 42300 583312 42306 583364
rect 299198 583312 299204 583364
rect 299256 583352 299262 583364
rect 325142 583352 325148 583364
rect 299256 583324 325148 583352
rect 299256 583312 299262 583324
rect 325142 583312 325148 583324
rect 325200 583312 325206 583364
rect 392118 583312 392124 583364
rect 392176 583352 392182 583364
rect 422570 583352 422576 583364
rect 392176 583324 422576 583352
rect 392176 583312 392182 583324
rect 422570 583312 422576 583324
rect 422628 583312 422634 583364
rect 19058 583244 19064 583296
rect 19116 583284 19122 583296
rect 44818 583284 44824 583296
rect 19116 583256 44824 583284
rect 19116 583244 19122 583256
rect 44818 583244 44824 583256
rect 44876 583244 44882 583296
rect 115014 583244 115020 583296
rect 115072 583284 115078 583296
rect 140774 583284 140780 583296
rect 115072 583256 140780 583284
rect 115072 583244 115078 583256
rect 140774 583244 140780 583256
rect 140832 583244 140838 583296
rect 300486 583244 300492 583296
rect 300544 583284 300550 583296
rect 330294 583284 330300 583296
rect 300544 583256 330300 583284
rect 300544 583244 300550 583256
rect 330294 583244 330300 583256
rect 330352 583244 330358 583296
rect 389542 583244 389548 583296
rect 389600 583284 389606 583296
rect 421374 583284 421380 583296
rect 389600 583256 421380 583284
rect 389600 583244 389606 583256
rect 421374 583244 421380 583256
rect 421432 583244 421438 583296
rect 17678 583176 17684 583228
rect 17736 583216 17742 583228
rect 49970 583216 49976 583228
rect 17736 583188 49976 583216
rect 17736 583176 17742 583188
rect 49970 583176 49976 583188
rect 50028 583176 50034 583228
rect 109862 583176 109868 583228
rect 109920 583216 109926 583228
rect 138290 583216 138296 583228
rect 109920 583188 138296 583216
rect 109920 583176 109926 583188
rect 138290 583176 138296 583188
rect 138348 583176 138354 583228
rect 297910 583176 297916 583228
rect 297968 583216 297974 583228
rect 340598 583216 340604 583228
rect 297968 583188 340604 583216
rect 297968 583176 297974 583188
rect 340598 583176 340604 583188
rect 340656 583176 340662 583228
rect 386966 583176 386972 583228
rect 387024 583216 387030 583228
rect 421190 583216 421196 583228
rect 387024 583188 421196 583216
rect 387024 583176 387030 583188
rect 421190 583176 421196 583188
rect 421248 583176 421254 583228
rect 18966 583108 18972 583160
rect 19024 583148 19030 583160
rect 57974 583148 57980 583160
rect 19024 583120 57980 583148
rect 19024 583108 19030 583120
rect 57974 583108 57980 583120
rect 58032 583108 58038 583160
rect 112438 583108 112444 583160
rect 112496 583148 112502 583160
rect 142154 583148 142160 583160
rect 112496 583120 142160 583148
rect 112496 583108 112502 583120
rect 142154 583108 142160 583120
rect 142212 583108 142218 583160
rect 296622 583108 296628 583160
rect 296680 583148 296686 583160
rect 343174 583148 343180 583160
rect 296680 583120 343180 583148
rect 296680 583108 296686 583120
rect 343174 583108 343180 583120
rect 343232 583108 343238 583160
rect 368934 583108 368940 583160
rect 368992 583148 368998 583160
rect 423674 583148 423680 583160
rect 368992 583120 423680 583148
rect 368992 583108 368998 583120
rect 423674 583108 423680 583120
rect 423732 583108 423738 583160
rect 15102 583040 15108 583092
rect 15160 583080 15166 583092
rect 73154 583080 73160 583092
rect 15160 583052 73160 583080
rect 15160 583040 15166 583052
rect 73154 583040 73160 583052
rect 73212 583040 73218 583092
rect 107286 583040 107292 583092
rect 107344 583080 107350 583092
rect 139762 583080 139768 583092
rect 107344 583052 139768 583080
rect 107344 583040 107350 583052
rect 139762 583040 139768 583052
rect 139820 583040 139826 583092
rect 296530 583040 296536 583092
rect 296588 583080 296594 583092
rect 353478 583080 353484 583092
rect 296588 583052 353484 583080
rect 296588 583040 296594 583052
rect 353478 583040 353484 583052
rect 353536 583040 353542 583092
rect 366358 583040 366364 583092
rect 366416 583080 366422 583092
rect 425146 583080 425152 583092
rect 366416 583052 425152 583080
rect 366416 583040 366422 583052
rect 425146 583040 425152 583052
rect 425204 583040 425210 583092
rect 16390 582972 16396 583024
rect 16448 583012 16454 583024
rect 75914 583012 75920 583024
rect 16448 582984 75920 583012
rect 16448 582972 16454 582984
rect 75914 582972 75920 582984
rect 75972 582972 75978 583024
rect 104710 582972 104716 583024
rect 104768 583012 104774 583024
rect 138474 583012 138480 583024
rect 104768 582984 138480 583012
rect 104768 582972 104774 582984
rect 138474 582972 138480 582984
rect 138532 582972 138538 583024
rect 297726 582972 297732 583024
rect 297784 583012 297790 583024
rect 356054 583012 356060 583024
rect 297784 582984 356060 583012
rect 297784 582972 297790 582984
rect 356054 582972 356060 582984
rect 356112 582972 356118 583024
rect 363782 582972 363788 583024
rect 363840 583012 363846 583024
rect 423858 583012 423864 583024
rect 363840 582984 423864 583012
rect 363840 582972 363846 582984
rect 423858 582972 423864 582984
rect 423916 582972 423922 583024
rect 85574 544348 85580 544400
rect 85632 544388 85638 544400
rect 142430 544388 142436 544400
rect 85632 544360 142436 544388
rect 85632 544348 85638 544360
rect 142430 544348 142436 544360
rect 142488 544348 142494 544400
rect 247034 544348 247040 544400
rect 247092 544388 247098 544400
rect 378134 544388 378140 544400
rect 247092 544360 378140 544388
rect 247092 544348 247098 544360
rect 378134 544348 378140 544360
rect 378192 544348 378198 544400
rect 71038 542988 71044 543040
rect 71096 543028 71102 543040
rect 262214 543028 262220 543040
rect 71096 543000 262220 543028
rect 71096 542988 71102 543000
rect 262214 542988 262220 543000
rect 262272 542988 262278 543040
rect 100754 542036 100760 542088
rect 100812 542076 100818 542088
rect 140958 542076 140964 542088
rect 100812 542048 140964 542076
rect 100812 542036 100818 542048
rect 140958 542036 140964 542048
rect 141016 542036 141022 542088
rect 96614 541968 96620 542020
rect 96672 542008 96678 542020
rect 142246 542008 142252 542020
rect 96672 541980 142252 542008
rect 96672 541968 96678 541980
rect 142246 541968 142252 541980
rect 142304 541968 142310 542020
rect 93854 541900 93860 541952
rect 93912 541940 93918 541952
rect 142338 541940 142344 541952
rect 93912 541912 142344 541940
rect 93912 541900 93918 541912
rect 142338 541900 142344 541912
rect 142396 541900 142402 541952
rect 17586 541832 17592 541884
rect 17644 541872 17650 541884
rect 59354 541872 59360 541884
rect 17644 541844 59360 541872
rect 17644 541832 17650 541844
rect 59354 541832 59360 541844
rect 59412 541832 59418 541884
rect 91094 541832 91100 541884
rect 91152 541872 91158 541884
rect 140866 541872 140872 541884
rect 91152 541844 140872 541872
rect 91152 541832 91158 541844
rect 140866 541832 140872 541844
rect 140924 541832 140930 541884
rect 380894 541832 380900 541884
rect 380952 541872 380958 541884
rect 421098 541872 421104 541884
rect 380952 541844 421104 541872
rect 380952 541832 380958 541844
rect 421098 541832 421104 541844
rect 421156 541832 421162 541884
rect 18874 541764 18880 541816
rect 18932 541804 18938 541816
rect 62114 541804 62120 541816
rect 18932 541776 62120 541804
rect 18932 541764 18938 541776
rect 62114 541764 62120 541776
rect 62172 541764 62178 541816
rect 82814 541764 82820 541816
rect 82872 541804 82878 541816
rect 142522 541804 142528 541816
rect 82872 541776 142528 541804
rect 82872 541764 82878 541776
rect 142522 541764 142528 541776
rect 142580 541764 142586 541816
rect 375374 541764 375380 541816
rect 375432 541804 375438 541816
rect 422386 541804 422392 541816
rect 375432 541776 422392 541804
rect 375432 541764 375438 541776
rect 422386 541764 422392 541776
rect 422444 541764 422450 541816
rect 20254 541696 20260 541748
rect 20312 541736 20318 541748
rect 64874 541736 64880 541748
rect 20312 541708 64880 541736
rect 20312 541696 20318 541708
rect 64874 541696 64880 541708
rect 64932 541696 64938 541748
rect 80054 541696 80060 541748
rect 80112 541736 80118 541748
rect 141050 541736 141056 541748
rect 80112 541708 141056 541736
rect 80112 541696 80118 541708
rect 141050 541696 141056 541708
rect 141108 541696 141114 541748
rect 297818 541696 297824 541748
rect 297876 541736 297882 541748
rect 345014 541736 345020 541748
rect 297876 541708 345020 541736
rect 297876 541696 297882 541708
rect 345014 541696 345020 541708
rect 345072 541696 345078 541748
rect 373994 541696 374000 541748
rect 374052 541736 374058 541748
rect 422478 541736 422484 541748
rect 374052 541708 422484 541736
rect 374052 541696 374058 541708
rect 422478 541696 422484 541708
rect 422536 541696 422542 541748
rect 16482 541628 16488 541680
rect 16540 541668 16546 541680
rect 77294 541668 77300 541680
rect 16540 541640 77300 541668
rect 16540 541628 16546 541640
rect 77294 541628 77300 541640
rect 77352 541628 77358 541680
rect 97994 541628 98000 541680
rect 98052 541668 98058 541680
rect 245654 541668 245660 541680
rect 98052 541640 245660 541668
rect 98052 541628 98058 541640
rect 245654 541628 245660 541640
rect 245712 541628 245718 541680
rect 263594 541628 263600 541680
rect 263652 541668 263658 541680
rect 348418 541668 348424 541680
rect 263652 541640 348424 541668
rect 263652 541628 263658 541640
rect 348418 541628 348424 541640
rect 348476 541628 348482 541680
rect 371234 541628 371240 541680
rect 371292 541668 371298 541680
rect 421282 541668 421288 541680
rect 371292 541640 421288 541668
rect 371292 541628 371298 541640
rect 421282 541628 421288 541640
rect 421340 541628 421346 541680
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 7558 514808 7564 514820
rect 3384 514780 7564 514808
rect 3384 514768 3390 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 420822 470568 420828 470620
rect 420880 470608 420886 470620
rect 579982 470608 579988 470620
rect 420880 470580 579988 470608
rect 420880 470568 420886 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 421190 465400 421196 465452
rect 421248 465400 421254 465452
rect 421208 465236 421236 465400
rect 421282 465236 421288 465248
rect 421208 465208 421288 465236
rect 421282 465196 421288 465208
rect 421340 465196 421346 465248
rect 421098 463060 421104 463072
rect 389146 463032 421104 463060
rect 389146 462992 389174 463032
rect 421098 463020 421104 463032
rect 421156 463060 421162 463072
rect 425054 463060 425060 463072
rect 421156 463032 425060 463060
rect 421156 463020 421162 463032
rect 425054 463020 425060 463032
rect 425112 463020 425118 463072
rect 421190 462992 421196 463004
rect 386386 462964 389174 462992
rect 393286 462964 421196 462992
rect 386386 462720 386414 462964
rect 393286 462924 393314 462964
rect 421190 462952 421196 462964
rect 421248 462952 421254 463004
rect 382108 462692 386414 462720
rect 389146 462896 393314 462924
rect 382108 462664 382136 462692
rect 20714 462612 20720 462664
rect 20772 462652 20778 462664
rect 21634 462652 21640 462664
rect 20772 462624 21640 462652
rect 20772 462612 20778 462624
rect 21634 462612 21640 462624
rect 21692 462612 21698 462664
rect 298922 462612 298928 462664
rect 298980 462652 298986 462664
rect 301222 462652 301228 462664
rect 298980 462624 301228 462652
rect 298980 462612 298986 462624
rect 301222 462612 301228 462624
rect 301280 462652 301286 462664
rect 314654 462652 314660 462664
rect 301280 462624 314660 462652
rect 301280 462612 301286 462624
rect 314654 462612 314660 462624
rect 314712 462612 314718 462664
rect 382090 462612 382096 462664
rect 382148 462612 382154 462664
rect 385494 462612 385500 462664
rect 385552 462652 385558 462664
rect 389146 462652 389174 462896
rect 385552 462624 389174 462652
rect 385552 462612 385558 462624
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 419626 462408 419632 462460
rect 419684 462408 419690 462460
rect 419644 462380 419672 462408
rect 419644 462352 419764 462380
rect 299106 462272 299112 462324
rect 299164 462312 299170 462324
rect 300394 462312 300400 462324
rect 299164 462284 300400 462312
rect 299164 462272 299170 462284
rect 300394 462272 300400 462284
rect 300452 462272 300458 462324
rect 418798 462272 418804 462324
rect 418856 462312 418862 462324
rect 419626 462312 419632 462324
rect 418856 462284 419632 462312
rect 418856 462272 418862 462284
rect 419626 462272 419632 462284
rect 419684 462272 419690 462324
rect 419736 462312 419764 462352
rect 421190 462340 421196 462392
rect 421248 462380 421254 462392
rect 423766 462380 423772 462392
rect 421248 462352 423772 462380
rect 421248 462340 421254 462352
rect 423766 462340 423772 462352
rect 423824 462340 423830 462392
rect 421098 462312 421104 462324
rect 419736 462284 421104 462312
rect 20622 462204 20628 462256
rect 20680 462244 20686 462256
rect 24210 462244 24216 462256
rect 20680 462216 24216 462244
rect 20680 462204 20686 462216
rect 24210 462204 24216 462216
rect 24268 462204 24274 462256
rect 418154 462204 418160 462256
rect 418212 462244 418218 462256
rect 419718 462244 419724 462256
rect 418212 462216 419724 462244
rect 418212 462204 418218 462216
rect 419718 462204 419724 462216
rect 419776 462204 419782 462256
rect 418062 462136 418068 462188
rect 418120 462176 418126 462188
rect 419828 462176 419856 462284
rect 421098 462272 421104 462284
rect 421156 462272 421162 462324
rect 418120 462148 419856 462176
rect 418120 462136 418126 462148
rect 418430 461728 418436 461780
rect 418488 461768 418494 461780
rect 419810 461768 419816 461780
rect 418488 461740 419816 461768
rect 418488 461728 418494 461740
rect 419810 461728 419816 461740
rect 419868 461728 419874 461780
rect 348602 461252 348608 461304
rect 348660 461292 348666 461304
rect 350534 461292 350540 461304
rect 348660 461264 350540 461292
rect 348660 461252 348666 461264
rect 350534 461252 350540 461264
rect 350592 461252 350598 461304
rect 115014 461116 115020 461168
rect 115072 461156 115078 461168
rect 140774 461156 140780 461168
rect 115072 461128 140780 461156
rect 115072 461116 115078 461128
rect 140774 461116 140780 461128
rect 140832 461116 140838 461168
rect 86356 461048 86362 461100
rect 86414 461088 86420 461100
rect 142430 461088 142436 461100
rect 86414 461060 142436 461088
rect 86414 461048 86420 461060
rect 142430 461048 142436 461060
rect 142488 461088 142494 461100
rect 143534 461088 143540 461100
rect 142488 461060 143540 461088
rect 142488 461048 142494 461060
rect 143534 461048 143540 461060
rect 143592 461048 143598 461100
rect 376662 461048 376668 461100
rect 376720 461088 376726 461100
rect 383562 461088 383568 461100
rect 376720 461060 383568 461088
rect 376720 461048 376726 461060
rect 383562 461048 383568 461060
rect 383620 461048 383626 461100
rect 83780 460980 83786 461032
rect 83838 461020 83844 461032
rect 142522 461020 142528 461032
rect 83838 460992 142528 461020
rect 83838 460980 83844 460992
rect 142522 460980 142528 460992
rect 142580 460980 142586 461032
rect 300394 460980 300400 461032
rect 300452 461020 300458 461032
rect 319990 461020 319996 461032
rect 300452 460992 319996 461020
rect 300452 460980 300458 460992
rect 319990 460980 319996 460992
rect 320048 460980 320054 461032
rect 371510 460980 371516 461032
rect 371568 461020 371574 461032
rect 385494 461020 385500 461032
rect 371568 460992 385500 461020
rect 371568 460980 371574 460992
rect 385494 460980 385500 460992
rect 385552 460980 385558 461032
rect 16482 460912 16488 460964
rect 16540 460952 16546 460964
rect 78306 460952 78312 460964
rect 16540 460924 78312 460952
rect 16540 460912 16546 460924
rect 78306 460912 78312 460924
rect 78364 460912 78370 460964
rect 81342 460912 81348 460964
rect 81400 460952 81406 460964
rect 141050 460952 141056 460964
rect 81400 460924 141056 460952
rect 81400 460912 81406 460924
rect 141050 460912 141056 460924
rect 141108 460952 141114 460964
rect 142062 460952 142068 460964
rect 141108 460924 142068 460952
rect 141108 460912 141114 460924
rect 142062 460912 142068 460924
rect 142120 460912 142126 460964
rect 301406 460912 301412 460964
rect 301464 460952 301470 460964
rect 332870 460952 332876 460964
rect 301464 460924 332876 460952
rect 301464 460912 301470 460924
rect 332870 460912 332876 460924
rect 332928 460912 332934 460964
rect 374086 460912 374092 460964
rect 374144 460952 374150 460964
rect 374144 460924 379514 460952
rect 374144 460912 374150 460924
rect 298002 460844 298008 460896
rect 298060 460884 298066 460896
rect 302694 460884 302700 460896
rect 298060 460856 302700 460884
rect 298060 460844 298066 460856
rect 302694 460844 302700 460856
rect 302752 460884 302758 460896
rect 358630 460884 358636 460896
rect 302752 460856 358636 460884
rect 302752 460844 302758 460856
rect 358630 460844 358636 460856
rect 358688 460844 358694 460896
rect 379486 460884 379514 460924
rect 404998 460912 405004 460964
rect 405056 460952 405062 460964
rect 418522 460952 418528 460964
rect 405056 460924 418528 460952
rect 405056 460912 405062 460924
rect 418522 460912 418528 460924
rect 418580 460952 418586 460964
rect 421006 460952 421012 460964
rect 418580 460924 421012 460952
rect 418580 460912 418586 460924
rect 421006 460912 421012 460924
rect 421064 460912 421070 460964
rect 422478 460884 422484 460896
rect 379486 460856 422484 460884
rect 422478 460844 422484 460856
rect 422536 460844 422542 460896
rect 383562 460776 383568 460828
rect 383620 460816 383626 460828
rect 422386 460816 422392 460828
rect 383620 460788 422392 460816
rect 383620 460776 383626 460788
rect 422386 460776 422392 460788
rect 422444 460776 422450 460828
rect 298830 460164 298836 460216
rect 298888 460204 298894 460216
rect 345750 460204 345756 460216
rect 298888 460176 345756 460204
rect 298888 460164 298894 460176
rect 345750 460164 345756 460176
rect 345808 460164 345814 460216
rect 297818 459892 297824 459944
rect 297876 459932 297882 459944
rect 298830 459932 298836 459944
rect 297876 459904 298836 459932
rect 297876 459892 297882 459904
rect 298830 459892 298836 459904
rect 298888 459892 298894 459944
rect 415210 459620 415216 459672
rect 415268 459660 415274 459672
rect 419534 459660 419540 459672
rect 415268 459632 419540 459660
rect 415268 459620 415274 459632
rect 419534 459620 419540 459632
rect 419592 459620 419598 459672
rect 418430 459592 418436 459604
rect 400232 459564 418436 459592
rect 41414 459484 41420 459536
rect 41472 459524 41478 459536
rect 47394 459524 47400 459536
rect 41472 459496 47400 459524
rect 41472 459484 41478 459496
rect 47394 459484 47400 459496
rect 47452 459484 47458 459536
rect 68646 459484 68652 459536
rect 68704 459524 68710 459536
rect 71038 459524 71044 459536
rect 68704 459496 71044 459524
rect 68704 459484 68710 459496
rect 71038 459484 71044 459496
rect 71096 459484 71102 459536
rect 135622 459484 135628 459536
rect 135680 459524 135686 459536
rect 138382 459524 138388 459536
rect 135680 459496 138388 459524
rect 135680 459484 135686 459496
rect 138382 459484 138388 459496
rect 138440 459484 138446 459536
rect 297910 459484 297916 459536
rect 297968 459524 297974 459536
rect 340598 459524 340604 459536
rect 297968 459496 340604 459524
rect 297968 459484 297974 459496
rect 340598 459484 340604 459496
rect 340656 459484 340662 459536
rect 397270 459484 397276 459536
rect 397328 459524 397334 459536
rect 400232 459524 400260 459564
rect 418430 459552 418436 459564
rect 418488 459552 418494 459604
rect 422386 459552 422392 459604
rect 422444 459592 422450 459604
rect 423950 459592 423956 459604
rect 422444 459564 423956 459592
rect 422444 459552 422450 459564
rect 423950 459552 423956 459564
rect 424008 459552 424014 459604
rect 397328 459496 400260 459524
rect 397328 459484 397334 459496
rect 402422 459484 402428 459536
rect 402480 459524 402486 459536
rect 407022 459524 407028 459536
rect 402480 459496 407028 459524
rect 402480 459484 402486 459496
rect 407022 459484 407028 459496
rect 407080 459484 407086 459536
rect 407574 459484 407580 459536
rect 407632 459524 407638 459536
rect 415210 459524 415216 459536
rect 407632 459496 415216 459524
rect 407632 459484 407638 459496
rect 415210 459484 415216 459496
rect 415268 459484 415274 459536
rect 415302 459484 415308 459536
rect 415360 459524 415366 459536
rect 418062 459524 418068 459536
rect 415360 459496 418068 459524
rect 415360 459484 415366 459496
rect 418062 459484 418068 459496
rect 418120 459484 418126 459536
rect 17310 459416 17316 459468
rect 17368 459456 17374 459468
rect 60274 459456 60280 459468
rect 17368 459428 60280 459456
rect 17368 459416 17374 459428
rect 60274 459416 60280 459428
rect 60332 459416 60338 459468
rect 94406 459416 94412 459468
rect 94464 459456 94470 459468
rect 142338 459456 142344 459468
rect 94464 459428 142344 459456
rect 94464 459416 94470 459428
rect 142338 459416 142344 459428
rect 142396 459416 142402 459468
rect 300486 459416 300492 459468
rect 300544 459456 300550 459468
rect 330294 459456 330300 459468
rect 300544 459428 330300 459456
rect 300544 459416 300550 459428
rect 330294 459416 330300 459428
rect 330352 459416 330358 459468
rect 392118 459416 392124 459468
rect 392176 459456 392182 459468
rect 422570 459456 422576 459468
rect 392176 459428 422576 459456
rect 392176 459416 392182 459428
rect 422570 459416 422576 459428
rect 422628 459416 422634 459468
rect 18966 459348 18972 459400
rect 19024 459388 19030 459400
rect 57974 459388 57980 459400
rect 19024 459360 57980 459388
rect 19024 459348 19030 459360
rect 57974 459348 57980 459360
rect 58032 459348 58038 459400
rect 102042 459348 102048 459400
rect 102100 459388 102106 459400
rect 140958 459388 140964 459400
rect 102100 459360 140964 459388
rect 102100 459348 102106 459360
rect 140958 459348 140964 459360
rect 141016 459348 141022 459400
rect 299106 459348 299112 459400
rect 299164 459388 299170 459400
rect 325142 459388 325148 459400
rect 299164 459360 325148 459388
rect 299164 459348 299170 459360
rect 325142 459348 325148 459360
rect 325200 459348 325206 459400
rect 410150 459348 410156 459400
rect 410208 459388 410214 459400
rect 419718 459388 419724 459400
rect 410208 459360 419724 459388
rect 410208 459348 410214 459360
rect 419718 459348 419724 459360
rect 419776 459348 419782 459400
rect 17678 459280 17684 459332
rect 17736 459320 17742 459332
rect 49970 459320 49976 459332
rect 17736 459292 49976 459320
rect 17736 459280 17742 459292
rect 49970 459280 49976 459292
rect 50028 459280 50034 459332
rect 91830 459280 91836 459332
rect 91888 459320 91894 459332
rect 140866 459320 140872 459332
rect 91888 459292 140872 459320
rect 91888 459280 91894 459292
rect 140866 459280 140872 459292
rect 140924 459280 140930 459332
rect 363782 459280 363788 459332
rect 363840 459320 363846 459332
rect 423858 459320 423864 459332
rect 363840 459292 423864 459320
rect 363840 459280 363846 459292
rect 423858 459280 423864 459292
rect 423916 459280 423922 459332
rect 19058 459212 19064 459264
rect 19116 459252 19122 459264
rect 23198 459252 23204 459264
rect 19116 459224 23204 459252
rect 19116 459212 19122 459224
rect 23198 459212 23204 459224
rect 23256 459252 23262 459264
rect 44818 459252 44824 459264
rect 23256 459224 44824 459252
rect 23256 459212 23262 459224
rect 44818 459212 44824 459224
rect 44876 459212 44882 459264
rect 417878 459212 417884 459264
rect 417936 459252 417942 459264
rect 421466 459252 421472 459264
rect 417936 459224 421472 459252
rect 417936 459212 417942 459224
rect 421466 459212 421472 459224
rect 421524 459212 421530 459264
rect 20254 459144 20260 459196
rect 20312 459184 20318 459196
rect 65426 459184 65432 459196
rect 20312 459156 65432 459184
rect 20312 459144 20318 459156
rect 65426 459144 65432 459156
rect 65484 459144 65490 459196
rect 300394 459144 300400 459196
rect 300452 459184 300458 459196
rect 300670 459184 300676 459196
rect 300452 459156 300676 459184
rect 300452 459144 300458 459156
rect 300670 459144 300676 459156
rect 300728 459144 300734 459196
rect 39114 459076 39120 459128
rect 39172 459116 39178 459128
rect 42242 459116 42248 459128
rect 39172 459088 42248 459116
rect 39172 459076 39178 459088
rect 42242 459076 42248 459088
rect 42300 459076 42306 459128
rect 112438 459008 112444 459060
rect 112496 459048 112502 459060
rect 141142 459048 141148 459060
rect 112496 459020 141148 459048
rect 112496 459008 112502 459020
rect 141142 459008 141148 459020
rect 141200 459048 141206 459060
rect 142154 459048 142160 459060
rect 141200 459020 142160 459048
rect 141200 459008 141206 459020
rect 142154 459008 142160 459020
rect 142212 459008 142218 459060
rect 300394 459008 300400 459060
rect 300452 459048 300458 459060
rect 327718 459048 327724 459060
rect 300452 459020 327724 459048
rect 300452 459008 300458 459020
rect 327718 459008 327724 459020
rect 327776 459008 327782 459060
rect 399846 459008 399852 459060
rect 399904 459048 399910 459060
rect 409874 459048 409880 459060
rect 399904 459020 409880 459048
rect 399904 459008 399910 459020
rect 409874 459008 409880 459020
rect 409932 459008 409938 459060
rect 96982 458940 96988 458992
rect 97040 458980 97046 458992
rect 140866 458980 140872 458992
rect 97040 458952 140872 458980
rect 97040 458940 97046 458952
rect 140866 458940 140872 458952
rect 140924 458940 140930 458992
rect 296622 458940 296628 458992
rect 296680 458980 296686 458992
rect 297910 458980 297916 458992
rect 296680 458952 297916 458980
rect 296680 458940 296686 458952
rect 297910 458940 297916 458952
rect 297968 458980 297974 458992
rect 343174 458980 343180 458992
rect 297968 458952 343180 458980
rect 297968 458940 297974 458952
rect 343174 458940 343180 458952
rect 343232 458940 343238 458992
rect 394694 458940 394700 458992
rect 394752 458980 394758 458992
rect 419810 458980 419816 458992
rect 394752 458952 419816 458980
rect 394752 458940 394758 458952
rect 419810 458940 419816 458952
rect 419868 458980 419874 458992
rect 420914 458980 420920 458992
rect 419868 458952 420920 458980
rect 419868 458940 419874 458952
rect 420914 458940 420920 458952
rect 420972 458940 420978 458992
rect 89254 458872 89260 458924
rect 89312 458912 89318 458924
rect 135714 458912 135720 458924
rect 89312 458884 135720 458912
rect 89312 458872 89318 458884
rect 135714 458872 135720 458884
rect 135772 458872 135778 458924
rect 296530 458872 296536 458924
rect 296588 458912 296594 458924
rect 297542 458912 297548 458924
rect 296588 458884 297548 458912
rect 296588 458872 296594 458884
rect 297542 458872 297548 458884
rect 297600 458912 297606 458924
rect 353478 458912 353484 458924
rect 297600 458884 353484 458912
rect 297600 458872 297606 458884
rect 353478 458872 353484 458884
rect 353536 458872 353542 458924
rect 366358 458872 366364 458924
rect 366416 458912 366422 458924
rect 418154 458912 418160 458924
rect 366416 458884 418160 458912
rect 366416 458872 366422 458884
rect 418154 458872 418160 458884
rect 418212 458872 418218 458924
rect 15102 458804 15108 458856
rect 15160 458844 15166 458856
rect 16206 458844 16212 458856
rect 15160 458816 16212 458844
rect 15160 458804 15166 458816
rect 16206 458804 16212 458816
rect 16264 458844 16270 458856
rect 73154 458844 73160 458856
rect 16264 458816 73160 458844
rect 16264 458804 16270 458816
rect 73154 458804 73160 458816
rect 73212 458804 73218 458856
rect 99282 458804 99288 458856
rect 99340 458844 99346 458856
rect 244274 458844 244280 458856
rect 99340 458816 244280 458844
rect 99340 458804 99346 458816
rect 244274 458804 244280 458816
rect 244332 458804 244338 458856
rect 264974 458804 264980 458856
rect 265032 458844 265038 458856
rect 348326 458844 348332 458856
rect 265032 458816 348332 458844
rect 265032 458804 265038 458816
rect 348326 458804 348332 458816
rect 348384 458804 348390 458856
rect 368934 458804 368940 458856
rect 368992 458844 368998 458856
rect 420914 458844 420920 458856
rect 368992 458816 420920 458844
rect 368992 458804 368998 458816
rect 420914 458804 420920 458816
rect 420972 458804 420978 458856
rect 140866 458736 140872 458788
rect 140924 458776 140930 458788
rect 141050 458776 141056 458788
rect 140924 458748 141056 458776
rect 140924 458736 140930 458748
rect 141050 458736 141056 458748
rect 141108 458776 141114 458788
rect 142246 458776 142252 458788
rect 141108 458748 142252 458776
rect 141108 458736 141114 458748
rect 142246 458736 142252 458748
rect 142304 458736 142310 458788
rect 140958 458192 140964 458244
rect 141016 458232 141022 458244
rect 141234 458232 141240 458244
rect 141016 458204 141240 458232
rect 141016 458192 141022 458204
rect 141234 458192 141240 458204
rect 141292 458192 141298 458244
rect 297634 458192 297640 458244
rect 297692 458232 297698 458244
rect 300486 458232 300492 458244
rect 297692 458204 300492 458232
rect 297692 458192 297698 458204
rect 300486 458192 300492 458204
rect 300544 458192 300550 458244
rect 19242 458124 19248 458176
rect 19300 458164 19306 458176
rect 34514 458164 34520 458176
rect 19300 458136 34520 458164
rect 19300 458124 19306 458136
rect 34514 458124 34520 458136
rect 34572 458124 34578 458176
rect 107286 458124 107292 458176
rect 107344 458164 107350 458176
rect 139762 458164 139768 458176
rect 107344 458136 139768 458164
rect 107344 458124 107350 458136
rect 139762 458124 139768 458136
rect 139820 458124 139826 458176
rect 299290 458124 299296 458176
rect 299348 458164 299354 458176
rect 322566 458164 322572 458176
rect 299348 458136 322572 458164
rect 299348 458124 299354 458136
rect 322566 458124 322572 458136
rect 322624 458124 322630 458176
rect 384390 458124 384396 458176
rect 384448 458164 384454 458176
rect 418062 458164 418068 458176
rect 384448 458136 418068 458164
rect 384448 458124 384454 458136
rect 418062 458124 418068 458136
rect 418120 458124 418126 458176
rect 418154 458124 418160 458176
rect 418212 458164 418218 458176
rect 418798 458164 418804 458176
rect 418212 458136 418804 458164
rect 418212 458124 418218 458136
rect 418798 458124 418804 458136
rect 418856 458164 418862 458176
rect 425146 458164 425152 458176
rect 418856 458136 425152 458164
rect 418856 458124 418862 458136
rect 425146 458124 425152 458136
rect 425204 458124 425210 458176
rect 21266 458056 21272 458108
rect 21324 458096 21330 458108
rect 26786 458096 26792 458108
rect 21324 458068 26792 458096
rect 21324 458056 21330 458068
rect 26786 458056 26792 458068
rect 26844 458056 26850 458108
rect 117222 458056 117228 458108
rect 117280 458096 117286 458108
rect 139670 458096 139676 458108
rect 117280 458068 139676 458096
rect 117280 458056 117286 458068
rect 139670 458056 139676 458068
rect 139728 458056 139734 458108
rect 299382 458056 299388 458108
rect 299440 458096 299446 458108
rect 317414 458096 317420 458108
rect 299440 458068 317420 458096
rect 299440 458056 299446 458068
rect 317414 458056 317420 458068
rect 317472 458056 317478 458108
rect 409874 458056 409880 458108
rect 409932 458096 409938 458108
rect 418338 458096 418344 458108
rect 409932 458068 418344 458096
rect 409932 458056 409938 458068
rect 418338 458056 418344 458068
rect 418396 458056 418402 458108
rect 420914 458056 420920 458108
rect 420972 458096 420978 458108
rect 421558 458096 421564 458108
rect 420972 458068 421564 458096
rect 420972 458056 420978 458068
rect 421558 458056 421564 458068
rect 421616 458096 421622 458108
rect 423674 458096 423680 458108
rect 421616 458068 423680 458096
rect 421616 458056 421622 458068
rect 423674 458056 423680 458068
rect 423732 458056 423738 458108
rect 125318 457988 125324 458040
rect 125376 458028 125382 458040
rect 139394 458028 139400 458040
rect 125376 458000 139400 458028
rect 125376 457988 125382 458000
rect 139394 457988 139400 458000
rect 139452 457988 139458 458040
rect 130470 457920 130476 457972
rect 130528 457960 130534 457972
rect 139578 457960 139584 457972
rect 130528 457932 139584 457960
rect 130528 457920 130534 457932
rect 139578 457920 139584 457932
rect 139636 457920 139642 457972
rect 21358 457648 21364 457700
rect 21416 457688 21422 457700
rect 31938 457688 31944 457700
rect 21416 457660 31944 457688
rect 21416 457648 21422 457660
rect 31938 457648 31944 457660
rect 31996 457648 32002 457700
rect 300578 457648 300584 457700
rect 300636 457688 300642 457700
rect 301222 457688 301228 457700
rect 300636 457660 301228 457688
rect 300636 457648 300642 457660
rect 301222 457648 301228 457660
rect 301280 457648 301286 457700
rect 17862 457580 17868 457632
rect 17920 457620 17926 457632
rect 17920 457592 26234 457620
rect 17920 457580 17926 457592
rect 19058 457512 19064 457564
rect 19116 457552 19122 457564
rect 21358 457552 21364 457564
rect 19116 457524 21364 457552
rect 19116 457512 19122 457524
rect 21358 457512 21364 457524
rect 21416 457512 21422 457564
rect 26206 457552 26234 457592
rect 37182 457552 37188 457564
rect 26206 457524 37188 457552
rect 37182 457512 37188 457524
rect 37240 457512 37246 457564
rect 20530 457444 20536 457496
rect 20588 457484 20594 457496
rect 21266 457484 21272 457496
rect 20588 457456 21272 457484
rect 20588 457444 20594 457456
rect 21266 457444 21272 457456
rect 21324 457444 21330 457496
rect 39114 457484 39120 457496
rect 26206 457456 39120 457484
rect 17770 457376 17776 457428
rect 17828 457416 17834 457428
rect 20438 457416 20444 457428
rect 17828 457388 20444 457416
rect 17828 457376 17834 457388
rect 20438 457376 20444 457388
rect 20496 457416 20502 457428
rect 26206 457416 26234 457456
rect 39114 457444 39120 457456
rect 39172 457444 39178 457496
rect 301222 457444 301228 457496
rect 301280 457484 301286 457496
rect 312262 457484 312268 457496
rect 301280 457456 312268 457484
rect 301280 457444 301286 457456
rect 312262 457444 312268 457456
rect 312320 457444 312326 457496
rect 20496 457388 26234 457416
rect 20496 457376 20502 457388
rect 139670 457104 139676 457156
rect 139728 457144 139734 457156
rect 139946 457144 139952 457156
rect 139728 457116 139952 457144
rect 139728 457104 139734 457116
rect 139946 457104 139952 457116
rect 140004 457104 140010 457156
rect 419534 457036 419540 457088
rect 419592 457076 419598 457088
rect 419810 457076 419816 457088
rect 419592 457048 419816 457076
rect 419592 457036 419598 457048
rect 419810 457036 419816 457048
rect 419868 457036 419874 457088
rect 139394 456832 139400 456884
rect 139452 456872 139458 456884
rect 140038 456872 140044 456884
rect 139452 456844 140044 456872
rect 139452 456832 139458 456844
rect 140038 456832 140044 456844
rect 140096 456832 140102 456884
rect 17862 456764 17868 456816
rect 17920 456804 17926 456816
rect 18874 456804 18880 456816
rect 17920 456776 18880 456804
rect 17920 456764 17926 456776
rect 18874 456764 18880 456776
rect 18932 456764 18938 456816
rect 18966 456764 18972 456816
rect 19024 456804 19030 456816
rect 19242 456804 19248 456816
rect 19024 456776 19248 456804
rect 19024 456764 19030 456776
rect 19242 456764 19248 456776
rect 19300 456764 19306 456816
rect 139578 456764 139584 456816
rect 139636 456804 139642 456816
rect 139762 456804 139768 456816
rect 139636 456776 139768 456804
rect 139636 456764 139642 456776
rect 139762 456764 139768 456776
rect 139820 456764 139826 456816
rect 299014 456764 299020 456816
rect 299072 456804 299078 456816
rect 299290 456804 299296 456816
rect 299072 456776 299296 456804
rect 299072 456764 299078 456776
rect 299290 456764 299296 456776
rect 299348 456764 299354 456816
rect 418246 456764 418252 456816
rect 418304 456804 418310 456816
rect 418522 456804 418528 456816
rect 418304 456776 418528 456804
rect 418304 456764 418310 456776
rect 418522 456764 418528 456776
rect 418580 456764 418586 456816
rect 300854 456696 300860 456748
rect 300912 456736 300918 456748
rect 301498 456736 301504 456748
rect 300912 456708 301504 456736
rect 300912 456696 300918 456708
rect 301498 456696 301504 456708
rect 301556 456736 301562 456748
rect 361206 456736 361212 456748
rect 301556 456708 361212 456736
rect 301556 456696 301562 456708
rect 361206 456696 361212 456708
rect 361264 456696 361270 456748
rect 297726 456628 297732 456680
rect 297784 456668 297790 456680
rect 356054 456668 356060 456680
rect 297784 456640 356060 456668
rect 297784 456628 297790 456640
rect 356054 456628 356060 456640
rect 356112 456628 356118 456680
rect 16390 455336 16396 455388
rect 16448 455376 16454 455388
rect 17862 455376 17868 455388
rect 16448 455348 17868 455376
rect 16448 455336 16454 455348
rect 17862 455336 17868 455348
rect 17920 455336 17926 455388
rect 17586 454656 17592 454708
rect 17644 454696 17650 454708
rect 17862 454696 17868 454708
rect 17644 454668 17868 454696
rect 17644 454656 17650 454668
rect 17862 454656 17868 454668
rect 17920 454696 17926 454708
rect 75914 454696 75920 454708
rect 17920 454668 75920 454696
rect 17920 454656 17926 454668
rect 75914 454656 75920 454668
rect 75972 454656 75978 454708
rect 248414 416032 248420 416084
rect 248472 416072 248478 416084
rect 378134 416072 378140 416084
rect 248472 416044 378140 416072
rect 248472 416032 248478 416044
rect 378134 416032 378140 416044
rect 378192 416032 378198 416084
rect 71038 413244 71044 413296
rect 71096 413284 71102 413296
rect 260834 413284 260840 413296
rect 71096 413256 260840 413284
rect 71096 413244 71102 413256
rect 260834 413244 260840 413256
rect 260892 413244 260898 413296
rect 2774 410048 2780 410100
rect 2832 410088 2838 410100
rect 4982 410088 4988 410100
rect 2832 410060 4988 410088
rect 2832 410048 2838 410060
rect 4982 410048 4988 410060
rect 5040 410048 5046 410100
rect 3694 398828 3700 398880
rect 3752 398868 3758 398880
rect 19978 398868 19984 398880
rect 3752 398840 19984 398868
rect 3752 398828 3758 398840
rect 19978 398828 19984 398840
rect 20036 398828 20042 398880
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 20070 345080 20076 345092
rect 3384 345052 20076 345080
rect 3384 345040 3390 345052
rect 20070 345040 20076 345052
rect 20128 345040 20134 345092
rect 16298 333208 16304 333260
rect 16356 333248 16362 333260
rect 18782 333248 18788 333260
rect 16356 333220 18788 333248
rect 16356 333208 16362 333220
rect 18782 333208 18788 333220
rect 18840 333248 18846 333260
rect 57698 333248 57704 333260
rect 18840 333220 57704 333248
rect 18840 333208 18846 333220
rect 57698 333208 57704 333220
rect 57756 333208 57762 333260
rect 96982 333004 96988 333056
rect 97040 333044 97046 333056
rect 141050 333044 141056 333056
rect 97040 333016 141056 333044
rect 97040 333004 97046 333016
rect 141050 333004 141056 333016
rect 141108 333004 141114 333056
rect 115014 332936 115020 332988
rect 115072 332976 115078 332988
rect 140774 332976 140780 332988
rect 115072 332948 140780 332976
rect 115072 332936 115078 332948
rect 140774 332936 140780 332948
rect 140832 332976 140838 332988
rect 142154 332976 142160 332988
rect 140832 332948 142160 332976
rect 140832 332936 140838 332948
rect 142154 332936 142160 332948
rect 142212 332936 142218 332988
rect 15010 332868 15016 332920
rect 15068 332908 15074 332920
rect 17770 332908 17776 332920
rect 15068 332880 17776 332908
rect 15068 332868 15074 332880
rect 17770 332868 17776 332880
rect 17828 332908 17834 332920
rect 47394 332908 47400 332920
rect 17828 332880 47400 332908
rect 17828 332868 17834 332880
rect 47394 332868 47400 332880
rect 47452 332868 47458 332920
rect 91830 332868 91836 332920
rect 91888 332908 91894 332920
rect 140866 332908 140872 332920
rect 91888 332880 140872 332908
rect 91888 332868 91894 332880
rect 140866 332868 140872 332880
rect 140924 332868 140930 332920
rect 300670 332868 300676 332920
rect 300728 332908 300734 332920
rect 318794 332908 318800 332920
rect 300728 332880 318800 332908
rect 300728 332868 300734 332880
rect 318794 332868 318800 332880
rect 318852 332908 318858 332920
rect 319990 332908 319996 332920
rect 318852 332880 319996 332908
rect 318852 332868 318858 332880
rect 319990 332868 319996 332880
rect 320048 332868 320054 332920
rect 17678 332800 17684 332852
rect 17736 332840 17742 332852
rect 49970 332840 49976 332852
rect 17736 332812 49976 332840
rect 17736 332800 17742 332812
rect 49970 332800 49976 332812
rect 50028 332800 50034 332852
rect 112438 332800 112444 332852
rect 112496 332840 112502 332852
rect 141142 332840 141148 332852
rect 112496 332812 141148 332840
rect 112496 332800 112502 332812
rect 141142 332800 141148 332812
rect 141200 332800 141206 332852
rect 299014 332800 299020 332852
rect 299072 332840 299078 332852
rect 321554 332840 321560 332852
rect 299072 332812 321560 332840
rect 299072 332800 299078 332812
rect 321554 332800 321560 332812
rect 321612 332840 321618 332852
rect 322566 332840 322572 332852
rect 321612 332812 322572 332840
rect 321612 332800 321618 332812
rect 322566 332800 322572 332812
rect 322624 332800 322630 332852
rect 327258 332840 327264 332852
rect 325666 332812 327264 332840
rect 16390 332732 16396 332784
rect 16448 332772 16454 332784
rect 73154 332772 73160 332784
rect 16448 332744 73160 332772
rect 16448 332732 16454 332744
rect 73154 332732 73160 332744
rect 73212 332732 73218 332784
rect 107286 332732 107292 332784
rect 107344 332772 107350 332784
rect 139302 332772 139308 332784
rect 107344 332744 139308 332772
rect 107344 332732 107350 332744
rect 139302 332732 139308 332744
rect 139360 332732 139366 332784
rect 299106 332732 299112 332784
rect 299164 332772 299170 332784
rect 324314 332772 324320 332784
rect 299164 332744 324320 332772
rect 299164 332732 299170 332744
rect 324314 332732 324320 332744
rect 324372 332772 324378 332784
rect 325142 332772 325148 332784
rect 324372 332744 325148 332772
rect 324372 332732 324378 332744
rect 325142 332732 325148 332744
rect 325200 332732 325206 332784
rect 17402 332664 17408 332716
rect 17460 332704 17466 332716
rect 17586 332704 17592 332716
rect 17460 332676 17592 332704
rect 17460 332664 17466 332676
rect 17586 332664 17592 332676
rect 17644 332704 17650 332716
rect 75914 332704 75920 332716
rect 17644 332676 75920 332704
rect 17644 332664 17650 332676
rect 75914 332664 75920 332676
rect 75972 332664 75978 332716
rect 109862 332664 109868 332716
rect 109920 332704 109926 332716
rect 142246 332704 142252 332716
rect 109920 332676 142252 332704
rect 109920 332664 109926 332676
rect 142246 332664 142252 332676
rect 142304 332664 142310 332716
rect 300394 332664 300400 332716
rect 300452 332704 300458 332716
rect 325666 332704 325694 332812
rect 327258 332800 327264 332812
rect 327316 332800 327322 332852
rect 416682 332840 416688 332852
rect 373966 332812 416688 332840
rect 373966 332772 373994 332812
rect 416682 332800 416688 332812
rect 416740 332840 416746 332852
rect 418798 332840 418804 332852
rect 416740 332812 418804 332840
rect 416740 332800 416746 332812
rect 418798 332800 418804 332812
rect 418856 332800 418862 332852
rect 300452 332676 325694 332704
rect 369780 332744 373994 332772
rect 300452 332664 300458 332676
rect 16482 332596 16488 332648
rect 16540 332636 16546 332648
rect 78306 332636 78312 332648
rect 16540 332608 78312 332636
rect 16540 332596 16546 332608
rect 78306 332596 78312 332608
rect 78364 332596 78370 332648
rect 104710 332596 104716 332648
rect 104768 332636 104774 332648
rect 138290 332636 138296 332648
rect 104768 332608 138296 332636
rect 104768 332596 104774 332608
rect 138290 332596 138296 332608
rect 138348 332636 138354 332648
rect 138566 332636 138572 332648
rect 138348 332608 138572 332636
rect 138348 332596 138354 332608
rect 138566 332596 138572 332608
rect 138624 332596 138630 332648
rect 297634 332596 297640 332648
rect 297692 332636 297698 332648
rect 329834 332636 329840 332648
rect 297692 332608 329840 332636
rect 297692 332596 297698 332608
rect 329834 332596 329840 332608
rect 329892 332596 329898 332648
rect 3602 332528 3608 332580
rect 3660 332568 3666 332580
rect 21634 332568 21640 332580
rect 3660 332540 21640 332568
rect 3660 332528 3666 332540
rect 21634 332528 21640 332540
rect 21692 332528 21698 332580
rect 68646 332528 68652 332580
rect 68704 332568 68710 332580
rect 71038 332568 71044 332580
rect 68704 332540 71044 332568
rect 68704 332528 68710 332540
rect 71038 332528 71044 332540
rect 71096 332528 71102 332580
rect 94406 332528 94412 332580
rect 94464 332568 94470 332580
rect 96522 332568 96528 332580
rect 94464 332540 96528 332568
rect 94464 332528 94470 332540
rect 96522 332528 96528 332540
rect 96580 332528 96586 332580
rect 135622 332528 135628 332580
rect 135680 332568 135686 332580
rect 138382 332568 138388 332580
rect 135680 332540 138388 332568
rect 135680 332528 135686 332540
rect 138382 332528 138388 332540
rect 138440 332528 138446 332580
rect 300302 332528 300308 332580
rect 300360 332568 300366 332580
rect 307110 332568 307116 332580
rect 300360 332540 307116 332568
rect 300360 332528 300366 332540
rect 307110 332528 307116 332540
rect 307168 332528 307174 332580
rect 335446 332568 335452 332580
rect 311084 332540 335452 332568
rect 19150 332460 19156 332512
rect 19208 332500 19214 332512
rect 39666 332500 39672 332512
rect 19208 332472 39672 332500
rect 19208 332460 19214 332472
rect 39666 332460 39672 332472
rect 39724 332460 39730 332512
rect 119982 332460 119988 332512
rect 120040 332500 120046 332512
rect 139762 332500 139768 332512
rect 120040 332472 139768 332500
rect 120040 332460 120046 332472
rect 139762 332460 139768 332472
rect 139820 332460 139826 332512
rect 303522 332460 303528 332512
rect 303580 332500 303586 332512
rect 310974 332500 310980 332512
rect 303580 332472 310980 332500
rect 303580 332460 303586 332472
rect 310974 332460 310980 332472
rect 311032 332460 311038 332512
rect 18874 332392 18880 332444
rect 18932 332432 18938 332444
rect 37274 332432 37280 332444
rect 18932 332404 37280 332432
rect 18932 332392 18938 332404
rect 37274 332392 37280 332404
rect 37332 332392 37338 332444
rect 122650 332392 122656 332444
rect 122708 332432 122714 332444
rect 138750 332432 138756 332444
rect 122708 332404 138756 332432
rect 122708 332392 122714 332404
rect 138750 332392 138756 332404
rect 138808 332392 138814 332444
rect 301314 332392 301320 332444
rect 301372 332432 301378 332444
rect 311084 332432 311112 332540
rect 335446 332528 335452 332540
rect 335504 332528 335510 332580
rect 348326 332528 348332 332580
rect 348384 332568 348390 332580
rect 350902 332568 350908 332580
rect 348384 332540 350908 332568
rect 348384 332528 348390 332540
rect 350902 332528 350908 332540
rect 350960 332528 350966 332580
rect 366358 332528 366364 332580
rect 366416 332568 366422 332580
rect 369780 332568 369808 332744
rect 386506 332732 386512 332784
rect 386564 332772 386570 332784
rect 421190 332772 421196 332784
rect 386564 332744 421196 332772
rect 386564 332732 386570 332744
rect 421190 332732 421196 332744
rect 421248 332732 421254 332784
rect 371510 332664 371516 332716
rect 371568 332704 371574 332716
rect 371568 332676 373994 332704
rect 371568 332664 371574 332676
rect 373966 332636 373994 332676
rect 383654 332664 383660 332716
rect 383712 332704 383718 332716
rect 384390 332704 384396 332716
rect 383712 332676 384396 332704
rect 383712 332664 383718 332676
rect 384390 332664 384396 332676
rect 384448 332704 384454 332716
rect 418522 332704 418528 332716
rect 384448 332676 418528 332704
rect 384448 332664 384454 332676
rect 418522 332664 418528 332676
rect 418580 332664 418586 332716
rect 423766 332636 423772 332648
rect 373966 332608 423772 332636
rect 423766 332596 423772 332608
rect 423824 332636 423830 332648
rect 424042 332636 424048 332648
rect 423824 332608 424048 332636
rect 423824 332596 423830 332608
rect 424042 332596 424048 332608
rect 424100 332596 424106 332648
rect 366416 332540 369808 332568
rect 366416 332528 366422 332540
rect 415302 332528 415308 332580
rect 415360 332568 415366 332580
rect 421098 332568 421104 332580
rect 415360 332540 421104 332568
rect 415360 332528 415366 332540
rect 421098 332528 421104 332540
rect 421156 332528 421162 332580
rect 338022 332500 338028 332512
rect 311268 332472 338028 332500
rect 301372 332404 311112 332432
rect 301372 332392 301378 332404
rect 311158 332392 311164 332444
rect 311216 332432 311222 332444
rect 311268 332432 311296 332472
rect 338022 332460 338028 332472
rect 338080 332460 338086 332512
rect 399846 332460 399852 332512
rect 399904 332500 399910 332512
rect 418430 332500 418436 332512
rect 399904 332472 418436 332500
rect 399904 332460 399910 332472
rect 418430 332460 418436 332472
rect 418488 332460 418494 332512
rect 332870 332432 332876 332444
rect 311216 332404 311296 332432
rect 316006 332404 332876 332432
rect 311216 332392 311222 332404
rect 21266 332324 21272 332376
rect 21324 332364 21330 332376
rect 26786 332364 26792 332376
rect 21324 332336 26792 332364
rect 21324 332324 21330 332336
rect 26786 332324 26792 332336
rect 26844 332324 26850 332376
rect 27522 332324 27528 332376
rect 27580 332364 27586 332376
rect 44818 332364 44824 332376
rect 27580 332336 44824 332364
rect 27580 332324 27586 332336
rect 44818 332324 44824 332336
rect 44876 332324 44882 332376
rect 125318 332324 125324 332376
rect 125376 332364 125382 332376
rect 140038 332364 140044 332376
rect 125376 332336 140044 332364
rect 125376 332324 125382 332336
rect 140038 332324 140044 332336
rect 140096 332324 140102 332376
rect 301038 332324 301044 332376
rect 301096 332364 301102 332376
rect 312262 332364 312268 332376
rect 301096 332336 312268 332364
rect 301096 332324 301102 332336
rect 312262 332324 312268 332336
rect 312320 332324 312326 332376
rect 18966 332256 18972 332308
rect 19024 332296 19030 332308
rect 34514 332296 34520 332308
rect 19024 332268 34520 332296
rect 19024 332256 19030 332268
rect 34514 332256 34520 332268
rect 34572 332256 34578 332308
rect 127894 332256 127900 332308
rect 127952 332296 127958 332308
rect 138842 332296 138848 332308
rect 127952 332268 138848 332296
rect 127952 332256 127958 332268
rect 138842 332256 138848 332268
rect 138900 332256 138906 332308
rect 301406 332256 301412 332308
rect 301464 332296 301470 332308
rect 316006 332296 316034 332404
rect 332870 332392 332876 332404
rect 332928 332392 332934 332444
rect 402422 332392 402428 332444
rect 402480 332432 402486 332444
rect 418706 332432 418712 332444
rect 402480 332404 418712 332432
rect 402480 332392 402486 332404
rect 418706 332392 418712 332404
rect 418764 332392 418770 332444
rect 407574 332324 407580 332376
rect 407632 332364 407638 332376
rect 419626 332364 419632 332376
rect 407632 332336 419632 332364
rect 407632 332324 407638 332336
rect 419626 332324 419632 332336
rect 419684 332324 419690 332376
rect 301464 332268 316034 332296
rect 301464 332256 301470 332268
rect 410150 332256 410156 332308
rect 410208 332296 410214 332308
rect 419902 332296 419908 332308
rect 410208 332268 419908 332296
rect 410208 332256 410214 332268
rect 419902 332256 419908 332268
rect 419960 332256 419966 332308
rect 19058 332188 19064 332240
rect 19116 332228 19122 332240
rect 31938 332228 31944 332240
rect 19116 332200 31944 332228
rect 19116 332188 19122 332200
rect 31938 332188 31944 332200
rect 31996 332188 32002 332240
rect 130470 332188 130476 332240
rect 130528 332228 130534 332240
rect 139670 332228 139676 332240
rect 130528 332200 139676 332228
rect 130528 332188 130534 332200
rect 139670 332188 139676 332200
rect 139728 332188 139734 332240
rect 397270 332188 397276 332240
rect 397328 332228 397334 332240
rect 418614 332228 418620 332240
rect 397328 332200 418620 332228
rect 397328 332188 397334 332200
rect 418614 332188 418620 332200
rect 418672 332188 418678 332240
rect 20346 332120 20352 332172
rect 20404 332160 20410 332172
rect 29362 332160 29368 332172
rect 20404 332132 29368 332160
rect 20404 332120 20410 332132
rect 29362 332120 29368 332132
rect 29420 332120 29426 332172
rect 117222 332120 117228 332172
rect 117280 332160 117286 332172
rect 139946 332160 139952 332172
rect 117280 332132 139952 332160
rect 117280 332120 117286 332132
rect 139946 332120 139952 332132
rect 140004 332120 140010 332172
rect 300578 332120 300584 332172
rect 300636 332160 300642 332172
rect 309686 332160 309692 332172
rect 300636 332132 309692 332160
rect 300636 332120 300642 332132
rect 309686 332120 309692 332132
rect 309744 332120 309750 332172
rect 20530 332052 20536 332104
rect 20588 332092 20594 332104
rect 42242 332092 42248 332104
rect 20588 332064 42248 332092
rect 20588 332052 20594 332064
rect 42242 332052 42248 332064
rect 42300 332052 42306 332104
rect 306742 331916 306748 331968
rect 306800 331956 306806 331968
rect 314838 331956 314844 331968
rect 306800 331928 314844 331956
rect 306800 331916 306806 331928
rect 314838 331916 314844 331928
rect 314896 331916 314902 331968
rect 266354 331848 266360 331900
rect 266412 331888 266418 331900
rect 348326 331888 348332 331900
rect 266412 331860 348332 331888
rect 266412 331848 266418 331860
rect 348326 331848 348332 331860
rect 348384 331848 348390 331900
rect 350534 331848 350540 331900
rect 350592 331888 350598 331900
rect 358630 331888 358636 331900
rect 350592 331860 358636 331888
rect 350592 331848 350598 331860
rect 358630 331848 358636 331860
rect 358688 331848 358694 331900
rect 404998 331848 405004 331900
rect 405056 331888 405062 331900
rect 419442 331888 419448 331900
rect 405056 331860 419448 331888
rect 405056 331848 405062 331860
rect 419442 331848 419448 331860
rect 419500 331848 419506 331900
rect 139486 331576 139492 331628
rect 139544 331616 139550 331628
rect 139946 331616 139952 331628
rect 139544 331588 139952 331616
rect 139544 331576 139550 331588
rect 139946 331576 139952 331588
rect 140004 331576 140010 331628
rect 376662 331372 376668 331424
rect 376720 331412 376726 331424
rect 382458 331412 382464 331424
rect 376720 331384 382464 331412
rect 376720 331372 376726 331384
rect 382458 331372 382464 331384
rect 382516 331372 382522 331424
rect 418614 331304 418620 331356
rect 418672 331344 418678 331356
rect 420086 331344 420092 331356
rect 418672 331316 420092 331344
rect 418672 331304 418678 331316
rect 420086 331304 420092 331316
rect 420144 331304 420150 331356
rect 19242 331236 19248 331288
rect 19300 331276 19306 331288
rect 20346 331276 20352 331288
rect 19300 331248 20352 331276
rect 19300 331236 19306 331248
rect 20346 331236 20352 331248
rect 20404 331236 20410 331288
rect 89254 331236 89260 331288
rect 89312 331276 89318 331288
rect 91002 331276 91008 331288
rect 89312 331248 91008 331276
rect 89312 331236 89318 331248
rect 91002 331236 91008 331248
rect 91060 331236 91066 331288
rect 138750 331236 138756 331288
rect 138808 331276 138814 331288
rect 139578 331276 139584 331288
rect 138808 331248 139584 331276
rect 138808 331236 138814 331248
rect 139578 331236 139584 331248
rect 139636 331236 139642 331288
rect 300210 331236 300216 331288
rect 300268 331276 300274 331288
rect 301406 331276 301412 331288
rect 300268 331248 301412 331276
rect 300268 331236 300274 331248
rect 301406 331236 301412 331248
rect 301464 331236 301470 331288
rect 311894 331236 311900 331288
rect 311952 331276 311958 331288
rect 317414 331276 317420 331288
rect 311952 331248 317420 331276
rect 311952 331236 311958 331248
rect 317414 331236 317420 331248
rect 317472 331236 317478 331288
rect 368934 331236 368940 331288
rect 368992 331276 368998 331288
rect 373258 331276 373264 331288
rect 368992 331248 373264 331276
rect 368992 331236 368998 331248
rect 373258 331236 373264 331248
rect 373316 331236 373322 331288
rect 374086 331236 374092 331288
rect 374144 331276 374150 331288
rect 379422 331276 379428 331288
rect 374144 331248 379428 331276
rect 374144 331236 374150 331248
rect 379422 331236 379428 331248
rect 379480 331236 379486 331288
rect 381814 331236 381820 331288
rect 381872 331276 381878 331288
rect 386322 331276 386328 331288
rect 381872 331248 386328 331276
rect 381872 331236 381878 331248
rect 386322 331236 386328 331248
rect 386380 331236 386386 331288
rect 418430 331236 418436 331288
rect 418488 331276 418494 331288
rect 419994 331276 420000 331288
rect 418488 331248 420000 331276
rect 418488 331236 418494 331248
rect 419994 331236 420000 331248
rect 420052 331236 420058 331288
rect 303522 331168 303528 331220
rect 303580 331208 303586 331220
rect 350534 331208 350540 331220
rect 303580 331180 350540 331208
rect 303580 331168 303586 331180
rect 350534 331168 350540 331180
rect 350592 331168 350598 331220
rect 363782 331168 363788 331220
rect 363840 331208 363846 331220
rect 363840 331180 412634 331208
rect 363840 331168 363846 331180
rect 299290 331100 299296 331152
rect 299348 331140 299354 331152
rect 311894 331140 311900 331152
rect 299348 331112 311900 331140
rect 299348 331100 299354 331112
rect 311894 331100 311900 331112
rect 311952 331100 311958 331152
rect 412606 331072 412634 331180
rect 418798 331100 418804 331152
rect 418856 331140 418862 331152
rect 419626 331140 419632 331152
rect 418856 331112 419632 331140
rect 418856 331100 418862 331112
rect 419626 331100 419632 331112
rect 419684 331100 419690 331152
rect 423766 331072 423772 331084
rect 412606 331044 423772 331072
rect 423766 331032 423772 331044
rect 423824 331032 423830 331084
rect 139486 330964 139492 331016
rect 139544 331004 139550 331016
rect 140038 331004 140044 331016
rect 139544 330976 140044 331004
rect 139544 330964 139550 330976
rect 140038 330964 140044 330976
rect 140096 330964 140102 331016
rect 419442 330964 419448 331016
rect 419500 331004 419506 331016
rect 421006 331004 421012 331016
rect 419500 330976 421012 331004
rect 419500 330964 419506 330976
rect 421006 330964 421012 330976
rect 421064 330964 421070 331016
rect 298830 330488 298836 330540
rect 298888 330528 298894 330540
rect 301222 330528 301228 330540
rect 298888 330500 301228 330528
rect 298888 330488 298894 330500
rect 301222 330488 301228 330500
rect 301280 330528 301286 330540
rect 345750 330528 345756 330540
rect 301280 330500 345756 330528
rect 301280 330488 301286 330500
rect 345750 330488 345756 330500
rect 345808 330488 345814 330540
rect 20180 329820 21128 329848
rect 17586 329740 17592 329792
rect 17644 329780 17650 329792
rect 20180 329780 20208 329820
rect 17644 329752 20208 329780
rect 17644 329740 17650 329752
rect 20254 329740 20260 329792
rect 20312 329780 20318 329792
rect 20990 329780 20996 329792
rect 20312 329752 20996 329780
rect 20312 329740 20318 329752
rect 20990 329740 20996 329752
rect 21048 329740 21054 329792
rect 21100 329780 21128 329820
rect 62850 329780 62856 329792
rect 21100 329752 62856 329780
rect 62850 329740 62856 329752
rect 62908 329740 62914 329792
rect 84010 329740 84016 329792
rect 84068 329780 84074 329792
rect 142430 329780 142436 329792
rect 84068 329752 142436 329780
rect 84068 329740 84074 329752
rect 142430 329740 142436 329752
rect 142488 329740 142494 329792
rect 382458 329740 382464 329792
rect 382516 329780 382522 329792
rect 417418 329780 417424 329792
rect 382516 329752 417424 329780
rect 382516 329740 382522 329752
rect 417418 329740 417424 329752
rect 417476 329740 417482 329792
rect 419810 329740 419816 329792
rect 419868 329780 419874 329792
rect 421558 329780 421564 329792
rect 419868 329752 421564 329780
rect 419868 329740 419874 329752
rect 421558 329740 421564 329752
rect 421616 329740 421622 329792
rect 21008 329712 21036 329740
rect 65426 329712 65432 329724
rect 21008 329684 65432 329712
rect 65426 329672 65432 329684
rect 65484 329672 65490 329724
rect 102134 329672 102140 329724
rect 102192 329712 102198 329724
rect 140958 329712 140964 329724
rect 102192 329684 140964 329712
rect 102192 329672 102198 329684
rect 140958 329672 140964 329684
rect 141016 329712 141022 329724
rect 142522 329712 142528 329724
rect 141016 329684 142528 329712
rect 141016 329672 141022 329684
rect 142522 329672 142528 329684
rect 142580 329672 142586 329724
rect 386322 329672 386328 329724
rect 386380 329712 386386 329724
rect 425054 329712 425060 329724
rect 386380 329684 425060 329712
rect 386380 329672 386386 329684
rect 425054 329672 425060 329684
rect 425112 329672 425118 329724
rect 16206 329604 16212 329656
rect 16264 329644 16270 329656
rect 17310 329644 17316 329656
rect 16264 329616 17316 329644
rect 16264 329604 16270 329616
rect 17310 329604 17316 329616
rect 17368 329644 17374 329656
rect 60274 329644 60280 329656
rect 17368 329616 60280 329644
rect 17368 329604 17374 329616
rect 60274 329604 60280 329616
rect 60332 329604 60338 329656
rect 392118 329604 392124 329656
rect 392176 329644 392182 329656
rect 393222 329644 393228 329656
rect 392176 329616 393228 329644
rect 392176 329604 392182 329616
rect 393222 329604 393228 329616
rect 393280 329644 393286 329656
rect 393314 329644 393320 329656
rect 393280 329616 393320 329644
rect 393280 329604 393286 329616
rect 393314 329604 393320 329616
rect 393372 329604 393378 329656
rect 422662 329644 422668 329656
rect 393424 329616 422668 329644
rect 389542 329536 389548 329588
rect 389600 329576 389606 329588
rect 390462 329576 390468 329588
rect 389600 329548 390468 329576
rect 389600 329536 389606 329548
rect 390462 329536 390468 329548
rect 390520 329576 390526 329588
rect 393424 329576 393452 329616
rect 422662 329604 422668 329616
rect 422720 329604 422726 329656
rect 390520 329548 393452 329576
rect 390520 329536 390526 329548
rect 393498 329536 393504 329588
rect 393556 329576 393562 329588
rect 422570 329576 422576 329588
rect 393556 329548 422576 329576
rect 393556 329536 393562 329548
rect 422570 329536 422576 329548
rect 422628 329536 422634 329588
rect 402946 329480 412634 329508
rect 394694 329400 394700 329452
rect 394752 329440 394758 329452
rect 395982 329440 395988 329452
rect 394752 329412 395988 329440
rect 394752 329400 394758 329412
rect 395982 329400 395988 329412
rect 396040 329440 396046 329452
rect 402946 329440 402974 329480
rect 396040 329412 402974 329440
rect 412606 329440 412634 329480
rect 417418 329468 417424 329520
rect 417476 329508 417482 329520
rect 423674 329508 423680 329520
rect 417476 329480 423680 329508
rect 417476 329468 417482 329480
rect 423674 329468 423680 329480
rect 423732 329508 423738 329520
rect 423950 329508 423956 329520
rect 423732 329480 423956 329508
rect 423732 329468 423738 329480
rect 423950 329468 423956 329480
rect 424008 329468 424014 329520
rect 419534 329440 419540 329452
rect 412606 329412 419540 329440
rect 396040 329400 396046 329412
rect 419534 329400 419540 329412
rect 419592 329400 419598 329452
rect 91002 329196 91008 329248
rect 91060 329236 91066 329248
rect 138658 329236 138664 329248
rect 91060 329208 138664 329236
rect 91060 329196 91066 329208
rect 138658 329196 138664 329208
rect 138716 329196 138722 329248
rect 86678 329128 86684 329180
rect 86736 329168 86742 329180
rect 140774 329168 140780 329180
rect 86736 329140 140780 329168
rect 86736 329128 86742 329140
rect 140774 329128 140780 329140
rect 140832 329128 140838 329180
rect 412726 329128 412732 329180
rect 412784 329168 412790 329180
rect 422478 329168 422484 329180
rect 412784 329140 422484 329168
rect 412784 329128 412790 329140
rect 422478 329128 422484 329140
rect 422536 329128 422542 329180
rect 81342 329060 81348 329112
rect 81400 329100 81406 329112
rect 141510 329100 141516 329112
rect 81400 329072 141516 329100
rect 81400 329060 81406 329072
rect 141510 329060 141516 329072
rect 141568 329060 141574 329112
rect 373258 329060 373264 329112
rect 373316 329100 373322 329112
rect 419810 329100 419816 329112
rect 373316 329072 419816 329100
rect 373316 329060 373322 329072
rect 419810 329060 419816 329072
rect 419868 329060 419874 329112
rect 140774 327700 140780 327752
rect 140832 327740 140838 327752
rect 142062 327740 142068 327752
rect 140832 327712 142068 327740
rect 140832 327700 140838 327712
rect 142062 327700 142068 327712
rect 142120 327740 142126 327752
rect 143534 327740 143540 327752
rect 142120 327712 143540 327740
rect 142120 327700 142126 327712
rect 143534 327700 143540 327712
rect 143592 327700 143598 327752
rect 140774 327564 140780 327616
rect 140832 327604 140838 327616
rect 141142 327604 141148 327616
rect 140832 327576 141148 327604
rect 140832 327564 140838 327576
rect 141142 327564 141148 327576
rect 141200 327564 141206 327616
rect 3602 318792 3608 318844
rect 3660 318832 3666 318844
rect 17218 318832 17224 318844
rect 3660 318804 17224 318832
rect 3660 318792 3666 318804
rect 17218 318792 17224 318804
rect 17276 318792 17282 318844
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4890 292856 4896 292868
rect 2832 292828 4896 292856
rect 2832 292816 2838 292828
rect 4890 292816 4896 292828
rect 4948 292816 4954 292868
rect 300762 288328 300768 288380
rect 300820 288368 300826 288380
rect 360194 288368 360200 288380
rect 300820 288340 360200 288368
rect 300820 288328 300826 288340
rect 360194 288328 360200 288340
rect 360252 288328 360258 288380
rect 297726 288260 297732 288312
rect 297784 288300 297790 288312
rect 356054 288300 356060 288312
rect 297784 288272 356060 288300
rect 297784 288260 297790 288272
rect 356054 288260 356060 288272
rect 356112 288260 356118 288312
rect 249794 287648 249800 287700
rect 249852 287688 249858 287700
rect 378134 287688 378140 287700
rect 249852 287660 378140 287688
rect 249852 287648 249858 287660
rect 378134 287648 378140 287660
rect 378192 287648 378198 287700
rect 296622 287036 296628 287088
rect 296680 287076 296686 287088
rect 297726 287076 297732 287088
rect 296680 287048 297732 287076
rect 296680 287036 296686 287048
rect 297726 287036 297732 287048
rect 297784 287036 297790 287088
rect 297818 285608 297824 285660
rect 297876 285648 297882 285660
rect 342254 285648 342260 285660
rect 297876 285620 342260 285648
rect 297876 285608 297882 285620
rect 342254 285608 342260 285620
rect 342312 285608 342318 285660
rect 298002 285540 298008 285592
rect 298060 285580 298066 285592
rect 339494 285580 339500 285592
rect 298060 285552 339500 285580
rect 298060 285540 298066 285552
rect 339494 285540 339500 285552
rect 339552 285540 339558 285592
rect 395982 285268 395988 285320
rect 396040 285308 396046 285320
rect 423950 285308 423956 285320
rect 396040 285280 423956 285308
rect 396040 285268 396046 285280
rect 423950 285268 423956 285280
rect 424008 285268 424014 285320
rect 300394 285200 300400 285252
rect 300452 285240 300458 285252
rect 318794 285240 318800 285252
rect 300452 285212 318800 285240
rect 300452 285200 300458 285212
rect 318794 285200 318800 285212
rect 318852 285200 318858 285252
rect 393222 285200 393228 285252
rect 393280 285240 393286 285252
rect 422570 285240 422576 285252
rect 393280 285212 422576 285240
rect 393280 285200 393286 285212
rect 422570 285200 422576 285212
rect 422628 285200 422634 285252
rect 299198 285132 299204 285184
rect 299256 285172 299262 285184
rect 321554 285172 321560 285184
rect 299256 285144 321560 285172
rect 299256 285132 299262 285144
rect 321554 285132 321560 285144
rect 321612 285132 321618 285184
rect 390462 285132 390468 285184
rect 390520 285172 390526 285184
rect 421006 285172 421012 285184
rect 390520 285144 421012 285172
rect 390520 285132 390526 285144
rect 421006 285132 421012 285144
rect 421064 285132 421070 285184
rect 297910 285064 297916 285116
rect 297968 285104 297974 285116
rect 324314 285104 324320 285116
rect 297968 285076 324320 285104
rect 297968 285064 297974 285076
rect 324314 285064 324320 285076
rect 324372 285064 324378 285116
rect 383654 285064 383660 285116
rect 383712 285104 383718 285116
rect 418246 285104 418252 285116
rect 383712 285076 418252 285104
rect 383712 285064 383718 285076
rect 418246 285064 418252 285076
rect 418304 285064 418310 285116
rect 136634 284996 136640 285048
rect 136692 285036 136698 285048
rect 296070 285036 296076 285048
rect 136692 285008 296076 285036
rect 136692 284996 136698 285008
rect 296070 284996 296076 285008
rect 296128 284996 296134 285048
rect 299014 284996 299020 285048
rect 299072 285036 299078 285048
rect 327074 285036 327080 285048
rect 299072 285008 327080 285036
rect 299072 284996 299078 285008
rect 327074 284996 327080 285008
rect 327132 284996 327138 285048
rect 386414 284996 386420 285048
rect 386472 285036 386478 285048
rect 421190 285036 421196 285048
rect 386472 285008 421196 285036
rect 386472 284996 386478 285008
rect 421190 284996 421196 285008
rect 421248 284996 421254 285048
rect 71038 284928 71044 284980
rect 71096 284968 71102 284980
rect 258074 284968 258080 284980
rect 71096 284940 258080 284968
rect 71096 284928 71102 284940
rect 258074 284928 258080 284940
rect 258132 284928 258138 284980
rect 299106 284928 299112 284980
rect 299164 284968 299170 284980
rect 329834 284968 329840 284980
rect 299164 284940 329840 284968
rect 299164 284928 299170 284940
rect 329834 284928 329840 284940
rect 329892 284928 329898 284980
rect 379422 284928 379428 284980
rect 379480 284968 379486 284980
rect 425146 284968 425152 284980
rect 379480 284940 425152 284968
rect 379480 284928 379486 284940
rect 425146 284928 425152 284940
rect 425204 284928 425210 284980
rect 297726 284316 297732 284368
rect 297784 284356 297790 284368
rect 298002 284356 298008 284368
rect 297784 284328 298008 284356
rect 297784 284316 297790 284328
rect 298002 284316 298008 284328
rect 298060 284316 298066 284368
rect 416682 284316 416688 284368
rect 416740 284356 416746 284368
rect 418522 284356 418528 284368
rect 416740 284328 418528 284356
rect 416740 284316 416746 284328
rect 418522 284316 418528 284328
rect 418580 284316 418586 284368
rect 2774 266364 2780 266416
rect 2832 266404 2838 266416
rect 6178 266404 6184 266416
rect 2832 266376 6184 266404
rect 2832 266364 2838 266376
rect 6178 266364 6184 266376
rect 6236 266364 6242 266416
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 5074 240224 5080 240236
rect 2832 240196 5080 240224
rect 2832 240184 2838 240196
rect 5074 240184 5080 240196
rect 5132 240184 5138 240236
rect 2774 213936 2780 213988
rect 2832 213976 2838 213988
rect 6270 213976 6276 213988
rect 2832 213948 6276 213976
rect 2832 213936 2838 213948
rect 6270 213936 6276 213948
rect 6328 213936 6334 213988
rect 300946 206592 300952 206644
rect 301004 206632 301010 206644
rect 301130 206632 301136 206644
rect 301004 206604 301136 206632
rect 301004 206592 301010 206604
rect 301130 206592 301136 206604
rect 301188 206592 301194 206644
rect 301038 206456 301044 206508
rect 301096 206496 301102 206508
rect 301406 206496 301412 206508
rect 301096 206468 301412 206496
rect 301096 206456 301102 206468
rect 301406 206456 301412 206468
rect 301464 206456 301470 206508
rect 140774 206320 140780 206372
rect 140832 206360 140838 206372
rect 142062 206360 142068 206372
rect 140832 206332 142068 206360
rect 140832 206320 140838 206332
rect 142062 206320 142068 206332
rect 142120 206360 142126 206372
rect 143534 206360 143540 206372
rect 142120 206332 143540 206360
rect 142120 206320 142126 206332
rect 143534 206320 143540 206332
rect 143592 206320 143598 206372
rect 371602 206252 371608 206304
rect 371660 206292 371666 206304
rect 424042 206292 424048 206304
rect 371660 206264 424048 206292
rect 371660 206252 371666 206264
rect 424042 206252 424048 206264
rect 424100 206252 424106 206304
rect 141234 205572 141240 205624
rect 141292 205612 141298 205624
rect 142522 205612 142528 205624
rect 141292 205584 142528 205612
rect 141292 205572 141298 205584
rect 142522 205572 142528 205584
rect 142580 205572 142586 205624
rect 420914 205368 420920 205420
rect 420972 205408 420978 205420
rect 422662 205408 422668 205420
rect 420972 205380 422668 205408
rect 420972 205368 420978 205380
rect 422662 205368 422668 205380
rect 422720 205368 422726 205420
rect 419534 205068 419540 205080
rect 412606 205040 419540 205068
rect 298922 204892 298928 204944
rect 298980 204932 298986 204944
rect 300394 204932 300400 204944
rect 298980 204904 300400 204932
rect 298980 204892 298986 204904
rect 300394 204892 300400 204904
rect 300452 204932 300458 204944
rect 309042 204932 309048 204944
rect 300452 204904 309048 204932
rect 300452 204892 300458 204904
rect 309042 204892 309048 204904
rect 309100 204892 309106 204944
rect 297542 204824 297548 204876
rect 297600 204864 297606 204876
rect 299014 204864 299020 204876
rect 297600 204836 299020 204864
rect 297600 204824 297606 204836
rect 299014 204824 299020 204836
rect 299072 204824 299078 204876
rect 297910 204756 297916 204808
rect 297968 204796 297974 204808
rect 300302 204796 300308 204808
rect 297968 204768 300308 204796
rect 297968 204756 297974 204768
rect 300302 204756 300308 204768
rect 300360 204756 300366 204808
rect 298002 204688 298008 204740
rect 298060 204728 298066 204740
rect 299106 204728 299112 204740
rect 298060 204700 299112 204728
rect 298060 204688 298066 204700
rect 299106 204688 299112 204700
rect 299164 204688 299170 204740
rect 372614 204688 372620 204740
rect 372672 204728 372678 204740
rect 412606 204728 412634 205040
rect 419534 205028 419540 205040
rect 419592 205028 419598 205080
rect 423950 205000 423956 205012
rect 372672 204700 412634 204728
rect 417436 204972 423956 205000
rect 372672 204688 372678 204700
rect 86678 204620 86684 204672
rect 86736 204660 86742 204672
rect 140774 204660 140780 204672
rect 86736 204632 140780 204660
rect 86736 204620 86742 204632
rect 140774 204620 140780 204632
rect 140832 204620 140838 204672
rect 394694 204620 394700 204672
rect 394752 204660 394758 204672
rect 417436 204660 417464 204972
rect 423950 204960 423956 204972
rect 424008 205000 424014 205012
rect 425238 205000 425244 205012
rect 424008 204972 425244 205000
rect 424008 204960 424014 204972
rect 425238 204960 425244 204972
rect 425296 204960 425302 205012
rect 421558 204892 421564 204944
rect 421616 204932 421622 204944
rect 425146 204932 425152 204944
rect 421616 204904 425152 204932
rect 421616 204892 421622 204904
rect 425146 204892 425152 204904
rect 425204 204892 425210 204944
rect 418246 204688 418252 204740
rect 418304 204728 418310 204740
rect 418430 204728 418436 204740
rect 418304 204700 418436 204728
rect 418304 204688 418310 204700
rect 418430 204688 418436 204700
rect 418488 204688 418494 204740
rect 394752 204632 417464 204660
rect 394752 204620 394758 204632
rect 115014 204552 115020 204604
rect 115072 204592 115078 204604
rect 142154 204592 142160 204604
rect 115072 204564 142160 204592
rect 115072 204552 115078 204564
rect 142154 204552 142160 204564
rect 142212 204552 142218 204604
rect 301406 204552 301412 204604
rect 301464 204592 301470 204604
rect 365622 204592 365628 204604
rect 301464 204564 365628 204592
rect 301464 204552 301470 204564
rect 365622 204552 365628 204564
rect 365680 204552 365686 204604
rect 392118 204552 392124 204604
rect 392176 204592 392182 204604
rect 422570 204592 422576 204604
rect 392176 204564 422576 204592
rect 392176 204552 392182 204564
rect 422570 204552 422576 204564
rect 422628 204592 422634 204604
rect 424042 204592 424048 204604
rect 422628 204564 424048 204592
rect 422628 204552 422634 204564
rect 424042 204552 424048 204564
rect 424100 204552 424106 204604
rect 102042 204484 102048 204536
rect 102100 204524 102106 204536
rect 141234 204524 141240 204536
rect 102100 204496 141240 204524
rect 102100 204484 102106 204496
rect 141234 204484 141240 204496
rect 141292 204484 141298 204536
rect 300302 204484 300308 204536
rect 300360 204524 300366 204536
rect 325142 204524 325148 204536
rect 300360 204496 325148 204524
rect 300360 204484 300366 204496
rect 325142 204484 325148 204496
rect 325200 204484 325206 204536
rect 389542 204484 389548 204536
rect 389600 204524 389606 204536
rect 420914 204524 420920 204536
rect 389600 204496 420920 204524
rect 389600 204484 389606 204496
rect 420914 204484 420920 204496
rect 420972 204484 420978 204536
rect 96982 204416 96988 204468
rect 97040 204456 97046 204468
rect 141142 204456 141148 204468
rect 97040 204428 141148 204456
rect 97040 204416 97046 204428
rect 141142 204416 141148 204428
rect 141200 204416 141206 204468
rect 299014 204416 299020 204468
rect 299072 204456 299078 204468
rect 327718 204456 327724 204468
rect 299072 204428 327724 204456
rect 299072 204416 299078 204428
rect 327718 204416 327724 204428
rect 327776 204416 327782 204468
rect 386966 204416 386972 204468
rect 387024 204456 387030 204468
rect 421190 204456 421196 204468
rect 387024 204428 421196 204456
rect 387024 204416 387030 204428
rect 421190 204416 421196 204428
rect 421248 204416 421254 204468
rect 19058 204348 19064 204400
rect 19116 204388 19122 204400
rect 31938 204388 31944 204400
rect 19116 204360 31944 204388
rect 19116 204348 19122 204360
rect 31938 204348 31944 204360
rect 31996 204348 32002 204400
rect 94406 204348 94412 204400
rect 94464 204388 94470 204400
rect 142338 204388 142344 204400
rect 94464 204360 142344 204388
rect 94464 204348 94470 204360
rect 142338 204348 142344 204360
rect 142396 204348 142402 204400
rect 299106 204348 299112 204400
rect 299164 204388 299170 204400
rect 330294 204388 330300 204400
rect 299164 204360 330300 204388
rect 299164 204348 299170 204360
rect 330294 204348 330300 204360
rect 330352 204348 330358 204400
rect 384390 204348 384396 204400
rect 384448 204388 384454 204400
rect 418430 204388 418436 204400
rect 384448 204360 418436 204388
rect 384448 204348 384454 204360
rect 418430 204348 418436 204360
rect 418488 204348 418494 204400
rect 19150 204280 19156 204332
rect 19208 204320 19214 204332
rect 39666 204320 39672 204332
rect 19208 204292 39672 204320
rect 19208 204280 19214 204292
rect 39666 204280 39672 204292
rect 39724 204280 39730 204332
rect 138014 204280 138020 204332
rect 138072 204320 138078 204332
rect 138658 204320 138664 204332
rect 138072 204292 138664 204320
rect 138072 204280 138078 204292
rect 138658 204280 138664 204292
rect 138716 204320 138722 204332
rect 143626 204320 143632 204332
rect 138716 204292 143632 204320
rect 138716 204280 138722 204292
rect 143626 204280 143632 204292
rect 143684 204280 143690 204332
rect 295242 204280 295248 204332
rect 295300 204320 295306 204332
rect 297634 204320 297640 204332
rect 295300 204292 297640 204320
rect 295300 204280 295306 204292
rect 297634 204280 297640 204292
rect 297692 204320 297698 204332
rect 353478 204320 353484 204332
rect 297692 204292 353484 204320
rect 297692 204280 297698 204292
rect 353478 204280 353484 204292
rect 353536 204280 353542 204332
rect 374086 204280 374092 204332
rect 374144 204320 374150 204332
rect 421374 204320 421380 204332
rect 374144 204292 421380 204320
rect 374144 204280 374150 204292
rect 421374 204280 421380 204292
rect 421432 204320 421438 204332
rect 421558 204320 421564 204332
rect 421432 204292 421564 204320
rect 421432 204280 421438 204292
rect 421558 204280 421564 204292
rect 421616 204280 421622 204332
rect 7558 204212 7564 204264
rect 7616 204252 7622 204264
rect 21634 204252 21640 204264
rect 7616 204224 21640 204252
rect 7616 204212 7622 204224
rect 21634 204212 21640 204224
rect 21692 204212 21698 204264
rect 22002 204212 22008 204264
rect 22060 204252 22066 204264
rect 22060 204224 31064 204252
rect 22060 204212 22066 204224
rect 16206 204144 16212 204196
rect 16264 204184 16270 204196
rect 30926 204184 30932 204196
rect 16264 204156 30932 204184
rect 16264 204144 16270 204156
rect 30926 204144 30932 204156
rect 30984 204144 30990 204196
rect 21450 204076 21456 204128
rect 21508 204116 21514 204128
rect 26786 204116 26792 204128
rect 21508 204088 26792 204116
rect 21508 204076 21514 204088
rect 26786 204076 26792 204088
rect 26844 204076 26850 204128
rect 31036 204116 31064 204224
rect 68646 204212 68652 204264
rect 68704 204252 68710 204264
rect 70578 204252 70584 204264
rect 68704 204224 70584 204252
rect 68704 204212 68710 204224
rect 70578 204212 70584 204224
rect 70636 204252 70642 204264
rect 71038 204252 71044 204264
rect 70636 204224 71044 204252
rect 70636 204212 70642 204224
rect 71038 204212 71044 204224
rect 71096 204212 71102 204264
rect 127894 204212 127900 204264
rect 127952 204252 127958 204264
rect 130010 204252 130016 204264
rect 127952 204224 130016 204252
rect 127952 204212 127958 204224
rect 130010 204212 130016 204224
rect 130068 204212 130074 204264
rect 130470 204212 130476 204264
rect 130528 204252 130534 204264
rect 133782 204252 133788 204264
rect 130528 204224 133788 204252
rect 130528 204212 130534 204224
rect 133782 204212 133788 204224
rect 133840 204212 133846 204264
rect 307110 204252 307116 204264
rect 302528 204224 307116 204252
rect 31110 204144 31116 204196
rect 31168 204184 31174 204196
rect 60274 204184 60280 204196
rect 31168 204156 60280 204184
rect 31168 204144 31174 204156
rect 60274 204144 60280 204156
rect 60332 204144 60338 204196
rect 84010 204144 84016 204196
rect 84068 204184 84074 204196
rect 142430 204184 142436 204196
rect 84068 204156 142436 204184
rect 84068 204144 84074 204156
rect 142430 204144 142436 204156
rect 142488 204144 142494 204196
rect 299106 204144 299112 204196
rect 299164 204184 299170 204196
rect 299382 204184 299388 204196
rect 299164 204156 299388 204184
rect 299164 204144 299170 204156
rect 299382 204144 299388 204156
rect 299440 204144 299446 204196
rect 300578 204144 300584 204196
rect 300636 204184 300642 204196
rect 302528 204184 302556 204224
rect 307110 204212 307116 204224
rect 307168 204212 307174 204264
rect 309042 204212 309048 204264
rect 309100 204252 309106 204264
rect 319990 204252 319996 204264
rect 309100 204224 319996 204252
rect 309100 204212 309106 204224
rect 319990 204212 319996 204224
rect 320048 204212 320054 204264
rect 348326 204212 348332 204264
rect 348384 204252 348390 204264
rect 350902 204252 350908 204264
rect 348384 204224 350908 204252
rect 348384 204212 348390 204224
rect 350902 204212 350908 204224
rect 350960 204212 350966 204264
rect 368934 204212 368940 204264
rect 368992 204252 368998 204264
rect 372614 204252 372620 204264
rect 368992 204224 372620 204252
rect 368992 204212 368998 204224
rect 372614 204212 372620 204224
rect 372672 204212 372678 204264
rect 397270 204212 397276 204264
rect 397328 204252 397334 204264
rect 411254 204252 411260 204264
rect 397328 204224 411260 204252
rect 397328 204212 397334 204224
rect 411254 204212 411260 204224
rect 411312 204212 411318 204264
rect 415302 204212 415308 204264
rect 415360 204252 415366 204264
rect 416774 204252 416780 204264
rect 415360 204224 416780 204252
rect 415360 204212 415366 204224
rect 416774 204212 416780 204224
rect 416832 204212 416838 204264
rect 419626 204252 419632 204264
rect 418448 204224 419632 204252
rect 332870 204184 332876 204196
rect 300636 204156 302556 204184
rect 302620 204156 332876 204184
rect 300636 204144 300642 204156
rect 65426 204116 65432 204128
rect 31036 204088 65432 204116
rect 65426 204076 65432 204088
rect 65484 204076 65490 204128
rect 89254 204076 89260 204128
rect 89312 204116 89318 204128
rect 138014 204116 138020 204128
rect 89312 204088 138020 204116
rect 89312 204076 89318 204088
rect 138014 204076 138020 204088
rect 138072 204076 138078 204128
rect 300486 204076 300492 204128
rect 300544 204116 300550 204128
rect 302620 204116 302648 204156
rect 332870 204144 332876 204156
rect 332928 204144 332934 204196
rect 365622 204144 365628 204196
rect 365680 204184 365686 204196
rect 371510 204184 371516 204196
rect 365680 204156 371516 204184
rect 365680 204144 365686 204156
rect 371510 204144 371516 204156
rect 371568 204144 371574 204196
rect 402422 204144 402428 204196
rect 402480 204184 402486 204196
rect 418338 204184 418344 204196
rect 402480 204156 418344 204184
rect 402480 204144 402486 204156
rect 418338 204144 418344 204156
rect 418396 204144 418402 204196
rect 317414 204116 317420 204128
rect 300544 204088 302648 204116
rect 302712 204088 317420 204116
rect 300544 204076 300550 204088
rect 16298 204008 16304 204060
rect 16356 204048 16362 204060
rect 57974 204048 57980 204060
rect 16356 204020 57980 204048
rect 16356 204008 16362 204020
rect 57974 204008 57980 204020
rect 58032 204008 58038 204060
rect 91830 204008 91836 204060
rect 91888 204048 91894 204060
rect 141050 204048 141056 204060
rect 91888 204020 141056 204048
rect 91888 204008 91894 204020
rect 141050 204008 141056 204020
rect 141108 204008 141114 204060
rect 299290 204008 299296 204060
rect 299348 204048 299354 204060
rect 302712 204048 302740 204088
rect 317414 204076 317420 204088
rect 317472 204076 317478 204128
rect 410150 204076 410156 204128
rect 410208 204116 410214 204128
rect 418448 204116 418476 204224
rect 419626 204212 419632 204224
rect 419684 204212 419690 204264
rect 419442 204144 419448 204196
rect 419500 204184 419506 204196
rect 419902 204184 419908 204196
rect 419500 204156 419908 204184
rect 419500 204144 419506 204156
rect 419902 204144 419908 204156
rect 419960 204144 419966 204196
rect 410208 204088 418476 204116
rect 410208 204076 410214 204088
rect 299348 204020 302740 204048
rect 299348 204008 299354 204020
rect 302786 204008 302792 204060
rect 302844 204048 302850 204060
rect 314838 204048 314844 204060
rect 302844 204020 314844 204048
rect 302844 204008 302850 204020
rect 314838 204008 314844 204020
rect 314896 204008 314902 204060
rect 404998 204008 405004 204060
rect 405056 204048 405062 204060
rect 419460 204048 419488 204144
rect 405056 204020 419488 204048
rect 405056 204008 405062 204020
rect 17678 203940 17684 203992
rect 17736 203980 17742 203992
rect 49970 203980 49976 203992
rect 17736 203952 49976 203980
rect 17736 203940 17742 203952
rect 49970 203940 49976 203952
rect 50028 203940 50034 203992
rect 112438 203940 112444 203992
rect 112496 203980 112502 203992
rect 140866 203980 140872 203992
rect 112496 203952 140872 203980
rect 112496 203940 112502 203952
rect 140866 203940 140872 203952
rect 140924 203940 140930 203992
rect 301314 203940 301320 203992
rect 301372 203980 301378 203992
rect 312262 203980 312268 203992
rect 301372 203952 312268 203980
rect 301372 203940 301378 203952
rect 312262 203940 312268 203952
rect 312320 203940 312326 203992
rect 319346 203940 319352 203992
rect 319404 203980 319410 203992
rect 322566 203980 322572 203992
rect 319404 203952 322572 203980
rect 319404 203940 319410 203952
rect 322566 203940 322572 203952
rect 322624 203940 322630 203992
rect 407574 203940 407580 203992
rect 407632 203980 407638 203992
rect 418798 203980 418804 203992
rect 407632 203952 418804 203980
rect 407632 203940 407638 203952
rect 418798 203940 418804 203952
rect 418856 203940 418862 203992
rect 17770 203872 17776 203924
rect 17828 203912 17834 203924
rect 47394 203912 47400 203924
rect 17828 203884 47400 203912
rect 17828 203872 17834 203884
rect 47394 203872 47400 203884
rect 47452 203872 47458 203924
rect 81342 203872 81348 203924
rect 81400 203912 81406 203924
rect 141510 203912 141516 203924
rect 81400 203884 141516 203912
rect 81400 203872 81406 203884
rect 141510 203872 141516 203884
rect 141568 203872 141574 203924
rect 300670 203872 300676 203924
rect 300728 203912 300734 203924
rect 309686 203912 309692 203924
rect 300728 203884 309692 203912
rect 300728 203872 300734 203884
rect 309686 203872 309692 203884
rect 309744 203872 309750 203924
rect 399846 203872 399852 203924
rect 399904 203912 399910 203924
rect 419718 203912 419724 203924
rect 399904 203884 419724 203912
rect 399904 203872 399910 203884
rect 419718 203872 419724 203884
rect 419776 203872 419782 203924
rect 16114 203804 16120 203856
rect 16172 203844 16178 203856
rect 16390 203844 16396 203856
rect 16172 203816 16396 203844
rect 16172 203804 16178 203816
rect 16390 203804 16396 203816
rect 16448 203844 16454 203856
rect 73154 203844 73160 203856
rect 16448 203816 73160 203844
rect 16448 203804 16454 203816
rect 73154 203804 73160 203816
rect 73212 203804 73218 203856
rect 299106 203804 299112 203856
rect 299164 203844 299170 203856
rect 302786 203844 302792 203856
rect 299164 203816 302792 203844
rect 299164 203804 299170 203816
rect 302786 203804 302792 203816
rect 302844 203804 302850 203856
rect 303522 203804 303528 203856
rect 303580 203844 303586 203856
rect 338022 203844 338028 203856
rect 303580 203816 338028 203844
rect 303580 203804 303586 203816
rect 338022 203804 338028 203816
rect 338080 203804 338086 203856
rect 99190 203600 99196 203652
rect 99248 203640 99254 203652
rect 240134 203640 240140 203652
rect 99248 203612 240140 203640
rect 99248 203600 99254 203612
rect 240134 203600 240140 203612
rect 240192 203600 240198 203652
rect 133046 203532 133052 203584
rect 133104 203572 133110 203584
rect 282178 203572 282184 203584
rect 133104 203544 282184 203572
rect 133104 203532 133110 203544
rect 282178 203532 282184 203544
rect 282236 203532 282242 203584
rect 352558 203532 352564 203584
rect 352616 203572 352622 203584
rect 358630 203572 358636 203584
rect 352616 203544 358636 203572
rect 352616 203532 352622 203544
rect 358630 203532 358636 203544
rect 358688 203532 358694 203584
rect 125318 203464 125324 203516
rect 125376 203504 125382 203516
rect 128262 203504 128268 203516
rect 125376 203476 128268 203504
rect 125376 203464 125382 203476
rect 128262 203464 128268 203476
rect 128320 203464 128326 203516
rect 117222 203396 117228 203448
rect 117280 203436 117286 203448
rect 119982 203436 119988 203448
rect 117280 203408 119988 203436
rect 117280 203396 117286 203408
rect 119982 203396 119988 203408
rect 120040 203396 120046 203448
rect 122558 203328 122564 203380
rect 122616 203368 122622 203380
rect 125502 203368 125508 203380
rect 122616 203340 125508 203368
rect 122616 203328 122622 203340
rect 125502 203328 125508 203340
rect 125560 203328 125566 203380
rect 141234 203260 141240 203312
rect 141292 203300 141298 203312
rect 141510 203300 141516 203312
rect 141292 203272 141516 203300
rect 141292 203260 141298 203272
rect 141510 203260 141516 203272
rect 141568 203260 141574 203312
rect 376662 203124 376668 203176
rect 376720 203164 376726 203176
rect 382642 203164 382648 203176
rect 376720 203136 382648 203164
rect 376720 203124 376726 203136
rect 382642 203124 382648 203136
rect 382700 203124 382706 203176
rect 366358 203056 366364 203108
rect 366416 203096 366422 203108
rect 370130 203096 370136 203108
rect 366416 203068 370136 203096
rect 366416 203056 366422 203068
rect 370130 203056 370136 203068
rect 370188 203056 370194 203108
rect 381814 202920 381820 202972
rect 381872 202960 381878 202972
rect 385402 202960 385408 202972
rect 381872 202932 385408 202960
rect 381872 202920 381878 202932
rect 385402 202920 385408 202932
rect 385460 202920 385466 202972
rect 412726 202852 412732 202904
rect 412784 202892 412790 202904
rect 421282 202892 421288 202904
rect 412784 202864 421288 202892
rect 412784 202852 412790 202864
rect 421282 202852 421288 202864
rect 421340 202852 421346 202904
rect 20530 202784 20536 202836
rect 20588 202824 20594 202836
rect 23290 202824 23296 202836
rect 20588 202796 23296 202824
rect 20588 202784 20594 202796
rect 23290 202784 23296 202796
rect 23348 202824 23354 202836
rect 42242 202824 42248 202836
rect 23348 202796 42248 202824
rect 23348 202784 23354 202796
rect 42242 202784 42248 202796
rect 42300 202784 42306 202836
rect 107286 202784 107292 202836
rect 107344 202824 107350 202836
rect 138014 202824 138020 202836
rect 107344 202796 138020 202824
rect 107344 202784 107350 202796
rect 138014 202784 138020 202796
rect 138072 202784 138078 202836
rect 138474 202784 138480 202836
rect 138532 202824 138538 202836
rect 139486 202824 139492 202836
rect 138532 202796 139492 202824
rect 138532 202784 138538 202796
rect 139486 202784 139492 202796
rect 139544 202784 139550 202836
rect 125502 202716 125508 202768
rect 125560 202756 125566 202768
rect 139578 202756 139584 202768
rect 125560 202728 139584 202756
rect 125560 202716 125566 202728
rect 139578 202716 139584 202728
rect 139636 202716 139642 202768
rect 138014 202648 138020 202700
rect 138072 202688 138078 202700
rect 139302 202688 139308 202700
rect 138072 202660 139308 202688
rect 138072 202648 138078 202660
rect 139302 202648 139308 202660
rect 139360 202688 139366 202700
rect 139670 202688 139676 202700
rect 139360 202660 139676 202688
rect 139360 202648 139366 202660
rect 139670 202648 139676 202660
rect 139728 202648 139734 202700
rect 128262 202104 128268 202156
rect 128320 202144 128326 202156
rect 138474 202144 138480 202156
rect 128320 202116 138480 202144
rect 128320 202104 128326 202116
rect 138474 202104 138480 202116
rect 138532 202104 138538 202156
rect 300762 201424 300768 201476
rect 300820 201464 300826 201476
rect 361206 201464 361212 201476
rect 300820 201436 361212 201464
rect 300820 201424 300826 201436
rect 361206 201424 361212 201436
rect 361264 201424 361270 201476
rect 363782 201424 363788 201476
rect 363840 201464 363846 201476
rect 423858 201464 423864 201476
rect 363840 201436 423864 201464
rect 363840 201424 363846 201436
rect 423858 201424 423864 201436
rect 423916 201424 423922 201476
rect 296622 201356 296628 201408
rect 296680 201396 296686 201408
rect 356054 201396 356060 201408
rect 296680 201368 356060 201396
rect 296680 201356 296686 201368
rect 356054 201356 356060 201368
rect 356112 201356 356118 201408
rect 370130 201356 370136 201408
rect 370188 201396 370194 201408
rect 418522 201396 418528 201408
rect 370188 201368 418528 201396
rect 370188 201356 370194 201368
rect 418522 201356 418528 201368
rect 418580 201356 418586 201408
rect 300946 201288 300952 201340
rect 301004 201328 301010 201340
rect 345750 201328 345756 201340
rect 301004 201300 345756 201328
rect 301004 201288 301010 201300
rect 345750 201288 345756 201300
rect 345808 201288 345814 201340
rect 382642 201288 382648 201340
rect 382700 201328 382706 201340
rect 423674 201328 423680 201340
rect 382700 201300 423680 201328
rect 382700 201288 382706 201300
rect 423674 201288 423680 201300
rect 423732 201288 423738 201340
rect 385402 201220 385408 201272
rect 385460 201260 385466 201272
rect 425054 201260 425060 201272
rect 385460 201232 425060 201260
rect 385460 201220 385466 201232
rect 425054 201220 425060 201232
rect 425112 201220 425118 201272
rect 299014 200608 299020 200660
rect 299072 200648 299078 200660
rect 300946 200648 300952 200660
rect 299072 200620 300952 200648
rect 299072 200608 299078 200620
rect 300946 200608 300952 200620
rect 301004 200608 301010 200660
rect 17586 200064 17592 200116
rect 17644 200104 17650 200116
rect 75914 200104 75920 200116
rect 17644 200076 75920 200104
rect 17644 200064 17650 200076
rect 75914 200064 75920 200076
rect 75972 200064 75978 200116
rect 16482 199384 16488 199436
rect 16540 199424 16546 199436
rect 20530 199424 20536 199436
rect 16540 199396 20536 199424
rect 16540 199384 16546 199396
rect 20530 199384 20536 199396
rect 20588 199424 20594 199436
rect 77294 199424 77300 199436
rect 20588 199396 77300 199424
rect 20588 199384 20594 199396
rect 77294 199384 77300 199396
rect 77352 199384 77358 199436
rect 252554 164840 252560 164892
rect 252612 164880 252618 164892
rect 378134 164880 378140 164892
rect 252612 164852 378140 164880
rect 252612 164840 252618 164852
rect 378134 164840 378140 164852
rect 378192 164840 378198 164892
rect 303522 158652 303528 158704
rect 303580 158692 303586 158704
rect 352558 158692 352564 158704
rect 303580 158664 352564 158692
rect 303580 158652 303586 158664
rect 352558 158652 352564 158664
rect 352616 158652 352622 158704
rect 297818 158584 297824 158636
rect 297876 158624 297882 158636
rect 342254 158624 342260 158636
rect 297876 158596 342260 158624
rect 297876 158584 297882 158596
rect 342254 158584 342260 158596
rect 342312 158584 342318 158636
rect 297726 158516 297732 158568
rect 297784 158556 297790 158568
rect 339494 158556 339500 158568
rect 297784 158528 339500 158556
rect 297784 158516 297790 158528
rect 339494 158516 339500 158528
rect 339552 158516 339558 158568
rect 136634 158040 136640 158092
rect 136692 158080 136698 158092
rect 297358 158080 297364 158092
rect 136692 158052 297364 158080
rect 136692 158040 136698 158052
rect 297358 158040 297364 158052
rect 297416 158040 297422 158092
rect 71038 157972 71044 158024
rect 71096 158012 71102 158024
rect 256694 158012 256700 158024
rect 71096 157984 256700 158012
rect 71096 157972 71102 157984
rect 256694 157972 256700 157984
rect 256752 157972 256758 158024
rect 269114 157972 269120 158024
rect 269172 158012 269178 158024
rect 348418 158012 348424 158024
rect 269172 157984 348424 158012
rect 269172 157972 269178 157984
rect 348418 157972 348424 157984
rect 348476 157972 348482 158024
rect 2774 149472 2780 149524
rect 2832 149512 2838 149524
rect 5166 149512 5172 149524
rect 2832 149484 5172 149512
rect 2832 149472 2838 149484
rect 5166 149472 5172 149484
rect 5224 149472 5230 149524
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 13078 136660 13084 136672
rect 3384 136632 13084 136660
rect 3384 136620 3390 136632
rect 13078 136620 13084 136632
rect 13136 136620 13142 136672
rect 135622 78616 135628 78668
rect 135680 78656 135686 78668
rect 138566 78656 138572 78668
rect 135680 78628 138572 78656
rect 135680 78616 135686 78628
rect 138566 78616 138572 78628
rect 138624 78616 138630 78668
rect 300578 78616 300584 78668
rect 300636 78656 300642 78668
rect 306650 78656 306656 78668
rect 300636 78628 306656 78656
rect 300636 78616 300642 78628
rect 306650 78616 306656 78628
rect 306708 78616 306714 78668
rect 410426 78276 410432 78328
rect 410484 78316 410490 78328
rect 419626 78316 419632 78328
rect 410484 78288 419632 78316
rect 410484 78276 410490 78288
rect 419626 78276 419632 78288
rect 419684 78276 419690 78328
rect 407850 78208 407856 78260
rect 407908 78248 407914 78260
rect 418614 78248 418620 78260
rect 407908 78220 418620 78248
rect 407908 78208 407914 78220
rect 418614 78208 418620 78220
rect 418672 78208 418678 78260
rect 405274 78140 405280 78192
rect 405332 78180 405338 78192
rect 419902 78180 419908 78192
rect 405332 78152 419908 78180
rect 405332 78140 405338 78152
rect 419902 78140 419908 78152
rect 419960 78140 419966 78192
rect 297542 78072 297548 78124
rect 297600 78112 297606 78124
rect 327166 78112 327172 78124
rect 297600 78084 327172 78112
rect 297600 78072 297606 78084
rect 327166 78072 327172 78084
rect 327224 78112 327230 78124
rect 327350 78112 327356 78124
rect 327224 78084 327356 78112
rect 327224 78072 327230 78084
rect 327350 78072 327356 78084
rect 327408 78072 327414 78124
rect 398834 78072 398840 78124
rect 398892 78112 398898 78124
rect 400122 78112 400128 78124
rect 398892 78084 400128 78112
rect 398892 78072 398898 78084
rect 400122 78072 400128 78084
rect 400180 78112 400186 78124
rect 419718 78112 419724 78124
rect 400180 78084 419724 78112
rect 400180 78072 400186 78084
rect 419718 78072 419724 78084
rect 419776 78072 419782 78124
rect 300394 78004 300400 78056
rect 300452 78044 300458 78056
rect 330478 78044 330484 78056
rect 300452 78016 330484 78044
rect 300452 78004 300458 78016
rect 330478 78004 330484 78016
rect 330536 78044 330542 78056
rect 332594 78044 332600 78056
rect 330536 78016 332600 78044
rect 330536 78004 330542 78016
rect 332594 78004 332600 78016
rect 332652 78004 332658 78056
rect 396166 78004 396172 78056
rect 396224 78044 396230 78056
rect 397362 78044 397368 78056
rect 396224 78016 397368 78044
rect 396224 78004 396230 78016
rect 397362 78004 397368 78016
rect 397420 78044 397426 78056
rect 419810 78044 419816 78056
rect 397420 78016 419816 78044
rect 397420 78004 397426 78016
rect 419810 78004 419816 78016
rect 419868 78004 419874 78056
rect 130470 77936 130476 77988
rect 130528 77976 130534 77988
rect 139762 77976 139768 77988
rect 130528 77948 139768 77976
rect 130528 77936 130534 77948
rect 139762 77936 139768 77948
rect 139820 77936 139826 77988
rect 269758 77936 269764 77988
rect 269816 77976 269822 77988
rect 369854 77976 369860 77988
rect 269816 77948 369860 77976
rect 269816 77936 269822 77948
rect 369854 77936 369860 77948
rect 369912 77936 369918 77988
rect 393314 77936 393320 77988
rect 393372 77976 393378 77988
rect 422386 77976 422392 77988
rect 393372 77948 422392 77976
rect 393372 77936 393378 77948
rect 422386 77936 422392 77948
rect 422444 77936 422450 77988
rect 68646 77324 68652 77376
rect 68704 77364 68710 77376
rect 70578 77364 70584 77376
rect 68704 77336 70584 77364
rect 68704 77324 68710 77336
rect 70578 77324 70584 77336
rect 70636 77324 70642 77376
rect 348602 77324 348608 77376
rect 348660 77364 348666 77376
rect 350534 77364 350540 77376
rect 348660 77336 350540 77364
rect 348660 77324 348666 77336
rect 350534 77324 350540 77336
rect 350592 77324 350598 77376
rect 77294 77052 77300 77104
rect 77352 77092 77358 77104
rect 78628 77092 78634 77104
rect 77352 77064 78634 77092
rect 77352 77052 77358 77064
rect 78628 77052 78634 77064
rect 78686 77052 78692 77104
rect 390554 76644 390560 76696
rect 390612 76684 390618 76696
rect 421466 76684 421472 76696
rect 390612 76656 421472 76684
rect 390612 76644 390618 76656
rect 421466 76644 421472 76656
rect 421524 76644 421530 76696
rect 301130 76576 301136 76628
rect 301188 76616 301194 76628
rect 329926 76616 329932 76628
rect 301188 76588 329932 76616
rect 301188 76576 301194 76588
rect 329926 76576 329932 76588
rect 329984 76576 329990 76628
rect 378226 76576 378232 76628
rect 378284 76616 378290 76628
rect 421282 76616 421288 76628
rect 378284 76588 421288 76616
rect 378284 76576 378290 76588
rect 421282 76576 421288 76588
rect 421340 76576 421346 76628
rect 299014 76508 299020 76560
rect 299072 76548 299078 76560
rect 336734 76548 336740 76560
rect 299072 76520 336740 76548
rect 299072 76508 299078 76520
rect 336734 76508 336740 76520
rect 336792 76508 336798 76560
rect 376754 76508 376760 76560
rect 376812 76548 376818 76560
rect 422478 76548 422484 76560
rect 376812 76520 422484 76548
rect 376812 76508 376818 76520
rect 422478 76508 422484 76520
rect 422536 76508 422542 76560
rect 20530 75964 20536 76016
rect 20588 76004 20594 76016
rect 77294 76004 77300 76016
rect 20588 75976 77300 76004
rect 20588 75964 20594 75976
rect 77294 75964 77300 75976
rect 77352 75964 77358 76016
rect 17586 75896 17592 75948
rect 17644 75936 17650 75948
rect 75914 75936 75920 75948
rect 17644 75908 75920 75936
rect 17644 75896 17650 75908
rect 75914 75896 75920 75908
rect 75972 75896 75978 75948
rect 304534 75896 304540 75948
rect 304592 75936 304598 75948
rect 580534 75936 580540 75948
rect 304592 75908 580540 75936
rect 304592 75896 304598 75908
rect 580534 75896 580540 75908
rect 580592 75896 580598 75948
rect 18966 75828 18972 75880
rect 19024 75868 19030 75880
rect 34514 75868 34520 75880
rect 19024 75840 34520 75868
rect 19024 75828 19030 75840
rect 34514 75828 34520 75840
rect 34572 75828 34578 75880
rect 91830 75828 91836 75880
rect 91888 75868 91894 75880
rect 140774 75868 140780 75880
rect 91888 75840 140780 75868
rect 91888 75828 91894 75840
rect 140774 75828 140780 75840
rect 140832 75868 140838 75880
rect 141050 75868 141056 75880
rect 140832 75840 141056 75868
rect 140832 75828 140838 75840
rect 141050 75828 141056 75840
rect 141108 75828 141114 75880
rect 333974 75828 333980 75880
rect 334032 75868 334038 75880
rect 334618 75868 334624 75880
rect 334032 75840 334624 75868
rect 334032 75828 334038 75840
rect 334618 75828 334624 75840
rect 334676 75868 334682 75880
rect 338022 75868 338028 75880
rect 334676 75840 338028 75868
rect 334676 75828 334682 75840
rect 338022 75828 338028 75840
rect 338080 75828 338086 75880
rect 345750 75868 345756 75880
rect 344986 75840 345756 75868
rect 17862 75760 17868 75812
rect 17920 75800 17926 75812
rect 63218 75800 63224 75812
rect 17920 75772 63224 75800
rect 17920 75760 17926 75772
rect 63218 75760 63224 75772
rect 63276 75760 63282 75812
rect 107286 75760 107292 75812
rect 107344 75800 107350 75812
rect 139486 75800 139492 75812
rect 107344 75772 139492 75800
rect 107344 75760 107350 75772
rect 139486 75760 139492 75772
rect 139544 75800 139550 75812
rect 139670 75800 139676 75812
rect 139544 75772 139676 75800
rect 139544 75760 139550 75772
rect 139670 75760 139676 75772
rect 139728 75760 139734 75812
rect 322934 75760 322940 75812
rect 322992 75800 322998 75812
rect 325142 75800 325148 75812
rect 322992 75772 325148 75800
rect 322992 75760 322998 75772
rect 325142 75760 325148 75772
rect 325200 75760 325206 75812
rect 327074 75760 327080 75812
rect 327132 75800 327138 75812
rect 330294 75800 330300 75812
rect 327132 75772 330300 75800
rect 327132 75760 327138 75772
rect 330294 75760 330300 75772
rect 330352 75760 330358 75812
rect 336734 75760 336740 75812
rect 336792 75800 336798 75812
rect 344986 75800 345014 75840
rect 345750 75828 345756 75840
rect 345808 75828 345814 75880
rect 363782 75828 363788 75880
rect 363840 75868 363846 75880
rect 423858 75868 423864 75880
rect 363840 75840 423864 75868
rect 363840 75828 363846 75840
rect 423858 75828 423864 75840
rect 423916 75828 423922 75880
rect 336792 75772 345014 75800
rect 336792 75760 336798 75772
rect 386966 75760 386972 75812
rect 387024 75800 387030 75812
rect 421190 75800 421196 75812
rect 387024 75772 421196 75800
rect 387024 75760 387030 75772
rect 421190 75760 421196 75772
rect 421248 75760 421254 75812
rect 16206 75692 16212 75744
rect 16264 75732 16270 75744
rect 60642 75732 60648 75744
rect 16264 75704 60648 75732
rect 16264 75692 16270 75704
rect 60642 75692 60648 75704
rect 60700 75692 60706 75744
rect 112438 75692 112444 75744
rect 112496 75732 112502 75744
rect 140866 75732 140872 75744
rect 112496 75704 140872 75732
rect 112496 75692 112502 75704
rect 140866 75692 140872 75704
rect 140924 75692 140930 75744
rect 329926 75692 329932 75744
rect 329984 75732 329990 75744
rect 335446 75732 335452 75744
rect 329984 75704 335452 75732
rect 329984 75692 329990 75704
rect 335446 75692 335452 75704
rect 335504 75692 335510 75744
rect 384942 75692 384948 75744
rect 385000 75732 385006 75744
rect 418430 75732 418436 75744
rect 385000 75704 418436 75732
rect 385000 75692 385006 75704
rect 418430 75692 418436 75704
rect 418488 75692 418494 75744
rect 16298 75624 16304 75676
rect 16356 75664 16362 75676
rect 57974 75664 57980 75676
rect 16356 75636 57980 75664
rect 16356 75624 16362 75636
rect 57974 75624 57980 75636
rect 58032 75624 58038 75676
rect 122558 75624 122564 75676
rect 122616 75664 122622 75676
rect 139578 75664 139584 75676
rect 122616 75636 139584 75664
rect 122616 75624 122622 75636
rect 139578 75624 139584 75636
rect 139636 75624 139642 75676
rect 389542 75624 389548 75676
rect 389600 75664 389606 75676
rect 422662 75664 422668 75676
rect 389600 75636 422668 75664
rect 389600 75624 389606 75636
rect 422662 75624 422668 75636
rect 422720 75624 422726 75676
rect 17678 75556 17684 75608
rect 17736 75596 17742 75608
rect 50338 75596 50344 75608
rect 17736 75568 50344 75596
rect 17736 75556 17742 75568
rect 50338 75556 50344 75568
rect 50396 75556 50402 75608
rect 125318 75556 125324 75608
rect 125376 75596 125382 75608
rect 138474 75596 138480 75608
rect 125376 75568 138480 75596
rect 125376 75556 125382 75568
rect 138474 75556 138480 75568
rect 138532 75556 138538 75608
rect 300302 75556 300308 75608
rect 300360 75596 300366 75608
rect 322934 75596 322940 75608
rect 300360 75568 322940 75596
rect 300360 75556 300366 75568
rect 322934 75556 322940 75568
rect 322992 75556 322998 75608
rect 17770 75488 17776 75540
rect 17828 75528 17834 75540
rect 47578 75528 47584 75540
rect 17828 75500 47584 75528
rect 17828 75488 17834 75500
rect 47578 75488 47584 75500
rect 47636 75488 47642 75540
rect 119982 75488 119988 75540
rect 120040 75528 120046 75540
rect 131114 75528 131120 75540
rect 120040 75500 131120 75528
rect 120040 75488 120046 75500
rect 131114 75488 131120 75500
rect 131172 75488 131178 75540
rect 298002 75488 298008 75540
rect 298060 75528 298066 75540
rect 327074 75528 327080 75540
rect 298060 75500 327080 75528
rect 298060 75488 298066 75500
rect 327074 75488 327080 75500
rect 327132 75488 327138 75540
rect 16114 75420 16120 75472
rect 16172 75460 16178 75472
rect 73522 75460 73528 75472
rect 16172 75432 73528 75460
rect 16172 75420 16178 75432
rect 73522 75420 73528 75432
rect 73580 75420 73586 75472
rect 127894 75420 127900 75472
rect 127952 75460 127958 75472
rect 138382 75460 138388 75472
rect 127952 75432 138388 75460
rect 127952 75420 127958 75432
rect 138382 75420 138388 75432
rect 138440 75420 138446 75472
rect 297726 75420 297732 75472
rect 297784 75460 297790 75472
rect 332594 75460 332600 75472
rect 297784 75432 332600 75460
rect 297784 75420 297790 75432
rect 332594 75420 332600 75432
rect 332652 75460 332658 75472
rect 340598 75460 340604 75472
rect 332652 75432 340604 75460
rect 332652 75420 332658 75432
rect 340598 75420 340604 75432
rect 340656 75420 340662 75472
rect 57974 75352 57980 75404
rect 58032 75392 58038 75404
rect 59262 75392 59268 75404
rect 58032 75364 59268 75392
rect 58032 75352 58038 75364
rect 59262 75352 59268 75364
rect 59320 75352 59326 75404
rect 140774 75352 140780 75404
rect 140832 75392 140838 75404
rect 210418 75392 210424 75404
rect 140832 75364 210424 75392
rect 140832 75352 140838 75364
rect 210418 75352 210424 75364
rect 210476 75352 210482 75404
rect 280798 75352 280804 75404
rect 280856 75392 280862 75404
rect 379238 75392 379244 75404
rect 280856 75364 379244 75392
rect 280856 75352 280862 75364
rect 379238 75352 379244 75364
rect 379296 75352 379302 75404
rect 379514 75352 379520 75404
rect 379572 75392 379578 75404
rect 412726 75392 412732 75404
rect 379572 75364 412732 75392
rect 379572 75352 379578 75364
rect 412726 75352 412732 75364
rect 412784 75352 412790 75404
rect 133046 75284 133052 75336
rect 133104 75324 133110 75336
rect 231118 75324 231124 75336
rect 133104 75296 231124 75324
rect 133104 75284 133110 75296
rect 231118 75284 231124 75296
rect 231176 75284 231182 75336
rect 273254 75284 273260 75336
rect 273312 75324 273318 75336
rect 384390 75324 384396 75336
rect 273312 75296 384396 75324
rect 273312 75284 273318 75296
rect 384390 75284 384396 75296
rect 384448 75324 384454 75336
rect 384942 75324 384948 75336
rect 384448 75296 384948 75324
rect 384448 75284 384454 75296
rect 384942 75284 384948 75296
rect 385000 75284 385006 75336
rect 71222 75216 71228 75268
rect 71280 75256 71286 75268
rect 77938 75256 77944 75268
rect 71280 75228 77944 75256
rect 71280 75216 71286 75228
rect 77938 75216 77944 75228
rect 77996 75216 78002 75268
rect 140866 75216 140872 75268
rect 140924 75256 140930 75268
rect 254578 75256 254584 75268
rect 140924 75228 254584 75256
rect 140924 75216 140930 75228
rect 254578 75216 254584 75228
rect 254636 75216 254642 75268
rect 277394 75216 277400 75268
rect 277452 75256 277458 75268
rect 389542 75256 389548 75268
rect 277452 75228 389548 75256
rect 277452 75216 277458 75228
rect 389542 75216 389548 75228
rect 389600 75216 389606 75268
rect 34514 75148 34520 75200
rect 34572 75188 34578 75200
rect 100018 75188 100024 75200
rect 34572 75160 100024 75188
rect 34572 75148 34578 75160
rect 100018 75148 100024 75160
rect 100076 75148 100082 75200
rect 139486 75148 139492 75200
rect 139544 75188 139550 75200
rect 285674 75188 285680 75200
rect 139544 75160 285680 75188
rect 139544 75148 139550 75160
rect 285674 75148 285680 75160
rect 285732 75148 285738 75200
rect 297818 75148 297824 75200
rect 297876 75188 297882 75200
rect 335354 75188 335360 75200
rect 297876 75160 335360 75188
rect 297876 75148 297882 75160
rect 335354 75148 335360 75160
rect 335412 75188 335418 75200
rect 343174 75188 343180 75200
rect 335412 75160 343180 75188
rect 335412 75148 335418 75160
rect 343174 75148 343180 75160
rect 343232 75148 343238 75200
rect 351178 75148 351184 75200
rect 351236 75188 351242 75200
rect 386966 75188 386972 75200
rect 351236 75160 386972 75188
rect 351236 75148 351242 75160
rect 386966 75148 386972 75160
rect 387024 75148 387030 75200
rect 396074 75148 396080 75200
rect 396132 75188 396138 75200
rect 417878 75188 417884 75200
rect 396132 75160 417884 75188
rect 396132 75148 396138 75160
rect 417878 75148 417884 75160
rect 417936 75148 417942 75200
rect 21450 74468 21456 74520
rect 21508 74508 21514 74520
rect 27154 74508 27160 74520
rect 21508 74480 27160 74508
rect 21508 74468 21514 74480
rect 27154 74468 27160 74480
rect 27212 74468 27218 74520
rect 300670 74468 300676 74520
rect 300728 74508 300734 74520
rect 309686 74508 309692 74520
rect 300728 74480 309692 74508
rect 300728 74468 300734 74480
rect 309686 74468 309692 74480
rect 309744 74468 309750 74520
rect 368934 74468 368940 74520
rect 368992 74508 368998 74520
rect 419534 74508 419540 74520
rect 368992 74480 419540 74508
rect 368992 74468 368998 74480
rect 419534 74468 419540 74480
rect 419592 74468 419598 74520
rect 16390 74400 16396 74452
rect 16448 74440 16454 74452
rect 44818 74440 44824 74452
rect 16448 74412 44824 74440
rect 16448 74400 16454 74412
rect 44818 74400 44824 74412
rect 44876 74400 44882 74452
rect 298922 74400 298928 74452
rect 298980 74440 298986 74452
rect 319438 74440 319444 74452
rect 298980 74412 319444 74440
rect 298980 74400 298986 74412
rect 319438 74400 319444 74412
rect 319496 74400 319502 74452
rect 376662 74400 376668 74452
rect 376720 74440 376726 74452
rect 423766 74440 423772 74452
rect 376720 74412 423772 74440
rect 376720 74400 376726 74412
rect 423766 74400 423772 74412
rect 423824 74400 423830 74452
rect 18782 74332 18788 74384
rect 18840 74372 18846 74384
rect 37458 74372 37464 74384
rect 18840 74344 37464 74372
rect 18840 74332 18846 74344
rect 37458 74332 37464 74344
rect 37516 74332 37522 74384
rect 299290 74332 299296 74384
rect 299348 74372 299354 74384
rect 318058 74372 318064 74384
rect 299348 74344 318064 74372
rect 299348 74332 299354 74344
rect 318058 74332 318064 74344
rect 318116 74332 318122 74384
rect 381446 74332 381452 74384
rect 381504 74372 381510 74384
rect 425146 74372 425152 74384
rect 381504 74344 425152 74372
rect 381504 74332 381510 74344
rect 425146 74332 425152 74344
rect 425204 74332 425210 74384
rect 19058 74264 19064 74316
rect 19116 74304 19122 74316
rect 32398 74304 32404 74316
rect 19116 74276 32404 74304
rect 19116 74264 19122 74276
rect 32398 74264 32404 74276
rect 32456 74264 32462 74316
rect 299106 74264 299112 74316
rect 299164 74304 299170 74316
rect 315298 74304 315304 74316
rect 299164 74276 315304 74304
rect 299164 74264 299170 74276
rect 315298 74264 315304 74276
rect 315356 74264 315362 74316
rect 392578 74264 392584 74316
rect 392636 74304 392642 74316
rect 424042 74304 424048 74316
rect 392636 74276 424048 74304
rect 392636 74264 392642 74276
rect 424042 74264 424048 74276
rect 424100 74264 424106 74316
rect 18874 74196 18880 74248
rect 18932 74236 18938 74248
rect 29638 74236 29644 74248
rect 18932 74208 29644 74236
rect 18932 74196 18938 74208
rect 29638 74196 29644 74208
rect 29696 74196 29702 74248
rect 301314 74196 301320 74248
rect 301372 74236 301378 74248
rect 312538 74236 312544 74248
rect 301372 74208 312544 74236
rect 301372 74196 301378 74208
rect 312538 74196 312544 74208
rect 312596 74196 312602 74248
rect 394694 74196 394700 74248
rect 394752 74236 394758 74248
rect 425238 74236 425244 74248
rect 394752 74208 425244 74236
rect 394752 74196 394758 74208
rect 425238 74196 425244 74208
rect 425296 74196 425302 74248
rect 21266 74128 21272 74180
rect 21324 74168 21330 74180
rect 55858 74168 55864 74180
rect 21324 74140 55864 74168
rect 21324 74128 21330 74140
rect 55858 74128 55864 74140
rect 55916 74168 55922 74180
rect 56502 74168 56508 74180
rect 55916 74140 56508 74168
rect 55916 74128 55922 74140
rect 56502 74128 56508 74140
rect 56560 74128 56566 74180
rect 299198 74128 299204 74180
rect 299256 74168 299262 74180
rect 322566 74168 322572 74180
rect 299256 74140 322572 74168
rect 299256 74128 299262 74140
rect 322566 74128 322572 74140
rect 322624 74128 322630 74180
rect 402238 74128 402244 74180
rect 402296 74168 402302 74180
rect 418338 74168 418344 74180
rect 402296 74140 418344 74168
rect 402296 74128 402302 74140
rect 418338 74128 418344 74140
rect 418396 74128 418402 74180
rect 415302 74060 415308 74112
rect 415360 74100 415366 74112
rect 421098 74100 421104 74112
rect 415360 74072 421104 74100
rect 415360 74060 415366 74072
rect 421098 74060 421104 74072
rect 421156 74060 421162 74112
rect 138382 73788 138388 73840
rect 138440 73828 138446 73840
rect 308674 73828 308680 73840
rect 138440 73800 308680 73828
rect 138440 73788 138446 73800
rect 308674 73788 308680 73800
rect 308732 73788 308738 73840
rect 394694 73516 394700 73568
rect 394752 73556 394758 73568
rect 395338 73556 395344 73568
rect 394752 73528 395344 73556
rect 394752 73516 394758 73528
rect 395338 73516 395344 73528
rect 395396 73516 395402 73568
rect 309686 73176 309692 73228
rect 309744 73216 309750 73228
rect 311158 73216 311164 73228
rect 309744 73188 311164 73216
rect 309744 73176 309750 73188
rect 311158 73176 311164 73188
rect 311216 73176 311222 73228
rect 321922 73176 321928 73228
rect 321980 73216 321986 73228
rect 322566 73216 322572 73228
rect 321980 73188 322572 73216
rect 321980 73176 321986 73188
rect 322566 73176 322572 73188
rect 322624 73176 322630 73228
rect 376018 73176 376024 73228
rect 376076 73216 376082 73228
rect 376662 73216 376668 73228
rect 376076 73188 376668 73216
rect 376076 73176 376082 73188
rect 376662 73176 376668 73188
rect 376720 73176 376726 73228
rect 414658 73176 414664 73228
rect 414716 73216 414722 73228
rect 415302 73216 415308 73228
rect 414716 73188 415308 73216
rect 414716 73176 414722 73188
rect 415302 73176 415308 73188
rect 415360 73176 415366 73228
rect 104618 73108 104624 73160
rect 104676 73148 104682 73160
rect 138290 73148 138296 73160
rect 104676 73120 138296 73148
rect 104676 73108 104682 73120
rect 138290 73108 138296 73120
rect 138348 73108 138354 73160
rect 138290 72700 138296 72752
rect 138348 72740 138354 72752
rect 283834 72740 283840 72752
rect 138348 72712 283840 72740
rect 138348 72700 138354 72712
rect 283834 72700 283840 72712
rect 283892 72700 283898 72752
rect 75914 72632 75920 72684
rect 75972 72672 75978 72684
rect 224218 72672 224224 72684
rect 75972 72644 224224 72672
rect 75972 72632 75978 72644
rect 224218 72632 224224 72644
rect 224276 72632 224282 72684
rect 300394 72632 300400 72684
rect 300452 72672 300458 72684
rect 409874 72672 409880 72684
rect 300452 72644 409880 72672
rect 300452 72632 300458 72644
rect 409874 72632 409880 72644
rect 409932 72632 409938 72684
rect 212626 72564 212632 72616
rect 212684 72604 212690 72616
rect 363782 72604 363788 72616
rect 212684 72576 363788 72604
rect 212684 72564 212690 72576
rect 363782 72564 363788 72576
rect 363840 72564 363846 72616
rect 139578 72496 139584 72548
rect 139636 72536 139642 72548
rect 305362 72536 305368 72548
rect 139636 72508 305368 72536
rect 139636 72496 139642 72508
rect 305362 72496 305368 72508
rect 305420 72496 305426 72548
rect 59262 72428 59268 72480
rect 59320 72468 59326 72480
rect 357434 72468 357440 72480
rect 59320 72440 357440 72468
rect 59320 72428 59326 72440
rect 357434 72428 357440 72440
rect 357492 72428 357498 72480
rect 270586 71204 270592 71256
rect 270644 71244 270650 71256
rect 348326 71244 348332 71256
rect 270644 71216 348332 71244
rect 270644 71204 270650 71216
rect 348326 71204 348332 71216
rect 348384 71204 348390 71256
rect 137922 71136 137928 71188
rect 137980 71176 137986 71188
rect 381538 71176 381544 71188
rect 137980 71148 381544 71176
rect 137980 71136 137986 71148
rect 381538 71136 381544 71148
rect 381596 71136 381602 71188
rect 37458 71068 37464 71120
rect 37516 71108 37522 71120
rect 345106 71108 345112 71120
rect 37516 71080 345112 71108
rect 37516 71068 37522 71080
rect 345106 71068 345112 71080
rect 345164 71068 345170 71120
rect 27154 71000 27160 71052
rect 27212 71040 27218 71052
rect 338482 71040 338488 71052
rect 27212 71012 338488 71040
rect 27212 71000 27218 71012
rect 338482 71000 338488 71012
rect 338540 71000 338546 71052
rect 3050 70388 3056 70440
rect 3108 70428 3114 70440
rect 199470 70428 199476 70440
rect 3108 70400 199476 70428
rect 3108 70388 3114 70400
rect 199470 70388 199476 70400
rect 199528 70388 199534 70440
rect 81342 70320 81348 70372
rect 81400 70360 81406 70372
rect 141142 70360 141148 70372
rect 81400 70332 141148 70360
rect 81400 70320 81406 70332
rect 141142 70320 141148 70332
rect 141200 70320 141206 70372
rect 141142 69912 141148 69964
rect 141200 69952 141206 69964
rect 227714 69952 227720 69964
rect 141200 69924 227720 69952
rect 141200 69912 141206 69924
rect 227714 69912 227720 69924
rect 227772 69912 227778 69964
rect 73522 69844 73528 69896
rect 73580 69884 73586 69896
rect 222562 69884 222568 69896
rect 73580 69856 222568 69884
rect 73580 69844 73586 69856
rect 222562 69844 222568 69856
rect 222620 69844 222626 69896
rect 298738 69844 298744 69896
rect 298796 69884 298802 69896
rect 407114 69884 407120 69896
rect 298796 69856 407120 69884
rect 298796 69844 298802 69856
rect 407114 69844 407120 69856
rect 407172 69844 407178 69896
rect 215938 69776 215944 69828
rect 215996 69816 216002 69828
rect 368934 69816 368940 69828
rect 215996 69788 368940 69816
rect 215996 69776 216002 69788
rect 368934 69776 368940 69788
rect 368992 69776 368998 69828
rect 139854 69708 139860 69760
rect 139912 69748 139918 69760
rect 303706 69748 303712 69760
rect 139912 69720 303712 69748
rect 139912 69708 139918 69720
rect 303706 69708 303712 69720
rect 303764 69708 303770 69760
rect 60642 69640 60648 69692
rect 60700 69680 60706 69692
rect 360194 69680 360200 69692
rect 60700 69652 360200 69680
rect 60700 69640 60706 69652
rect 360194 69640 360200 69652
rect 360252 69640 360258 69692
rect 84010 68960 84016 69012
rect 84068 69000 84074 69012
rect 142430 69000 142436 69012
rect 84068 68972 142436 69000
rect 84068 68960 84074 68972
rect 142430 68960 142436 68972
rect 142488 69000 142494 69012
rect 143442 69000 143448 69012
rect 142488 68972 143448 69000
rect 142488 68960 142494 68972
rect 143442 68960 143448 68972
rect 143500 68960 143506 69012
rect 117222 68892 117228 68944
rect 117280 68932 117286 68944
rect 139394 68932 139400 68944
rect 117280 68904 139400 68932
rect 117280 68892 117286 68904
rect 139394 68892 139400 68904
rect 139452 68892 139458 68944
rect 143442 68484 143448 68536
rect 143500 68524 143506 68536
rect 229186 68524 229192 68536
rect 143500 68496 229192 68524
rect 143500 68484 143506 68496
rect 229186 68484 229192 68496
rect 229244 68484 229250 68536
rect 229738 68484 229744 68536
rect 229796 68524 229802 68536
rect 368474 68524 368480 68536
rect 229796 68496 368480 68524
rect 229796 68484 229802 68496
rect 368474 68484 368480 68496
rect 368532 68484 368538 68536
rect 138474 68416 138480 68468
rect 138532 68456 138538 68468
rect 290458 68456 290464 68468
rect 138532 68428 290464 68456
rect 138532 68416 138538 68428
rect 290458 68416 290464 68428
rect 290516 68416 290522 68468
rect 297082 68416 297088 68468
rect 297140 68456 297146 68468
rect 404354 68456 404360 68468
rect 297140 68428 404360 68456
rect 297140 68416 297146 68428
rect 404354 68416 404360 68428
rect 404412 68416 404418 68468
rect 139394 68348 139400 68400
rect 139452 68388 139458 68400
rect 302234 68388 302240 68400
rect 139452 68360 302240 68388
rect 139452 68348 139458 68360
rect 302234 68348 302240 68360
rect 302292 68348 302298 68400
rect 63218 68280 63224 68332
rect 63276 68320 63282 68332
rect 361666 68320 361672 68332
rect 63276 68292 361672 68320
rect 63276 68280 63282 68292
rect 361666 68280 361672 68292
rect 361724 68280 361730 68332
rect 77938 66988 77944 67040
rect 77996 67028 78002 67040
rect 255682 67028 255688 67040
rect 77996 67000 255688 67028
rect 77996 66988 78002 67000
rect 255682 66988 255688 67000
rect 255740 66988 255746 67040
rect 292114 66988 292120 67040
rect 292172 67028 292178 67040
rect 396166 67028 396172 67040
rect 292172 67000 396172 67028
rect 292172 66988 292178 67000
rect 396166 66988 396172 67000
rect 396224 66988 396230 67040
rect 56502 66920 56508 66972
rect 56560 66960 56566 66972
rect 356698 66960 356704 66972
rect 56560 66932 356704 66960
rect 56560 66920 56566 66932
rect 356698 66920 356704 66932
rect 356756 66920 356762 66972
rect 42058 66852 42064 66904
rect 42116 66892 42122 66904
rect 348418 66892 348424 66904
rect 42116 66864 348424 66892
rect 42116 66852 42122 66864
rect 348418 66852 348424 66864
rect 348476 66852 348482 66904
rect 88334 66172 88340 66224
rect 88392 66212 88398 66224
rect 143626 66212 143632 66224
rect 88392 66184 143632 66212
rect 88392 66172 88398 66184
rect 143626 66172 143632 66184
rect 143684 66212 143690 66224
rect 144822 66212 144828 66224
rect 143684 66184 144828 66212
rect 143684 66172 143690 66184
rect 144822 66172 144828 66184
rect 144880 66172 144886 66224
rect 295334 66172 295340 66224
rect 295392 66212 295398 66224
rect 296622 66212 296628 66224
rect 295392 66184 296628 66212
rect 295392 66172 295398 66184
rect 296622 66172 296628 66184
rect 296680 66212 296686 66224
rect 356054 66212 356060 66224
rect 296680 66184 356060 66212
rect 296680 66172 296686 66184
rect 356054 66172 356060 66184
rect 356112 66172 356118 66224
rect 93854 66104 93860 66156
rect 93912 66144 93918 66156
rect 142338 66144 142344 66156
rect 93912 66116 142344 66144
rect 93912 66104 93918 66116
rect 142338 66104 142344 66116
rect 142396 66144 142402 66156
rect 143442 66144 143448 66156
rect 142396 66116 143448 66144
rect 142396 66104 142402 66116
rect 143442 66104 143448 66116
rect 143500 66104 143506 66156
rect 96614 66036 96620 66088
rect 96672 66076 96678 66088
rect 140774 66076 140780 66088
rect 96672 66048 140780 66076
rect 96672 66036 96678 66048
rect 140774 66036 140780 66048
rect 140832 66076 140838 66088
rect 141050 66076 141056 66088
rect 140832 66048 141056 66076
rect 140832 66036 140838 66048
rect 141050 66036 141056 66048
rect 141108 66036 141114 66088
rect 144822 65696 144828 65748
rect 144880 65736 144886 65748
rect 232498 65736 232504 65748
rect 144880 65708 232504 65736
rect 144880 65696 144886 65708
rect 232498 65696 232504 65708
rect 232556 65696 232562 65748
rect 207658 65628 207664 65680
rect 207716 65668 207722 65680
rect 295334 65668 295340 65680
rect 207716 65640 295340 65668
rect 207716 65628 207722 65640
rect 295334 65628 295340 65640
rect 295392 65628 295398 65680
rect 143442 65560 143448 65612
rect 143500 65600 143506 65612
rect 235994 65600 236000 65612
rect 143500 65572 236000 65600
rect 143500 65560 143506 65572
rect 235994 65560 236000 65572
rect 236052 65560 236058 65612
rect 254026 65560 254032 65612
rect 254084 65600 254090 65612
rect 280798 65600 280804 65612
rect 254084 65572 280804 65600
rect 254084 65560 254090 65572
rect 280798 65560 280804 65572
rect 280856 65560 280862 65612
rect 293954 65560 293960 65612
rect 294012 65600 294018 65612
rect 398834 65600 398840 65612
rect 294012 65572 398840 65600
rect 294012 65560 294018 65572
rect 398834 65560 398840 65572
rect 398892 65560 398898 65612
rect 140774 65492 140780 65544
rect 140832 65532 140838 65544
rect 237466 65532 237472 65544
rect 140832 65504 237472 65532
rect 140832 65492 140838 65504
rect 237466 65492 237472 65504
rect 237524 65492 237530 65544
rect 272242 65492 272248 65544
rect 272300 65532 272306 65544
rect 381446 65532 381452 65544
rect 272300 65504 381452 65532
rect 272300 65492 272306 65504
rect 381446 65492 381452 65504
rect 381504 65492 381510 65544
rect 214282 64336 214288 64388
rect 214340 64376 214346 64388
rect 366358 64376 366364 64388
rect 214340 64348 366364 64376
rect 214340 64336 214346 64348
rect 366358 64336 366364 64348
rect 366416 64336 366422 64388
rect 50338 64268 50344 64320
rect 50396 64308 50402 64320
rect 353386 64308 353392 64320
rect 50396 64280 353392 64308
rect 50396 64268 50402 64280
rect 353386 64268 353392 64280
rect 353444 64268 353450 64320
rect 47578 64200 47584 64252
rect 47636 64240 47642 64252
rect 351914 64240 351920 64252
rect 47636 64212 351920 64240
rect 47636 64200 47642 64212
rect 351914 64200 351920 64212
rect 351972 64200 351978 64252
rect 44818 64132 44824 64184
rect 44876 64172 44882 64184
rect 350074 64172 350080 64184
rect 44876 64144 350080 64172
rect 44876 64132 44882 64144
rect 350074 64132 350080 64144
rect 350132 64132 350138 64184
rect 300762 63452 300768 63504
rect 300820 63492 300826 63504
rect 360286 63492 360292 63504
rect 300820 63464 360292 63492
rect 300820 63452 300826 63464
rect 360286 63452 360292 63464
rect 360344 63452 360350 63504
rect 211154 62976 211160 63028
rect 211212 63016 211218 63028
rect 300762 63016 300768 63028
rect 211212 62988 300768 63016
rect 211212 62976 211218 62988
rect 300762 62976 300768 62988
rect 300820 62976 300826 63028
rect 65518 62908 65524 62960
rect 65576 62948 65582 62960
rect 322934 62948 322940 62960
rect 65576 62920 322940 62948
rect 65576 62908 65582 62920
rect 322934 62908 322940 62920
rect 322992 62908 322998 62960
rect 32398 62840 32404 62892
rect 32456 62880 32462 62892
rect 341794 62880 341800 62892
rect 32456 62852 341800 62880
rect 32456 62840 32462 62852
rect 341794 62840 341800 62852
rect 341852 62840 341858 62892
rect 29638 62772 29644 62824
rect 29696 62812 29702 62824
rect 340138 62812 340144 62824
rect 29696 62784 340144 62812
rect 29696 62772 29702 62784
rect 340138 62772 340144 62784
rect 340196 62772 340202 62824
rect 340230 62772 340236 62824
rect 340288 62812 340294 62824
rect 392578 62812 392584 62824
rect 340288 62784 392584 62812
rect 340288 62772 340294 62784
rect 392578 62772 392584 62784
rect 392636 62772 392642 62824
rect 13078 62024 13084 62076
rect 13136 62064 13142 62076
rect 57054 62064 57060 62076
rect 13136 62036 57060 62064
rect 13136 62024 13142 62036
rect 57054 62024 57060 62036
rect 57112 62024 57118 62076
rect 100754 62024 100760 62076
rect 100812 62064 100818 62076
rect 140774 62064 140780 62076
rect 100812 62036 140780 62064
rect 100812 62024 100818 62036
rect 140774 62024 140780 62036
rect 140832 62024 140838 62076
rect 301406 62024 301412 62076
rect 301464 62064 301470 62076
rect 371326 62064 371332 62076
rect 301464 62036 371332 62064
rect 301464 62024 301470 62036
rect 371326 62024 371332 62036
rect 371384 62024 371390 62076
rect 98362 61684 98368 61736
rect 98420 61724 98426 61736
rect 239122 61724 239128 61736
rect 98420 61696 239128 61724
rect 98420 61684 98426 61696
rect 239122 61684 239128 61696
rect 239180 61684 239186 61736
rect 217594 61548 217600 61600
rect 217652 61588 217658 61600
rect 301406 61588 301412 61600
rect 217652 61560 301412 61588
rect 217652 61548 217658 61560
rect 301406 61548 301412 61560
rect 301464 61548 301470 61600
rect 280522 61480 280528 61532
rect 280580 61520 280586 61532
rect 395338 61520 395344 61532
rect 280580 61492 395344 61520
rect 280580 61480 280586 61492
rect 395338 61480 395344 61492
rect 395396 61480 395402 61532
rect 140774 61412 140780 61464
rect 140832 61452 140838 61464
rect 141418 61452 141424 61464
rect 140832 61424 141424 61452
rect 140832 61412 140838 61424
rect 141418 61412 141424 61424
rect 141476 61452 141482 61464
rect 282086 61452 282092 61464
rect 141476 61424 282092 61452
rect 141476 61412 141482 61424
rect 282086 61412 282092 61424
rect 282144 61412 282150 61464
rect 282178 61412 282184 61464
rect 282236 61452 282242 61464
rect 366634 61452 366640 61464
rect 282236 61424 366640 61452
rect 282236 61412 282242 61424
rect 366634 61412 366640 61424
rect 366692 61412 366698 61464
rect 220906 61344 220912 61396
rect 220964 61384 220970 61396
rect 376018 61384 376024 61396
rect 220964 61356 376024 61384
rect 220964 61344 220970 61356
rect 376018 61344 376024 61356
rect 376076 61344 376082 61396
rect 294046 60664 294052 60716
rect 294104 60704 294110 60716
rect 295242 60704 295248 60716
rect 294104 60676 295248 60704
rect 294104 60664 294110 60676
rect 295242 60664 295248 60676
rect 295300 60704 295306 60716
rect 353294 60704 353300 60716
rect 295300 60676 353300 60704
rect 295300 60664 295306 60676
rect 353294 60664 353300 60676
rect 353352 60664 353358 60716
rect 302326 60596 302332 60648
rect 302384 60636 302390 60648
rect 357526 60636 357532 60648
rect 302384 60608 357532 60636
rect 302384 60596 302390 60608
rect 357526 60596 357532 60608
rect 357584 60596 357590 60648
rect 206002 60120 206008 60172
rect 206060 60160 206066 60172
rect 294046 60160 294052 60172
rect 206060 60132 294052 60160
rect 206060 60120 206066 60132
rect 294046 60120 294052 60132
rect 294104 60120 294110 60172
rect 231118 60052 231124 60104
rect 231176 60092 231182 60104
rect 364978 60092 364984 60104
rect 231176 60064 364984 60092
rect 231176 60052 231182 60064
rect 364978 60052 364984 60064
rect 365036 60052 365042 60104
rect 219434 59984 219440 60036
rect 219492 60024 219498 60036
rect 374638 60024 374644 60036
rect 219492 59996 374644 60024
rect 219492 59984 219498 59996
rect 374638 59984 374644 59996
rect 374696 59984 374702 60036
rect 209314 59372 209320 59424
rect 209372 59412 209378 59424
rect 302326 59412 302332 59424
rect 209372 59384 302332 59412
rect 209372 59372 209378 59384
rect 302326 59372 302332 59384
rect 302384 59372 302390 59424
rect 135254 58828 135260 58880
rect 135312 58868 135318 58880
rect 204346 58868 204352 58880
rect 135312 58840 204352 58868
rect 135312 58828 135318 58840
rect 204346 58828 204352 58840
rect 204404 58828 204410 58880
rect 210418 58828 210424 58880
rect 210476 58868 210482 58880
rect 234154 58868 234160 58880
rect 210476 58840 234160 58868
rect 210476 58828 210482 58840
rect 234154 58828 234160 58840
rect 234212 58828 234218 58880
rect 254578 58828 254584 58880
rect 254636 58868 254642 58880
rect 288802 58868 288808 58880
rect 254636 58840 288808 58868
rect 254636 58828 254642 58840
rect 288802 58828 288808 58840
rect 288860 58828 288866 58880
rect 295426 58828 295432 58880
rect 295484 58868 295490 58880
rect 402238 58868 402244 58880
rect 295484 58840 402244 58868
rect 295484 58828 295490 58840
rect 402238 58828 402244 58840
rect 402296 58828 402302 58880
rect 129734 58760 129740 58812
rect 129792 58800 129798 58812
rect 307110 58800 307116 58812
rect 129792 58772 307116 58800
rect 129792 58760 129798 58772
rect 307110 58760 307116 58772
rect 307168 58760 307174 58812
rect 202874 58692 202880 58744
rect 202932 58732 202938 58744
rect 414658 58732 414664 58744
rect 202932 58704 414664 58732
rect 202932 58692 202938 58704
rect 414658 58692 414664 58704
rect 414716 58692 414722 58744
rect 100018 58624 100024 58676
rect 100076 58664 100082 58676
rect 343634 58664 343640 58676
rect 100076 58636 343640 58664
rect 100076 58624 100082 58636
rect 343634 58624 343640 58636
rect 343692 58624 343698 58676
rect 109034 57876 109040 57928
rect 109092 57916 109098 57928
rect 142246 57916 142252 57928
rect 109092 57888 142252 57916
rect 109092 57876 109098 57888
rect 142246 57876 142252 57888
rect 142304 57916 142310 57928
rect 143442 57916 143448 57928
rect 142304 57888 143448 57916
rect 142304 57876 142310 57888
rect 143442 57876 143448 57888
rect 143500 57876 143506 57928
rect 311158 57876 311164 57928
rect 311216 57916 311222 57928
rect 314010 57916 314016 57928
rect 311216 57888 314016 57916
rect 311216 57876 311222 57888
rect 314010 57876 314016 57888
rect 314068 57876 314074 57928
rect 318058 57876 318064 57928
rect 318116 57916 318122 57928
rect 318978 57916 318984 57928
rect 318116 57888 318984 57916
rect 318116 57876 318122 57888
rect 318978 57876 318984 57888
rect 319036 57876 319042 57928
rect 319438 57876 319444 57928
rect 319496 57916 319502 57928
rect 320634 57916 320640 57928
rect 319496 57888 320640 57916
rect 319496 57876 319502 57888
rect 320634 57876 320640 57888
rect 320692 57876 320698 57928
rect 328914 57876 328920 57928
rect 328972 57916 328978 57928
rect 330478 57916 330484 57928
rect 328972 57888 330484 57916
rect 328972 57876 328978 57888
rect 330478 57876 330484 57888
rect 330536 57876 330542 57928
rect 114554 57808 114560 57860
rect 114612 57848 114618 57860
rect 142154 57848 142160 57860
rect 114612 57820 142160 57848
rect 114612 57808 114618 57820
rect 142154 57808 142160 57820
rect 142212 57848 142218 57860
rect 143350 57848 143356 57860
rect 142212 57820 143356 57848
rect 142212 57808 142218 57820
rect 143350 57808 143356 57820
rect 143408 57808 143414 57860
rect 306374 57808 306380 57860
rect 306432 57848 306438 57860
rect 312354 57848 312360 57860
rect 306432 57820 312360 57848
rect 306432 57808 306438 57820
rect 312354 57808 312360 57820
rect 312412 57808 312418 57860
rect 312538 57808 312544 57860
rect 312596 57848 312602 57860
rect 315666 57848 315672 57860
rect 312596 57820 315672 57848
rect 312596 57808 312602 57820
rect 315666 57808 315672 57820
rect 315724 57808 315730 57860
rect 332226 57740 332232 57792
rect 332284 57780 332290 57792
rect 334618 57780 334624 57792
rect 332284 57752 334624 57780
rect 332284 57740 332290 57752
rect 334618 57740 334624 57752
rect 334676 57740 334682 57792
rect 307386 57644 307392 57656
rect 296686 57616 307392 57644
rect 290458 57536 290464 57588
rect 290516 57576 290522 57588
rect 296686 57576 296714 57616
rect 307386 57604 307392 57616
rect 307444 57604 307450 57656
rect 290516 57548 296714 57576
rect 290516 57536 290522 57548
rect 322934 57536 322940 57588
rect 322992 57576 322998 57588
rect 363690 57576 363696 57588
rect 322992 57548 363696 57576
rect 322992 57536 322998 57548
rect 363690 57536 363696 57548
rect 363748 57536 363754 57588
rect 279234 57468 279240 57520
rect 279292 57508 279298 57520
rect 340230 57508 340236 57520
rect 279292 57480 340236 57508
rect 279292 57468 279298 57480
rect 340230 57468 340236 57480
rect 340288 57468 340294 57520
rect 275922 57400 275928 57452
rect 275980 57440 275986 57452
rect 351178 57440 351184 57452
rect 275980 57412 351184 57440
rect 275980 57400 275986 57412
rect 351178 57400 351184 57412
rect 351236 57400 351242 57452
rect 297358 57332 297364 57384
rect 297416 57372 297422 57384
rect 383562 57372 383568 57384
rect 297416 57344 383568 57372
rect 297416 57332 297422 57344
rect 383562 57332 383568 57344
rect 383620 57332 383626 57384
rect 143442 57264 143448 57316
rect 143500 57304 143506 57316
rect 287514 57304 287520 57316
rect 143500 57276 287520 57304
rect 143500 57264 143506 57276
rect 287514 57264 287520 57276
rect 287572 57264 287578 57316
rect 296070 57264 296076 57316
rect 296128 57304 296134 57316
rect 385218 57304 385224 57316
rect 296128 57276 385224 57304
rect 296128 57264 296134 57276
rect 385218 57264 385224 57276
rect 385276 57264 385282 57316
rect 395154 57264 395160 57316
rect 395212 57304 395218 57316
rect 418246 57304 418252 57316
rect 395212 57276 418252 57304
rect 395212 57264 395218 57276
rect 418246 57264 418252 57276
rect 418304 57264 418310 57316
rect 143350 57196 143356 57248
rect 143408 57236 143414 57248
rect 290826 57236 290832 57248
rect 143408 57208 290832 57236
rect 143408 57196 143414 57208
rect 290826 57196 290832 57208
rect 290884 57196 290890 57248
rect 295978 57196 295984 57248
rect 296036 57236 296042 57248
rect 388530 57236 388536 57248
rect 296036 57208 388536 57236
rect 296036 57196 296042 57208
rect 388530 57196 388536 57208
rect 388588 57196 388594 57248
rect 390186 57196 390192 57248
rect 390244 57236 390250 57248
rect 422294 57236 422300 57248
rect 390244 57208 422300 57236
rect 390244 57196 390250 57208
rect 422294 57196 422300 57208
rect 422352 57196 422358 57248
rect 307110 56924 307116 56976
rect 307168 56964 307174 56976
rect 310698 56964 310704 56976
rect 307168 56936 310704 56964
rect 307168 56924 307174 56936
rect 310698 56924 310704 56936
rect 310756 56924 310762 56976
rect 315298 56584 315304 56636
rect 315356 56624 315362 56636
rect 317322 56624 317328 56636
rect 315356 56596 317328 56624
rect 315356 56584 315362 56596
rect 317322 56584 317328 56596
rect 317380 56584 317386 56636
rect 325602 56584 325608 56636
rect 325660 56624 325666 56636
rect 327166 56624 327172 56636
rect 325660 56596 327172 56624
rect 325660 56584 325666 56596
rect 327166 56584 327172 56596
rect 327224 56584 327230 56636
rect 5166 56516 5172 56568
rect 5224 56556 5230 56568
rect 57514 56556 57520 56568
rect 5224 56528 57520 56556
rect 5224 56516 5230 56528
rect 57514 56516 57520 56528
rect 57572 56516 57578 56568
rect 102134 55224 102140 55276
rect 102192 55264 102198 55276
rect 196618 55264 196624 55276
rect 102192 55236 196624 55264
rect 102192 55224 102198 55236
rect 196618 55224 196624 55236
rect 196676 55224 196682 55276
rect 102134 53864 102140 53916
rect 102192 53904 102198 53916
rect 103882 53904 103888 53916
rect 102192 53876 103888 53904
rect 102192 53864 102198 53876
rect 103882 53864 103888 53876
rect 103940 53864 103946 53916
rect 399478 53048 399484 53100
rect 399536 53088 399542 53100
rect 580258 53088 580264 53100
rect 399536 53060 580264 53088
rect 399536 53048 399542 53060
rect 580258 53048 580264 53060
rect 580316 53048 580322 53100
rect 102134 52504 102140 52556
rect 102192 52544 102198 52556
rect 196158 52544 196164 52556
rect 102192 52516 196164 52544
rect 102192 52504 102198 52516
rect 196158 52504 196164 52516
rect 196216 52504 196222 52556
rect 102226 52436 102232 52488
rect 102284 52476 102290 52488
rect 103974 52476 103980 52488
rect 102284 52448 103980 52476
rect 102284 52436 102290 52448
rect 103974 52436 103980 52448
rect 104032 52436 104038 52488
rect 5074 52368 5080 52420
rect 5132 52408 5138 52420
rect 57054 52408 57060 52420
rect 5132 52380 57060 52408
rect 5132 52368 5138 52380
rect 57054 52368 57060 52380
rect 57112 52368 57118 52420
rect 102870 52368 102876 52420
rect 102928 52408 102934 52420
rect 195974 52408 195980 52420
rect 102928 52380 195980 52408
rect 102928 52368 102934 52380
rect 195974 52368 195980 52380
rect 196032 52368 196038 52420
rect 103146 52300 103152 52352
rect 103204 52340 103210 52352
rect 196066 52340 196072 52352
rect 103204 52312 196072 52340
rect 103204 52300 103210 52312
rect 196066 52300 196072 52312
rect 196124 52300 196130 52352
rect 103054 51008 103060 51060
rect 103112 51048 103118 51060
rect 195974 51048 195980 51060
rect 103112 51020 195980 51048
rect 103112 51008 103118 51020
rect 195974 51008 195980 51020
rect 196032 51008 196038 51060
rect 102134 49784 102140 49836
rect 102192 49824 102198 49836
rect 104342 49824 104348 49836
rect 102192 49796 104348 49824
rect 102192 49784 102198 49796
rect 104342 49784 104348 49796
rect 104400 49784 104406 49836
rect 102778 49648 102784 49700
rect 102836 49688 102842 49700
rect 195974 49688 195980 49700
rect 102836 49660 195980 49688
rect 102836 49648 102842 49660
rect 195974 49648 195980 49660
rect 196032 49648 196038 49700
rect 102594 49580 102600 49632
rect 102652 49620 102658 49632
rect 196066 49620 196072 49632
rect 102652 49592 196072 49620
rect 102652 49580 102658 49592
rect 196066 49580 196072 49592
rect 196124 49580 196130 49632
rect 103882 48220 103888 48272
rect 103940 48260 103946 48272
rect 195974 48260 195980 48272
rect 103940 48232 195980 48260
rect 103940 48220 103946 48232
rect 195974 48220 195980 48232
rect 196032 48220 196038 48272
rect 6178 46860 6184 46912
rect 6236 46900 6242 46912
rect 57514 46900 57520 46912
rect 6236 46872 57520 46900
rect 6236 46860 6242 46872
rect 57514 46860 57520 46872
rect 57572 46860 57578 46912
rect 103974 46860 103980 46912
rect 104032 46900 104038 46912
rect 195974 46900 195980 46912
rect 104032 46872 195980 46900
rect 104032 46860 104038 46872
rect 195974 46860 195980 46872
rect 196032 46860 196038 46912
rect 103238 45500 103244 45552
rect 103296 45540 103302 45552
rect 195974 45540 195980 45552
rect 103296 45512 195980 45540
rect 103296 45500 103302 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 3326 44140 3332 44192
rect 3384 44180 3390 44192
rect 59998 44180 60004 44192
rect 3384 44152 60004 44180
rect 3384 44140 3390 44152
rect 59998 44140 60004 44152
rect 60056 44140 60062 44192
rect 102870 44072 102876 44124
rect 102928 44112 102934 44124
rect 196066 44112 196072 44124
rect 102928 44084 196072 44112
rect 102928 44072 102934 44084
rect 196066 44072 196072 44084
rect 196124 44072 196130 44124
rect 104342 44004 104348 44056
rect 104400 44044 104406 44056
rect 195974 44044 195980 44056
rect 104400 44016 195980 44044
rect 104400 44004 104406 44016
rect 195974 44004 195980 44016
rect 196032 44004 196038 44056
rect 3510 42712 3516 42764
rect 3568 42752 3574 42764
rect 57146 42752 57152 42764
rect 3568 42724 57152 42752
rect 3568 42712 3574 42724
rect 57146 42712 57152 42724
rect 57204 42712 57210 42764
rect 102594 42712 102600 42764
rect 102652 42752 102658 42764
rect 196066 42752 196072 42764
rect 102652 42724 196072 42752
rect 102652 42712 102658 42724
rect 196066 42712 196072 42724
rect 196124 42712 196130 42764
rect 102962 42644 102968 42696
rect 103020 42684 103026 42696
rect 195974 42684 195980 42696
rect 103020 42656 195980 42684
rect 103020 42644 103026 42656
rect 195974 42644 195980 42656
rect 196032 42644 196038 42696
rect 103514 41352 103520 41404
rect 103572 41392 103578 41404
rect 195974 41392 195980 41404
rect 103572 41364 195980 41392
rect 103572 41352 103578 41364
rect 195974 41352 195980 41364
rect 196032 41352 196038 41404
rect 102134 40672 102140 40724
rect 102192 40712 102198 40724
rect 196158 40712 196164 40724
rect 102192 40684 196164 40712
rect 102192 40672 102198 40684
rect 196158 40672 196164 40684
rect 196216 40672 196222 40724
rect 102318 39992 102324 40044
rect 102376 40032 102382 40044
rect 196066 40032 196072 40044
rect 102376 40004 196072 40032
rect 102376 39992 102382 40004
rect 196066 39992 196072 40004
rect 196124 39992 196130 40044
rect 103606 39924 103612 39976
rect 103664 39964 103670 39976
rect 195974 39964 195980 39976
rect 103664 39936 195980 39964
rect 103664 39924 103670 39936
rect 195974 39924 195980 39936
rect 196032 39924 196038 39976
rect 102226 38564 102232 38616
rect 102284 38604 102290 38616
rect 195974 38604 195980 38616
rect 102284 38576 195980 38604
rect 102284 38564 102290 38576
rect 195974 38564 195980 38576
rect 196032 38564 196038 38616
rect 6270 37204 6276 37256
rect 6328 37244 6334 37256
rect 57054 37244 57060 37256
rect 6328 37216 57060 37244
rect 6328 37204 6334 37216
rect 57054 37204 57060 37216
rect 57112 37204 57118 37256
rect 102134 37204 102140 37256
rect 102192 37244 102198 37256
rect 195974 37244 195980 37256
rect 102192 37216 195980 37244
rect 102192 37204 102198 37216
rect 195974 37204 195980 37216
rect 196032 37204 196038 37256
rect 102778 35844 102784 35896
rect 102836 35884 102842 35896
rect 195974 35884 195980 35896
rect 102836 35856 195980 35884
rect 102836 35844 102842 35856
rect 195974 35844 195980 35856
rect 196032 35844 196038 35896
rect 102594 35776 102600 35828
rect 102652 35816 102658 35828
rect 196066 35816 196072 35828
rect 102652 35788 196072 35816
rect 102652 35776 102658 35788
rect 196066 35776 196072 35788
rect 196124 35776 196130 35828
rect 102686 34416 102692 34468
rect 102744 34456 102750 34468
rect 196066 34456 196072 34468
rect 102744 34428 196072 34456
rect 102744 34416 102750 34428
rect 196066 34416 196072 34428
rect 196124 34416 196130 34468
rect 102870 34348 102876 34400
rect 102928 34388 102934 34400
rect 195974 34388 195980 34400
rect 102928 34360 195980 34388
rect 102928 34348 102934 34360
rect 195974 34348 195980 34360
rect 196032 34348 196038 34400
rect 102134 33056 102140 33108
rect 102192 33096 102198 33108
rect 195974 33096 195980 33108
rect 102192 33068 195980 33096
rect 102192 33056 102198 33068
rect 195974 33056 195980 33068
rect 196032 33056 196038 33108
rect 4890 31696 4896 31748
rect 4948 31736 4954 31748
rect 57606 31736 57612 31748
rect 4948 31708 57612 31736
rect 4948 31696 4954 31708
rect 57606 31696 57612 31708
rect 57664 31696 57670 31748
rect 102134 31696 102140 31748
rect 102192 31736 102198 31748
rect 196066 31736 196072 31748
rect 102192 31708 196072 31736
rect 102192 31696 102198 31708
rect 196066 31696 196072 31708
rect 196124 31696 196130 31748
rect 102318 31628 102324 31680
rect 102376 31668 102382 31680
rect 195974 31668 195980 31680
rect 102376 31640 195980 31668
rect 102376 31628 102382 31640
rect 195974 31628 195980 31640
rect 196032 31628 196038 31680
rect 102134 30268 102140 30320
rect 102192 30308 102198 30320
rect 196066 30308 196072 30320
rect 102192 30280 196072 30308
rect 102192 30268 102198 30280
rect 196066 30268 196072 30280
rect 196124 30268 196130 30320
rect 102226 30200 102232 30252
rect 102284 30240 102290 30252
rect 195974 30240 195980 30252
rect 102284 30212 195980 30240
rect 102284 30200 102290 30212
rect 195974 30200 195980 30212
rect 196032 30200 196038 30252
rect 102134 28908 102140 28960
rect 102192 28948 102198 28960
rect 195974 28948 195980 28960
rect 102192 28920 195980 28948
rect 102192 28908 102198 28920
rect 195974 28908 195980 28920
rect 196032 28908 196038 28960
rect 102134 28228 102140 28280
rect 102192 28268 102198 28280
rect 195974 28268 195980 28280
rect 102192 28240 195980 28268
rect 102192 28228 102198 28240
rect 195974 28228 195980 28240
rect 196032 28228 196038 28280
rect 17218 27548 17224 27600
rect 17276 27588 17282 27600
rect 57238 27588 57244 27600
rect 17276 27560 57244 27588
rect 17276 27548 17282 27560
rect 57238 27548 57244 27560
rect 57296 27548 57302 27600
rect 102134 27548 102140 27600
rect 102192 27588 102198 27600
rect 195974 27588 195980 27600
rect 102192 27560 195980 27588
rect 102192 27548 102198 27560
rect 195974 27548 195980 27560
rect 196032 27548 196038 27600
rect 102778 26188 102784 26240
rect 102836 26228 102842 26240
rect 195974 26228 195980 26240
rect 102836 26200 195980 26228
rect 102836 26188 102842 26200
rect 195974 26188 195980 26200
rect 196032 26188 196038 26240
rect 397178 24624 397184 24676
rect 397236 24664 397242 24676
rect 399478 24664 399484 24676
rect 397236 24636 399484 24664
rect 397236 24624 397242 24636
rect 399478 24624 399484 24636
rect 399536 24624 399542 24676
rect 20622 24216 20628 24268
rect 20680 24256 20686 24268
rect 356974 24256 356980 24268
rect 20680 24228 356980 24256
rect 20680 24216 20686 24228
rect 356974 24216 356980 24228
rect 357032 24216 357038 24268
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 360654 24188 360660 24200
rect 20128 24160 360660 24188
rect 20128 24148 20134 24160
rect 360654 24148 360660 24160
rect 360712 24148 360718 24200
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 371326 24120 371332 24132
rect 3476 24092 371332 24120
rect 3476 24080 3482 24092
rect 371326 24080 371332 24092
rect 371384 24080 371390 24132
rect 85482 23468 85488 23520
rect 85540 23508 85546 23520
rect 266354 23508 266360 23520
rect 85540 23480 266360 23508
rect 85540 23468 85546 23480
rect 266354 23468 266360 23480
rect 266412 23508 266418 23520
rect 267366 23508 267372 23520
rect 266412 23480 267372 23508
rect 266412 23468 266418 23480
rect 267366 23468 267372 23480
rect 267424 23468 267430 23520
rect 59998 22244 60004 22296
rect 60056 22284 60062 22296
rect 353754 22284 353760 22296
rect 60056 22256 353760 22284
rect 60056 22244 60062 22256
rect 353754 22244 353760 22256
rect 353812 22244 353818 22296
rect 3510 22176 3516 22228
rect 3568 22216 3574 22228
rect 335814 22216 335820 22228
rect 3568 22188 335820 22216
rect 3568 22176 3574 22188
rect 335814 22176 335820 22188
rect 335872 22176 335878 22228
rect 3694 22108 3700 22160
rect 3752 22148 3758 22160
rect 346578 22148 346584 22160
rect 3752 22120 346584 22148
rect 3752 22108 3758 22120
rect 346578 22108 346584 22120
rect 346636 22108 346642 22160
rect 62298 22040 62304 22092
rect 62356 22080 62362 22092
rect 85482 22080 85488 22092
rect 62356 22052 85488 22080
rect 62356 22040 62362 22052
rect 85482 22040 85488 22052
rect 85540 22040 85546 22092
rect 200022 22040 200028 22092
rect 200080 22080 200086 22092
rect 378870 22080 378876 22092
rect 200080 22052 378876 22080
rect 200080 22040 200086 22052
rect 378870 22040 378876 22052
rect 378928 22040 378934 22092
rect 386046 22040 386052 22092
rect 386104 22080 386110 22092
rect 527818 22080 527824 22092
rect 386104 22052 527824 22080
rect 386104 22040 386110 22052
rect 527818 22040 527824 22052
rect 527876 22040 527882 22092
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 364518 22012 364524 22024
rect 20036 21984 364524 22012
rect 20036 21972 20042 21984
rect 364518 21972 364524 21984
rect 364576 21972 364582 22024
rect 3602 21904 3608 21956
rect 3660 21944 3666 21956
rect 342990 21944 342996 21956
rect 3660 21916 342996 21944
rect 3660 21904 3666 21916
rect 342990 21904 342996 21916
rect 343048 21904 343054 21956
rect 199378 21836 199384 21888
rect 199436 21876 199442 21888
rect 375282 21876 375288 21888
rect 199436 21848 375288 21876
rect 199436 21836 199442 21848
rect 375282 21836 375288 21848
rect 375340 21836 375346 21888
rect 199470 21768 199476 21820
rect 199528 21808 199534 21820
rect 350166 21808 350172 21820
rect 199528 21780 350172 21808
rect 199528 21768 199534 21780
rect 350166 21768 350172 21780
rect 350224 21768 350230 21820
rect 184842 21428 184848 21480
rect 184900 21468 184906 21480
rect 303522 21468 303528 21480
rect 184900 21440 303528 21468
rect 184900 21428 184906 21440
rect 303522 21428 303528 21440
rect 303580 21428 303586 21480
rect 151814 21360 151820 21412
rect 151872 21400 151878 21412
rect 296346 21400 296352 21412
rect 151872 21372 296352 21400
rect 151872 21360 151878 21372
rect 296346 21360 296352 21372
rect 296404 21360 296410 21412
rect 132494 20068 132500 20120
rect 132552 20108 132558 20120
rect 210234 20108 210240 20120
rect 132552 20080 210240 20108
rect 132552 20068 132558 20080
rect 210234 20068 210240 20080
rect 210292 20068 210298 20120
rect 142798 20000 142804 20052
rect 142856 20040 142862 20052
rect 281994 20040 282000 20052
rect 142856 20012 282000 20040
rect 142856 20000 142862 20012
rect 281994 20000 282000 20012
rect 282052 20000 282058 20052
rect 166994 19932 167000 19984
rect 167052 19972 167058 19984
rect 310698 19972 310704 19984
rect 167052 19944 310704 19972
rect 167052 19932 167058 19944
rect 310698 19932 310704 19944
rect 310756 19932 310762 19984
rect 175274 18708 175280 18760
rect 175332 18748 175338 18760
rect 253290 18748 253296 18760
rect 175332 18720 253296 18748
rect 175332 18708 175338 18720
rect 253290 18708 253296 18720
rect 253348 18708 253354 18760
rect 135254 18640 135260 18692
rect 135312 18680 135318 18692
rect 213822 18680 213828 18692
rect 135312 18652 213828 18680
rect 135312 18640 135318 18652
rect 213822 18640 213828 18652
rect 213880 18640 213886 18692
rect 160094 18572 160100 18624
rect 160152 18612 160158 18624
rect 184842 18612 184848 18624
rect 160152 18584 184848 18612
rect 160152 18572 160158 18584
rect 184842 18572 184848 18584
rect 184900 18572 184906 18624
rect 184934 18572 184940 18624
rect 184992 18612 184998 18624
rect 328638 18612 328644 18624
rect 184992 18584 328644 18612
rect 184992 18572 184998 18584
rect 328638 18572 328644 18584
rect 328696 18572 328702 18624
rect 171134 17348 171140 17400
rect 171192 17388 171198 17400
rect 249702 17388 249708 17400
rect 171192 17360 249708 17388
rect 171192 17348 171198 17360
rect 249702 17348 249708 17360
rect 249760 17348 249766 17400
rect 131114 17280 131120 17332
rect 131172 17320 131178 17332
rect 274818 17320 274824 17332
rect 131172 17292 274824 17320
rect 131172 17280 131178 17292
rect 274818 17280 274824 17292
rect 274876 17280 274882 17332
rect 71130 17212 71136 17264
rect 71188 17252 71194 17264
rect 242894 17252 242900 17264
rect 71188 17224 242900 17252
rect 71188 17212 71194 17224
rect 242894 17212 242900 17224
rect 242952 17212 242958 17264
rect 168374 15988 168380 16040
rect 168432 16028 168438 16040
rect 245654 16028 245660 16040
rect 168432 16000 245660 16028
rect 168432 15988 168438 16000
rect 245654 15988 245660 16000
rect 245712 15988 245718 16040
rect 135346 15920 135352 15972
rect 135404 15960 135410 15972
rect 277394 15960 277400 15972
rect 135404 15932 277400 15960
rect 135404 15920 135410 15932
rect 277394 15920 277400 15932
rect 277452 15920 277458 15972
rect 74534 15852 74540 15904
rect 74592 15892 74598 15904
rect 245930 15892 245936 15904
rect 74592 15864 245936 15892
rect 74592 15852 74598 15864
rect 245930 15852 245936 15864
rect 245988 15852 245994 15904
rect 164418 14560 164424 14612
rect 164476 14600 164482 14612
rect 241514 14600 241520 14612
rect 164476 14572 241520 14600
rect 164476 14560 164482 14572
rect 241514 14560 241520 14572
rect 241572 14560 241578 14612
rect 178586 14492 178592 14544
rect 178644 14532 178650 14544
rect 256694 14532 256700 14544
rect 178644 14504 256700 14532
rect 178644 14492 178650 14504
rect 256694 14492 256700 14504
rect 256752 14492 256758 14544
rect 173894 14424 173900 14476
rect 173952 14464 173958 14476
rect 317414 14464 317420 14476
rect 173952 14436 317420 14464
rect 173952 14424 173958 14436
rect 317414 14424 317420 14436
rect 317472 14424 317478 14476
rect 139578 13200 139584 13252
rect 139636 13240 139642 13252
rect 216674 13240 216680 13252
rect 139636 13212 216680 13240
rect 139636 13200 139642 13212
rect 216674 13200 216680 13212
rect 216732 13200 216738 13252
rect 217318 13200 217324 13252
rect 217376 13240 217382 13252
rect 284294 13240 284300 13252
rect 217376 13212 284300 13240
rect 217376 13200 217382 13212
rect 284294 13200 284300 13212
rect 284352 13200 284358 13252
rect 161290 13132 161296 13184
rect 161348 13172 161354 13184
rect 238754 13172 238760 13184
rect 161348 13144 238760 13172
rect 161348 13132 161354 13144
rect 238754 13132 238760 13144
rect 238812 13132 238818 13184
rect 176654 13064 176660 13116
rect 176712 13104 176718 13116
rect 320174 13104 320180 13116
rect 176712 13076 320180 13104
rect 176712 13064 176718 13076
rect 320174 13064 320180 13076
rect 320232 13064 320238 13116
rect 150618 11908 150624 11960
rect 150676 11948 150682 11960
rect 227714 11948 227720 11960
rect 150676 11920 227720 11948
rect 150676 11908 150682 11920
rect 227714 11908 227720 11920
rect 227772 11908 227778 11960
rect 125594 11840 125600 11892
rect 125652 11880 125658 11892
rect 202874 11880 202880 11892
rect 125652 11852 202880 11880
rect 125652 11840 125658 11852
rect 202874 11840 202880 11852
rect 202932 11840 202938 11892
rect 186130 11772 186136 11824
rect 186188 11812 186194 11824
rect 263594 11812 263600 11824
rect 186188 11784 263600 11812
rect 186188 11772 186194 11784
rect 263594 11772 263600 11784
rect 263652 11772 263658 11824
rect 145466 11704 145472 11756
rect 145524 11744 145530 11756
rect 288434 11744 288440 11756
rect 145524 11716 288440 11744
rect 145524 11704 145530 11716
rect 288434 11704 288440 11716
rect 288492 11704 288498 11756
rect 147122 10480 147128 10532
rect 147180 10520 147186 10532
rect 223574 10520 223580 10532
rect 147180 10492 223580 10520
rect 147180 10480 147186 10492
rect 223574 10480 223580 10492
rect 223632 10480 223638 10532
rect 188522 10412 188528 10464
rect 188580 10452 188586 10464
rect 331214 10452 331220 10464
rect 188580 10424 331220 10452
rect 188580 10412 188586 10424
rect 331214 10412 331220 10424
rect 331272 10412 331278 10464
rect 149514 10344 149520 10396
rect 149572 10384 149578 10396
rect 292574 10384 292580 10396
rect 149572 10356 292580 10384
rect 149572 10344 149578 10356
rect 292574 10344 292580 10356
rect 292632 10344 292638 10396
rect 3418 10276 3424 10328
rect 3476 10316 3482 10328
rect 338114 10316 338120 10328
rect 3476 10288 338120 10316
rect 3476 10276 3482 10288
rect 338114 10276 338120 10288
rect 338172 10276 338178 10328
rect 170766 9052 170772 9104
rect 170824 9092 170830 9104
rect 313274 9092 313280 9104
rect 170824 9064 313280 9092
rect 170824 9052 170830 9064
rect 313274 9052 313280 9064
rect 313332 9052 313338 9104
rect 163682 8984 163688 9036
rect 163740 9024 163746 9036
rect 306374 9024 306380 9036
rect 163740 8996 306380 9024
rect 163740 8984 163746 8996
rect 306374 8984 306380 8996
rect 306432 8984 306438 9036
rect 84194 8916 84200 8968
rect 84252 8956 84258 8968
rect 241698 8956 241704 8968
rect 84252 8928 241704 8956
rect 84252 8916 84258 8928
rect 241698 8916 241704 8928
rect 241756 8916 241762 8968
rect 157794 7692 157800 7744
rect 157852 7732 157858 7744
rect 234614 7732 234620 7744
rect 157852 7704 234620 7732
rect 157852 7692 157858 7704
rect 234614 7692 234620 7704
rect 234672 7692 234678 7744
rect 128170 7624 128176 7676
rect 128228 7664 128234 7676
rect 270494 7664 270500 7676
rect 128228 7636 270500 7664
rect 128228 7624 128234 7636
rect 270494 7624 270500 7636
rect 270552 7624 270558 7676
rect 88334 7556 88340 7608
rect 88392 7596 88398 7608
rect 245194 7596 245200 7608
rect 88392 7568 245200 7596
rect 88392 7556 88398 7568
rect 245194 7556 245200 7568
rect 245252 7556 245258 7608
rect 143534 6332 143540 6384
rect 143592 6372 143598 6384
rect 220814 6372 220820 6384
rect 143592 6344 220820 6372
rect 143592 6332 143598 6344
rect 220814 6332 220820 6344
rect 220872 6332 220878 6384
rect 181438 6264 181444 6316
rect 181496 6304 181502 6316
rect 324314 6304 324320 6316
rect 181496 6276 324320 6304
rect 181496 6264 181502 6276
rect 324314 6264 324320 6276
rect 324372 6264 324378 6316
rect 92474 6196 92480 6248
rect 92532 6236 92538 6248
rect 248782 6236 248788 6248
rect 92532 6208 248788 6236
rect 92532 6196 92538 6208
rect 248782 6196 248788 6208
rect 248840 6196 248846 6248
rect 78674 6128 78680 6180
rect 78732 6168 78738 6180
rect 249978 6168 249984 6180
rect 78732 6140 249984 6168
rect 78732 6128 78738 6140
rect 249978 6128 249984 6140
rect 250036 6128 250042 6180
rect 182542 4972 182548 5024
rect 182600 5012 182606 5024
rect 259454 5012 259460 5024
rect 182600 4984 259460 5012
rect 182600 4972 182606 4984
rect 259454 4972 259460 4984
rect 259512 4972 259518 5024
rect 154206 4904 154212 4956
rect 154264 4944 154270 4956
rect 230474 4944 230480 4956
rect 154264 4916 230480 4944
rect 154264 4904 154270 4916
rect 230474 4904 230480 4916
rect 230532 4904 230538 4956
rect 129366 4836 129372 4888
rect 129424 4876 129430 4888
rect 205634 4876 205640 4888
rect 129424 4848 205640 4876
rect 129424 4836 129430 4848
rect 205634 4836 205640 4848
rect 205692 4836 205698 4888
rect 96614 4768 96620 4820
rect 96672 4808 96678 4820
rect 252370 4808 252376 4820
rect 96672 4780 252376 4808
rect 96672 4768 96678 4780
rect 252370 4768 252376 4780
rect 252428 4768 252434 4820
rect 138842 3952 138848 4004
rect 138900 3992 138906 4004
rect 142798 3992 142804 4004
rect 138900 3964 142804 3992
rect 138900 3952 138906 3964
rect 142798 3952 142804 3964
rect 142856 3952 142862 4004
rect 135254 3544 135260 3596
rect 135312 3584 135318 3596
rect 136450 3584 136456 3596
rect 135312 3556 136456 3584
rect 135312 3544 135318 3556
rect 136450 3544 136456 3556
rect 136508 3544 136514 3596
rect 142430 3544 142436 3596
rect 142488 3584 142494 3596
rect 217318 3584 217324 3596
rect 142488 3556 217324 3584
rect 142488 3544 142494 3556
rect 217318 3544 217324 3556
rect 217376 3544 217382 3596
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153010 3516 153016 3528
rect 151872 3488 153016 3516
rect 151872 3476 151878 3488
rect 153010 3476 153016 3488
rect 153068 3476 153074 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 299474 3516 299480 3528
rect 156656 3488 299480 3516
rect 156656 3476 156662 3488
rect 299474 3476 299480 3488
rect 299532 3476 299538 3528
rect 66254 3408 66260 3460
rect 66312 3448 66318 3460
rect 239306 3448 239312 3460
rect 66312 3420 239312 3448
rect 66312 3408 66318 3420
rect 239306 3408 239312 3420
rect 239364 3408 239370 3460
rect 266354 3408 266360 3460
rect 266412 3448 266418 3460
rect 579798 3448 579804 3460
rect 266412 3420 579804 3448
rect 266412 3408 266418 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 177850 3380 177856 3392
rect 176712 3352 177856 3380
rect 176712 3340 176718 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
<< via1 >>
rect 8116 700952 8168 701004
rect 72976 700952 73028 701004
rect 397460 700952 397512 701004
rect 418160 700952 418212 701004
rect 462320 700952 462372 701004
rect 20628 700340 20680 700392
rect 89168 700340 89220 700392
rect 137836 700340 137888 700392
rect 198740 700340 198792 700392
rect 72976 700272 73028 700324
rect 199384 700272 199436 700324
rect 198740 699796 198792 699848
rect 200028 699796 200080 699848
rect 202788 699796 202840 699848
rect 20720 699660 20772 699712
rect 24308 699660 24360 699712
rect 527180 697552 527232 697604
rect 527824 697552 527876 697604
rect 580172 697552 580224 697604
rect 300860 667156 300912 667208
rect 412640 667156 412692 667208
rect 304540 586508 304592 586560
rect 477500 586508 477552 586560
rect 22008 586440 22060 586492
rect 153200 586440 153252 586492
rect 348424 586440 348476 586492
rect 350908 586440 350960 586492
rect 68652 586372 68704 586424
rect 71044 586372 71096 586424
rect 300768 586100 300820 586152
rect 309692 586100 309744 586152
rect 410156 586100 410208 586152
rect 418804 586100 418856 586152
rect 20352 586032 20404 586084
rect 29368 586032 29420 586084
rect 130476 586032 130528 586084
rect 139492 586032 139544 586084
rect 300584 586032 300636 586084
rect 312268 586032 312320 586084
rect 407580 586032 407632 586084
rect 419540 586032 419592 586084
rect 21364 585964 21416 586016
rect 31944 585964 31996 586016
rect 127900 585964 127952 586016
rect 138664 585964 138716 586016
rect 301228 585964 301280 586016
rect 314844 585964 314896 586016
rect 405004 585964 405056 586016
rect 19248 585896 19300 585948
rect 34520 585896 34572 585948
rect 125324 585896 125376 585948
rect 139400 585896 139452 585948
rect 299388 585896 299440 585948
rect 317420 585896 317472 585948
rect 402428 585896 402480 585948
rect 415124 585896 415176 585948
rect 415308 585964 415360 586016
rect 419632 585964 419684 586016
rect 418436 585896 418488 585948
rect 17868 585828 17920 585880
rect 37280 585828 37332 585880
rect 122748 585828 122800 585880
rect 138572 585828 138624 585880
rect 299112 585828 299164 585880
rect 319996 585828 320048 585880
rect 399852 585828 399904 585880
rect 418344 585828 418396 585880
rect 19156 585760 19208 585812
rect 39672 585760 39724 585812
rect 119988 585760 120040 585812
rect 139860 585760 139912 585812
rect 301412 585760 301464 585812
rect 332876 585760 332928 585812
rect 397276 585760 397328 585812
rect 419816 585760 419868 585812
rect 415124 585692 415176 585744
rect 419724 585692 419776 585744
rect 20536 585148 20588 585200
rect 26792 585148 26844 585200
rect 135628 585148 135680 585200
rect 138388 585148 138440 585200
rect 300400 585148 300452 585200
rect 307116 585148 307168 585200
rect 299296 583380 299348 583432
rect 322572 583380 322624 583432
rect 394700 583380 394752 583432
rect 420920 583380 420972 583432
rect 17776 583312 17828 583364
rect 42248 583312 42300 583364
rect 299204 583312 299256 583364
rect 325148 583312 325200 583364
rect 392124 583312 392176 583364
rect 422576 583312 422628 583364
rect 19064 583244 19116 583296
rect 44824 583244 44876 583296
rect 115020 583244 115072 583296
rect 140780 583244 140832 583296
rect 300492 583244 300544 583296
rect 330300 583244 330352 583296
rect 389548 583244 389600 583296
rect 421380 583244 421432 583296
rect 17684 583176 17736 583228
rect 49976 583176 50028 583228
rect 109868 583176 109920 583228
rect 138296 583176 138348 583228
rect 297916 583176 297968 583228
rect 340604 583176 340656 583228
rect 386972 583176 387024 583228
rect 421196 583176 421248 583228
rect 18972 583108 19024 583160
rect 57980 583108 58032 583160
rect 112444 583108 112496 583160
rect 142160 583108 142212 583160
rect 296628 583108 296680 583160
rect 343180 583108 343232 583160
rect 368940 583108 368992 583160
rect 423680 583108 423732 583160
rect 15108 583040 15160 583092
rect 73160 583040 73212 583092
rect 107292 583040 107344 583092
rect 139768 583040 139820 583092
rect 296536 583040 296588 583092
rect 353484 583040 353536 583092
rect 366364 583040 366416 583092
rect 425152 583040 425204 583092
rect 16396 582972 16448 583024
rect 75920 582972 75972 583024
rect 104716 582972 104768 583024
rect 138480 582972 138532 583024
rect 297732 582972 297784 583024
rect 356060 582972 356112 583024
rect 363788 582972 363840 583024
rect 423864 582972 423916 583024
rect 85580 544348 85632 544400
rect 142436 544348 142488 544400
rect 247040 544348 247092 544400
rect 378140 544348 378192 544400
rect 71044 542988 71096 543040
rect 262220 542988 262272 543040
rect 100760 542036 100812 542088
rect 140964 542036 141016 542088
rect 96620 541968 96672 542020
rect 142252 541968 142304 542020
rect 93860 541900 93912 541952
rect 142344 541900 142396 541952
rect 17592 541832 17644 541884
rect 59360 541832 59412 541884
rect 91100 541832 91152 541884
rect 140872 541832 140924 541884
rect 380900 541832 380952 541884
rect 421104 541832 421156 541884
rect 18880 541764 18932 541816
rect 62120 541764 62172 541816
rect 82820 541764 82872 541816
rect 142528 541764 142580 541816
rect 375380 541764 375432 541816
rect 422392 541764 422444 541816
rect 20260 541696 20312 541748
rect 64880 541696 64932 541748
rect 80060 541696 80112 541748
rect 141056 541696 141108 541748
rect 297824 541696 297876 541748
rect 345020 541696 345072 541748
rect 374000 541696 374052 541748
rect 422484 541696 422536 541748
rect 16488 541628 16540 541680
rect 77300 541628 77352 541680
rect 98000 541628 98052 541680
rect 245660 541628 245712 541680
rect 263600 541628 263652 541680
rect 348424 541628 348476 541680
rect 371240 541628 371292 541680
rect 421288 541628 421340 541680
rect 3332 514768 3384 514820
rect 7564 514768 7616 514820
rect 420828 470568 420880 470620
rect 579988 470568 580040 470620
rect 421196 465400 421248 465452
rect 421288 465196 421340 465248
rect 421104 463020 421156 463072
rect 425060 463020 425112 463072
rect 421196 462952 421248 463004
rect 20720 462612 20772 462664
rect 21640 462612 21692 462664
rect 298928 462612 298980 462664
rect 301228 462612 301280 462664
rect 314660 462612 314712 462664
rect 382096 462612 382148 462664
rect 385500 462612 385552 462664
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 419632 462408 419684 462460
rect 299112 462272 299164 462324
rect 300400 462272 300452 462324
rect 418804 462272 418856 462324
rect 419632 462272 419684 462324
rect 421196 462340 421248 462392
rect 423772 462340 423824 462392
rect 20628 462204 20680 462256
rect 24216 462204 24268 462256
rect 418160 462204 418212 462256
rect 419724 462204 419776 462256
rect 418068 462136 418120 462188
rect 421104 462272 421156 462324
rect 418436 461728 418488 461780
rect 419816 461728 419868 461780
rect 348608 461252 348660 461304
rect 350540 461252 350592 461304
rect 115020 461116 115072 461168
rect 140780 461116 140832 461168
rect 86362 461048 86414 461100
rect 142436 461048 142488 461100
rect 143540 461048 143592 461100
rect 376668 461048 376720 461100
rect 383568 461048 383620 461100
rect 83786 460980 83838 461032
rect 142528 460980 142580 461032
rect 300400 460980 300452 461032
rect 319996 460980 320048 461032
rect 371516 460980 371568 461032
rect 385500 460980 385552 461032
rect 16488 460912 16540 460964
rect 78312 460912 78364 460964
rect 81348 460912 81400 460964
rect 141056 460912 141108 460964
rect 142068 460912 142120 460964
rect 301412 460912 301464 460964
rect 332876 460912 332928 460964
rect 374092 460912 374144 460964
rect 298008 460844 298060 460896
rect 302700 460844 302752 460896
rect 358636 460844 358688 460896
rect 405004 460912 405056 460964
rect 418528 460912 418580 460964
rect 421012 460912 421064 460964
rect 422484 460844 422536 460896
rect 383568 460776 383620 460828
rect 422392 460776 422444 460828
rect 298836 460164 298888 460216
rect 345756 460164 345808 460216
rect 297824 459892 297876 459944
rect 298836 459892 298888 459944
rect 415216 459620 415268 459672
rect 419540 459620 419592 459672
rect 41420 459484 41472 459536
rect 47400 459484 47452 459536
rect 68652 459484 68704 459536
rect 71044 459484 71096 459536
rect 135628 459484 135680 459536
rect 138388 459484 138440 459536
rect 297916 459484 297968 459536
rect 340604 459484 340656 459536
rect 397276 459484 397328 459536
rect 418436 459552 418488 459604
rect 422392 459552 422444 459604
rect 423956 459552 424008 459604
rect 402428 459484 402480 459536
rect 407028 459484 407080 459536
rect 407580 459484 407632 459536
rect 415216 459484 415268 459536
rect 415308 459484 415360 459536
rect 418068 459484 418120 459536
rect 17316 459416 17368 459468
rect 60280 459416 60332 459468
rect 94412 459416 94464 459468
rect 142344 459416 142396 459468
rect 300492 459416 300544 459468
rect 330300 459416 330352 459468
rect 392124 459416 392176 459468
rect 422576 459416 422628 459468
rect 18972 459348 19024 459400
rect 57980 459348 58032 459400
rect 102048 459348 102100 459400
rect 140964 459348 141016 459400
rect 299112 459348 299164 459400
rect 325148 459348 325200 459400
rect 410156 459348 410208 459400
rect 419724 459348 419776 459400
rect 17684 459280 17736 459332
rect 49976 459280 50028 459332
rect 91836 459280 91888 459332
rect 140872 459280 140924 459332
rect 363788 459280 363840 459332
rect 423864 459280 423916 459332
rect 19064 459212 19116 459264
rect 23204 459212 23256 459264
rect 44824 459212 44876 459264
rect 417884 459212 417936 459264
rect 421472 459212 421524 459264
rect 20260 459144 20312 459196
rect 65432 459144 65484 459196
rect 300400 459144 300452 459196
rect 300676 459144 300728 459196
rect 39120 459076 39172 459128
rect 42248 459076 42300 459128
rect 112444 459008 112496 459060
rect 141148 459008 141200 459060
rect 142160 459008 142212 459060
rect 300400 459008 300452 459060
rect 327724 459008 327776 459060
rect 399852 459008 399904 459060
rect 409880 459008 409932 459060
rect 96988 458940 97040 458992
rect 140872 458940 140924 458992
rect 296628 458940 296680 458992
rect 297916 458940 297968 458992
rect 343180 458940 343232 458992
rect 394700 458940 394752 458992
rect 419816 458940 419868 458992
rect 420920 458940 420972 458992
rect 89260 458872 89312 458924
rect 135720 458872 135772 458924
rect 296536 458872 296588 458924
rect 297548 458872 297600 458924
rect 353484 458872 353536 458924
rect 366364 458872 366416 458924
rect 418160 458872 418212 458924
rect 15108 458804 15160 458856
rect 16212 458804 16264 458856
rect 73160 458804 73212 458856
rect 99288 458804 99340 458856
rect 244280 458804 244332 458856
rect 264980 458804 265032 458856
rect 348332 458804 348384 458856
rect 368940 458804 368992 458856
rect 420920 458804 420972 458856
rect 140872 458736 140924 458788
rect 141056 458736 141108 458788
rect 142252 458736 142304 458788
rect 140964 458192 141016 458244
rect 141240 458192 141292 458244
rect 297640 458192 297692 458244
rect 300492 458192 300544 458244
rect 19248 458124 19300 458176
rect 34520 458124 34572 458176
rect 107292 458124 107344 458176
rect 139768 458124 139820 458176
rect 299296 458124 299348 458176
rect 322572 458124 322624 458176
rect 384396 458124 384448 458176
rect 418068 458124 418120 458176
rect 418160 458124 418212 458176
rect 418804 458124 418856 458176
rect 425152 458124 425204 458176
rect 21272 458056 21324 458108
rect 26792 458056 26844 458108
rect 117228 458056 117280 458108
rect 139676 458056 139728 458108
rect 299388 458056 299440 458108
rect 317420 458056 317472 458108
rect 409880 458056 409932 458108
rect 418344 458056 418396 458108
rect 420920 458056 420972 458108
rect 421564 458056 421616 458108
rect 423680 458056 423732 458108
rect 125324 457988 125376 458040
rect 139400 457988 139452 458040
rect 130476 457920 130528 457972
rect 139584 457920 139636 457972
rect 21364 457648 21416 457700
rect 31944 457648 31996 457700
rect 300584 457648 300636 457700
rect 301228 457648 301280 457700
rect 17868 457580 17920 457632
rect 19064 457512 19116 457564
rect 21364 457512 21416 457564
rect 37188 457512 37240 457564
rect 20536 457444 20588 457496
rect 21272 457444 21324 457496
rect 17776 457376 17828 457428
rect 20444 457376 20496 457428
rect 39120 457444 39172 457496
rect 301228 457444 301280 457496
rect 312268 457444 312320 457496
rect 139676 457104 139728 457156
rect 139952 457104 140004 457156
rect 419540 457036 419592 457088
rect 419816 457036 419868 457088
rect 139400 456832 139452 456884
rect 140044 456832 140096 456884
rect 17868 456764 17920 456816
rect 18880 456764 18932 456816
rect 18972 456764 19024 456816
rect 19248 456764 19300 456816
rect 139584 456764 139636 456816
rect 139768 456764 139820 456816
rect 299020 456764 299072 456816
rect 299296 456764 299348 456816
rect 418252 456764 418304 456816
rect 418528 456764 418580 456816
rect 300860 456696 300912 456748
rect 301504 456696 301556 456748
rect 361212 456696 361264 456748
rect 297732 456628 297784 456680
rect 356060 456628 356112 456680
rect 16396 455336 16448 455388
rect 17868 455336 17920 455388
rect 17592 454656 17644 454708
rect 17868 454656 17920 454708
rect 75920 454656 75972 454708
rect 248420 416032 248472 416084
rect 378140 416032 378192 416084
rect 71044 413244 71096 413296
rect 260840 413244 260892 413296
rect 2780 410048 2832 410100
rect 4988 410048 5040 410100
rect 3700 398828 3752 398880
rect 19984 398828 20036 398880
rect 3332 345040 3384 345092
rect 20076 345040 20128 345092
rect 16304 333208 16356 333260
rect 18788 333208 18840 333260
rect 57704 333208 57756 333260
rect 96988 333004 97040 333056
rect 141056 333004 141108 333056
rect 115020 332936 115072 332988
rect 140780 332936 140832 332988
rect 142160 332936 142212 332988
rect 15016 332868 15068 332920
rect 17776 332868 17828 332920
rect 47400 332868 47452 332920
rect 91836 332868 91888 332920
rect 140872 332868 140924 332920
rect 300676 332868 300728 332920
rect 318800 332868 318852 332920
rect 319996 332868 320048 332920
rect 17684 332800 17736 332852
rect 49976 332800 50028 332852
rect 112444 332800 112496 332852
rect 141148 332800 141200 332852
rect 299020 332800 299072 332852
rect 321560 332800 321612 332852
rect 322572 332800 322624 332852
rect 16396 332732 16448 332784
rect 73160 332732 73212 332784
rect 107292 332732 107344 332784
rect 139308 332732 139360 332784
rect 299112 332732 299164 332784
rect 324320 332732 324372 332784
rect 325148 332732 325200 332784
rect 17408 332664 17460 332716
rect 17592 332664 17644 332716
rect 75920 332664 75972 332716
rect 109868 332664 109920 332716
rect 142252 332664 142304 332716
rect 300400 332664 300452 332716
rect 327264 332800 327316 332852
rect 416688 332800 416740 332852
rect 418804 332800 418856 332852
rect 16488 332596 16540 332648
rect 78312 332596 78364 332648
rect 104716 332596 104768 332648
rect 138296 332596 138348 332648
rect 138572 332596 138624 332648
rect 297640 332596 297692 332648
rect 329840 332596 329892 332648
rect 3608 332528 3660 332580
rect 21640 332528 21692 332580
rect 68652 332528 68704 332580
rect 71044 332528 71096 332580
rect 94412 332528 94464 332580
rect 96528 332528 96580 332580
rect 135628 332528 135680 332580
rect 138388 332528 138440 332580
rect 300308 332528 300360 332580
rect 307116 332528 307168 332580
rect 19156 332460 19208 332512
rect 39672 332460 39724 332512
rect 119988 332460 120040 332512
rect 139768 332460 139820 332512
rect 303528 332460 303580 332512
rect 310980 332460 311032 332512
rect 18880 332392 18932 332444
rect 37280 332392 37332 332444
rect 122656 332392 122708 332444
rect 138756 332392 138808 332444
rect 301320 332392 301372 332444
rect 335452 332528 335504 332580
rect 348332 332528 348384 332580
rect 350908 332528 350960 332580
rect 366364 332528 366416 332580
rect 386512 332732 386564 332784
rect 421196 332732 421248 332784
rect 371516 332664 371568 332716
rect 383660 332664 383712 332716
rect 384396 332664 384448 332716
rect 418528 332664 418580 332716
rect 423772 332596 423824 332648
rect 424048 332596 424100 332648
rect 415308 332528 415360 332580
rect 421104 332528 421156 332580
rect 311164 332392 311216 332444
rect 338028 332460 338080 332512
rect 399852 332460 399904 332512
rect 418436 332460 418488 332512
rect 21272 332324 21324 332376
rect 26792 332324 26844 332376
rect 27528 332324 27580 332376
rect 44824 332324 44876 332376
rect 125324 332324 125376 332376
rect 140044 332324 140096 332376
rect 301044 332324 301096 332376
rect 312268 332324 312320 332376
rect 18972 332256 19024 332308
rect 34520 332256 34572 332308
rect 127900 332256 127952 332308
rect 138848 332256 138900 332308
rect 301412 332256 301464 332308
rect 332876 332392 332928 332444
rect 402428 332392 402480 332444
rect 418712 332392 418764 332444
rect 407580 332324 407632 332376
rect 419632 332324 419684 332376
rect 410156 332256 410208 332308
rect 419908 332256 419960 332308
rect 19064 332188 19116 332240
rect 31944 332188 31996 332240
rect 130476 332188 130528 332240
rect 139676 332188 139728 332240
rect 397276 332188 397328 332240
rect 418620 332188 418672 332240
rect 20352 332120 20404 332172
rect 29368 332120 29420 332172
rect 117228 332120 117280 332172
rect 139952 332120 140004 332172
rect 300584 332120 300636 332172
rect 309692 332120 309744 332172
rect 20536 332052 20588 332104
rect 42248 332052 42300 332104
rect 306748 331916 306800 331968
rect 314844 331916 314896 331968
rect 266360 331848 266412 331900
rect 348332 331848 348384 331900
rect 350540 331848 350592 331900
rect 358636 331848 358688 331900
rect 405004 331848 405056 331900
rect 419448 331848 419500 331900
rect 139492 331576 139544 331628
rect 139952 331576 140004 331628
rect 376668 331372 376720 331424
rect 382464 331372 382516 331424
rect 418620 331304 418672 331356
rect 420092 331304 420144 331356
rect 19248 331236 19300 331288
rect 20352 331236 20404 331288
rect 89260 331236 89312 331288
rect 91008 331236 91060 331288
rect 138756 331236 138808 331288
rect 139584 331236 139636 331288
rect 300216 331236 300268 331288
rect 301412 331236 301464 331288
rect 311900 331236 311952 331288
rect 317420 331236 317472 331288
rect 368940 331236 368992 331288
rect 373264 331236 373316 331288
rect 374092 331236 374144 331288
rect 379428 331236 379480 331288
rect 381820 331236 381872 331288
rect 386328 331236 386380 331288
rect 418436 331236 418488 331288
rect 420000 331236 420052 331288
rect 303528 331168 303580 331220
rect 350540 331168 350592 331220
rect 363788 331168 363840 331220
rect 299296 331100 299348 331152
rect 311900 331100 311952 331152
rect 418804 331100 418856 331152
rect 419632 331100 419684 331152
rect 423772 331032 423824 331084
rect 139492 330964 139544 331016
rect 140044 330964 140096 331016
rect 419448 330964 419500 331016
rect 421012 330964 421064 331016
rect 298836 330488 298888 330540
rect 301228 330488 301280 330540
rect 345756 330488 345808 330540
rect 17592 329740 17644 329792
rect 20260 329740 20312 329792
rect 20996 329740 21048 329792
rect 62856 329740 62908 329792
rect 84016 329740 84068 329792
rect 142436 329740 142488 329792
rect 382464 329740 382516 329792
rect 417424 329740 417476 329792
rect 419816 329740 419868 329792
rect 421564 329740 421616 329792
rect 65432 329672 65484 329724
rect 102140 329672 102192 329724
rect 140964 329672 141016 329724
rect 142528 329672 142580 329724
rect 386328 329672 386380 329724
rect 425060 329672 425112 329724
rect 16212 329604 16264 329656
rect 17316 329604 17368 329656
rect 60280 329604 60332 329656
rect 392124 329604 392176 329656
rect 393228 329604 393280 329656
rect 393320 329604 393372 329656
rect 389548 329536 389600 329588
rect 390468 329536 390520 329588
rect 422668 329604 422720 329656
rect 393504 329536 393556 329588
rect 422576 329536 422628 329588
rect 394700 329400 394752 329452
rect 395988 329400 396040 329452
rect 417424 329468 417476 329520
rect 423680 329468 423732 329520
rect 423956 329468 424008 329520
rect 419540 329400 419592 329452
rect 91008 329196 91060 329248
rect 138664 329196 138716 329248
rect 86684 329128 86736 329180
rect 140780 329128 140832 329180
rect 412732 329128 412784 329180
rect 422484 329128 422536 329180
rect 81348 329060 81400 329112
rect 141516 329060 141568 329112
rect 373264 329060 373316 329112
rect 419816 329060 419868 329112
rect 140780 327700 140832 327752
rect 142068 327700 142120 327752
rect 143540 327700 143592 327752
rect 140780 327564 140832 327616
rect 141148 327564 141200 327616
rect 3608 318792 3660 318844
rect 17224 318792 17276 318844
rect 2780 292816 2832 292868
rect 4896 292816 4948 292868
rect 300768 288328 300820 288380
rect 360200 288328 360252 288380
rect 297732 288260 297784 288312
rect 356060 288260 356112 288312
rect 249800 287648 249852 287700
rect 378140 287648 378192 287700
rect 296628 287036 296680 287088
rect 297732 287036 297784 287088
rect 297824 285608 297876 285660
rect 342260 285608 342312 285660
rect 298008 285540 298060 285592
rect 339500 285540 339552 285592
rect 395988 285268 396040 285320
rect 423956 285268 424008 285320
rect 300400 285200 300452 285252
rect 318800 285200 318852 285252
rect 393228 285200 393280 285252
rect 422576 285200 422628 285252
rect 299204 285132 299256 285184
rect 321560 285132 321612 285184
rect 390468 285132 390520 285184
rect 421012 285132 421064 285184
rect 297916 285064 297968 285116
rect 324320 285064 324372 285116
rect 383660 285064 383712 285116
rect 418252 285064 418304 285116
rect 136640 284996 136692 285048
rect 296076 284996 296128 285048
rect 299020 284996 299072 285048
rect 327080 284996 327132 285048
rect 386420 284996 386472 285048
rect 421196 284996 421248 285048
rect 71044 284928 71096 284980
rect 258080 284928 258132 284980
rect 299112 284928 299164 284980
rect 329840 284928 329892 284980
rect 379428 284928 379480 284980
rect 425152 284928 425204 284980
rect 297732 284316 297784 284368
rect 298008 284316 298060 284368
rect 416688 284316 416740 284368
rect 418528 284316 418580 284368
rect 2780 266364 2832 266416
rect 6184 266364 6236 266416
rect 2780 240184 2832 240236
rect 5080 240184 5132 240236
rect 2780 213936 2832 213988
rect 6276 213936 6328 213988
rect 300952 206592 301004 206644
rect 301136 206592 301188 206644
rect 301044 206456 301096 206508
rect 301412 206456 301464 206508
rect 140780 206320 140832 206372
rect 142068 206320 142120 206372
rect 143540 206320 143592 206372
rect 371608 206252 371660 206304
rect 424048 206252 424100 206304
rect 141240 205572 141292 205624
rect 142528 205572 142580 205624
rect 420920 205368 420972 205420
rect 422668 205368 422720 205420
rect 298928 204892 298980 204944
rect 300400 204892 300452 204944
rect 309048 204892 309100 204944
rect 297548 204824 297600 204876
rect 299020 204824 299072 204876
rect 297916 204756 297968 204808
rect 300308 204756 300360 204808
rect 298008 204688 298060 204740
rect 299112 204688 299164 204740
rect 372620 204688 372672 204740
rect 419540 205028 419592 205080
rect 86684 204620 86736 204672
rect 140780 204620 140832 204672
rect 394700 204620 394752 204672
rect 423956 204960 424008 205012
rect 425244 204960 425296 205012
rect 421564 204892 421616 204944
rect 425152 204892 425204 204944
rect 418252 204688 418304 204740
rect 418436 204688 418488 204740
rect 115020 204552 115072 204604
rect 142160 204552 142212 204604
rect 301412 204552 301464 204604
rect 365628 204552 365680 204604
rect 392124 204552 392176 204604
rect 422576 204552 422628 204604
rect 424048 204552 424100 204604
rect 102048 204484 102100 204536
rect 141240 204484 141292 204536
rect 300308 204484 300360 204536
rect 325148 204484 325200 204536
rect 389548 204484 389600 204536
rect 420920 204484 420972 204536
rect 96988 204416 97040 204468
rect 141148 204416 141200 204468
rect 299020 204416 299072 204468
rect 327724 204416 327776 204468
rect 386972 204416 387024 204468
rect 421196 204416 421248 204468
rect 19064 204348 19116 204400
rect 31944 204348 31996 204400
rect 94412 204348 94464 204400
rect 142344 204348 142396 204400
rect 299112 204348 299164 204400
rect 330300 204348 330352 204400
rect 384396 204348 384448 204400
rect 418436 204348 418488 204400
rect 19156 204280 19208 204332
rect 39672 204280 39724 204332
rect 138020 204280 138072 204332
rect 138664 204280 138716 204332
rect 143632 204280 143684 204332
rect 295248 204280 295300 204332
rect 297640 204280 297692 204332
rect 353484 204280 353536 204332
rect 374092 204280 374144 204332
rect 421380 204280 421432 204332
rect 421564 204280 421616 204332
rect 7564 204212 7616 204264
rect 21640 204212 21692 204264
rect 22008 204212 22060 204264
rect 16212 204144 16264 204196
rect 30932 204144 30984 204196
rect 21456 204076 21508 204128
rect 26792 204076 26844 204128
rect 68652 204212 68704 204264
rect 70584 204212 70636 204264
rect 71044 204212 71096 204264
rect 127900 204212 127952 204264
rect 130016 204212 130068 204264
rect 130476 204212 130528 204264
rect 133788 204212 133840 204264
rect 31116 204144 31168 204196
rect 60280 204144 60332 204196
rect 84016 204144 84068 204196
rect 142436 204144 142488 204196
rect 299112 204144 299164 204196
rect 299388 204144 299440 204196
rect 300584 204144 300636 204196
rect 307116 204212 307168 204264
rect 309048 204212 309100 204264
rect 319996 204212 320048 204264
rect 348332 204212 348384 204264
rect 350908 204212 350960 204264
rect 368940 204212 368992 204264
rect 372620 204212 372672 204264
rect 397276 204212 397328 204264
rect 411260 204212 411312 204264
rect 415308 204212 415360 204264
rect 416780 204212 416832 204264
rect 65432 204076 65484 204128
rect 89260 204076 89312 204128
rect 138020 204076 138072 204128
rect 300492 204076 300544 204128
rect 332876 204144 332928 204196
rect 365628 204144 365680 204196
rect 371516 204144 371568 204196
rect 402428 204144 402480 204196
rect 418344 204144 418396 204196
rect 16304 204008 16356 204060
rect 57980 204008 58032 204060
rect 91836 204008 91888 204060
rect 141056 204008 141108 204060
rect 299296 204008 299348 204060
rect 317420 204076 317472 204128
rect 410156 204076 410208 204128
rect 419632 204212 419684 204264
rect 419448 204144 419500 204196
rect 419908 204144 419960 204196
rect 302792 204008 302844 204060
rect 314844 204008 314896 204060
rect 405004 204008 405056 204060
rect 17684 203940 17736 203992
rect 49976 203940 50028 203992
rect 112444 203940 112496 203992
rect 140872 203940 140924 203992
rect 301320 203940 301372 203992
rect 312268 203940 312320 203992
rect 319352 203940 319404 203992
rect 322572 203940 322624 203992
rect 407580 203940 407632 203992
rect 418804 203940 418856 203992
rect 17776 203872 17828 203924
rect 47400 203872 47452 203924
rect 81348 203872 81400 203924
rect 141516 203872 141568 203924
rect 300676 203872 300728 203924
rect 309692 203872 309744 203924
rect 399852 203872 399904 203924
rect 419724 203872 419776 203924
rect 16120 203804 16172 203856
rect 16396 203804 16448 203856
rect 73160 203804 73212 203856
rect 299112 203804 299164 203856
rect 302792 203804 302844 203856
rect 303528 203804 303580 203856
rect 338028 203804 338080 203856
rect 99196 203600 99248 203652
rect 240140 203600 240192 203652
rect 133052 203532 133104 203584
rect 282184 203532 282236 203584
rect 352564 203532 352616 203584
rect 358636 203532 358688 203584
rect 125324 203464 125376 203516
rect 128268 203464 128320 203516
rect 117228 203396 117280 203448
rect 119988 203396 120040 203448
rect 122564 203328 122616 203380
rect 125508 203328 125560 203380
rect 141240 203260 141292 203312
rect 141516 203260 141568 203312
rect 376668 203124 376720 203176
rect 382648 203124 382700 203176
rect 366364 203056 366416 203108
rect 370136 203056 370188 203108
rect 381820 202920 381872 202972
rect 385408 202920 385460 202972
rect 412732 202852 412784 202904
rect 421288 202852 421340 202904
rect 20536 202784 20588 202836
rect 23296 202784 23348 202836
rect 42248 202784 42300 202836
rect 107292 202784 107344 202836
rect 138020 202784 138072 202836
rect 138480 202784 138532 202836
rect 139492 202784 139544 202836
rect 125508 202716 125560 202768
rect 139584 202716 139636 202768
rect 138020 202648 138072 202700
rect 139308 202648 139360 202700
rect 139676 202648 139728 202700
rect 128268 202104 128320 202156
rect 138480 202104 138532 202156
rect 300768 201424 300820 201476
rect 361212 201424 361264 201476
rect 363788 201424 363840 201476
rect 423864 201424 423916 201476
rect 296628 201356 296680 201408
rect 356060 201356 356112 201408
rect 370136 201356 370188 201408
rect 418528 201356 418580 201408
rect 300952 201288 301004 201340
rect 345756 201288 345808 201340
rect 382648 201288 382700 201340
rect 423680 201288 423732 201340
rect 385408 201220 385460 201272
rect 425060 201220 425112 201272
rect 299020 200608 299072 200660
rect 300952 200608 301004 200660
rect 17592 200064 17644 200116
rect 75920 200064 75972 200116
rect 16488 199384 16540 199436
rect 20536 199384 20588 199436
rect 77300 199384 77352 199436
rect 252560 164840 252612 164892
rect 378140 164840 378192 164892
rect 303528 158652 303580 158704
rect 352564 158652 352616 158704
rect 297824 158584 297876 158636
rect 342260 158584 342312 158636
rect 297732 158516 297784 158568
rect 339500 158516 339552 158568
rect 136640 158040 136692 158092
rect 297364 158040 297416 158092
rect 71044 157972 71096 158024
rect 256700 157972 256752 158024
rect 269120 157972 269172 158024
rect 348424 157972 348476 158024
rect 2780 149472 2832 149524
rect 5172 149472 5224 149524
rect 3332 136620 3384 136672
rect 13084 136620 13136 136672
rect 135628 78616 135680 78668
rect 138572 78616 138624 78668
rect 300584 78616 300636 78668
rect 306656 78616 306708 78668
rect 410432 78276 410484 78328
rect 419632 78276 419684 78328
rect 407856 78208 407908 78260
rect 418620 78208 418672 78260
rect 405280 78140 405332 78192
rect 419908 78140 419960 78192
rect 297548 78072 297600 78124
rect 327172 78072 327224 78124
rect 327356 78072 327408 78124
rect 398840 78072 398892 78124
rect 400128 78072 400180 78124
rect 419724 78072 419776 78124
rect 300400 78004 300452 78056
rect 330484 78004 330536 78056
rect 332600 78004 332652 78056
rect 396172 78004 396224 78056
rect 397368 78004 397420 78056
rect 419816 78004 419868 78056
rect 130476 77936 130528 77988
rect 139768 77936 139820 77988
rect 269764 77936 269816 77988
rect 369860 77936 369912 77988
rect 393320 77936 393372 77988
rect 422392 77936 422444 77988
rect 68652 77324 68704 77376
rect 70584 77324 70636 77376
rect 348608 77324 348660 77376
rect 350540 77324 350592 77376
rect 77300 77052 77352 77104
rect 78634 77052 78686 77104
rect 390560 76644 390612 76696
rect 421472 76644 421524 76696
rect 301136 76576 301188 76628
rect 329932 76576 329984 76628
rect 378232 76576 378284 76628
rect 421288 76576 421340 76628
rect 299020 76508 299072 76560
rect 336740 76508 336792 76560
rect 376760 76508 376812 76560
rect 422484 76508 422536 76560
rect 20536 75964 20588 76016
rect 77300 75964 77352 76016
rect 17592 75896 17644 75948
rect 75920 75896 75972 75948
rect 304540 75896 304592 75948
rect 580540 75896 580592 75948
rect 18972 75828 19024 75880
rect 34520 75828 34572 75880
rect 91836 75828 91888 75880
rect 140780 75828 140832 75880
rect 141056 75828 141108 75880
rect 333980 75828 334032 75880
rect 334624 75828 334676 75880
rect 338028 75828 338080 75880
rect 17868 75760 17920 75812
rect 63224 75760 63276 75812
rect 107292 75760 107344 75812
rect 139492 75760 139544 75812
rect 139676 75760 139728 75812
rect 322940 75760 322992 75812
rect 325148 75760 325200 75812
rect 327080 75760 327132 75812
rect 330300 75760 330352 75812
rect 336740 75760 336792 75812
rect 345756 75828 345808 75880
rect 363788 75828 363840 75880
rect 423864 75828 423916 75880
rect 386972 75760 387024 75812
rect 421196 75760 421248 75812
rect 16212 75692 16264 75744
rect 60648 75692 60700 75744
rect 112444 75692 112496 75744
rect 140872 75692 140924 75744
rect 329932 75692 329984 75744
rect 335452 75692 335504 75744
rect 384948 75692 385000 75744
rect 418436 75692 418488 75744
rect 16304 75624 16356 75676
rect 57980 75624 58032 75676
rect 122564 75624 122616 75676
rect 139584 75624 139636 75676
rect 389548 75624 389600 75676
rect 422668 75624 422720 75676
rect 17684 75556 17736 75608
rect 50344 75556 50396 75608
rect 125324 75556 125376 75608
rect 138480 75556 138532 75608
rect 300308 75556 300360 75608
rect 322940 75556 322992 75608
rect 17776 75488 17828 75540
rect 47584 75488 47636 75540
rect 119988 75488 120040 75540
rect 131120 75488 131172 75540
rect 298008 75488 298060 75540
rect 327080 75488 327132 75540
rect 16120 75420 16172 75472
rect 73528 75420 73580 75472
rect 127900 75420 127952 75472
rect 138388 75420 138440 75472
rect 297732 75420 297784 75472
rect 332600 75420 332652 75472
rect 340604 75420 340656 75472
rect 57980 75352 58032 75404
rect 59268 75352 59320 75404
rect 140780 75352 140832 75404
rect 210424 75352 210476 75404
rect 280804 75352 280856 75404
rect 379244 75352 379296 75404
rect 379520 75352 379572 75404
rect 412732 75352 412784 75404
rect 133052 75284 133104 75336
rect 231124 75284 231176 75336
rect 273260 75284 273312 75336
rect 384396 75284 384448 75336
rect 384948 75284 385000 75336
rect 71228 75216 71280 75268
rect 77944 75216 77996 75268
rect 140872 75216 140924 75268
rect 254584 75216 254636 75268
rect 277400 75216 277452 75268
rect 389548 75216 389600 75268
rect 34520 75148 34572 75200
rect 100024 75148 100076 75200
rect 139492 75148 139544 75200
rect 285680 75148 285732 75200
rect 297824 75148 297876 75200
rect 335360 75148 335412 75200
rect 343180 75148 343232 75200
rect 351184 75148 351236 75200
rect 386972 75148 387024 75200
rect 396080 75148 396132 75200
rect 417884 75148 417936 75200
rect 21456 74468 21508 74520
rect 27160 74468 27212 74520
rect 300676 74468 300728 74520
rect 309692 74468 309744 74520
rect 368940 74468 368992 74520
rect 419540 74468 419592 74520
rect 16396 74400 16448 74452
rect 44824 74400 44876 74452
rect 298928 74400 298980 74452
rect 319444 74400 319496 74452
rect 376668 74400 376720 74452
rect 423772 74400 423824 74452
rect 18788 74332 18840 74384
rect 37464 74332 37516 74384
rect 299296 74332 299348 74384
rect 318064 74332 318116 74384
rect 381452 74332 381504 74384
rect 425152 74332 425204 74384
rect 19064 74264 19116 74316
rect 32404 74264 32456 74316
rect 299112 74264 299164 74316
rect 315304 74264 315356 74316
rect 392584 74264 392636 74316
rect 424048 74264 424100 74316
rect 18880 74196 18932 74248
rect 29644 74196 29696 74248
rect 301320 74196 301372 74248
rect 312544 74196 312596 74248
rect 394700 74196 394752 74248
rect 425244 74196 425296 74248
rect 21272 74128 21324 74180
rect 55864 74128 55916 74180
rect 56508 74128 56560 74180
rect 299204 74128 299256 74180
rect 322572 74128 322624 74180
rect 402244 74128 402296 74180
rect 418344 74128 418396 74180
rect 415308 74060 415360 74112
rect 421104 74060 421156 74112
rect 138388 73788 138440 73840
rect 308680 73788 308732 73840
rect 394700 73516 394752 73568
rect 395344 73516 395396 73568
rect 309692 73176 309744 73228
rect 311164 73176 311216 73228
rect 321928 73176 321980 73228
rect 322572 73176 322624 73228
rect 376024 73176 376076 73228
rect 376668 73176 376720 73228
rect 414664 73176 414716 73228
rect 415308 73176 415360 73228
rect 104624 73108 104676 73160
rect 138296 73108 138348 73160
rect 138296 72700 138348 72752
rect 283840 72700 283892 72752
rect 75920 72632 75972 72684
rect 224224 72632 224276 72684
rect 300400 72632 300452 72684
rect 409880 72632 409932 72684
rect 212632 72564 212684 72616
rect 363788 72564 363840 72616
rect 139584 72496 139636 72548
rect 305368 72496 305420 72548
rect 59268 72428 59320 72480
rect 357440 72428 357492 72480
rect 270592 71204 270644 71256
rect 348332 71204 348384 71256
rect 137928 71136 137980 71188
rect 381544 71136 381596 71188
rect 37464 71068 37516 71120
rect 345112 71068 345164 71120
rect 27160 71000 27212 71052
rect 338488 71000 338540 71052
rect 3056 70388 3108 70440
rect 199476 70388 199528 70440
rect 81348 70320 81400 70372
rect 141148 70320 141200 70372
rect 141148 69912 141200 69964
rect 227720 69912 227772 69964
rect 73528 69844 73580 69896
rect 222568 69844 222620 69896
rect 298744 69844 298796 69896
rect 407120 69844 407172 69896
rect 215944 69776 215996 69828
rect 368940 69776 368992 69828
rect 139860 69708 139912 69760
rect 303712 69708 303764 69760
rect 60648 69640 60700 69692
rect 360200 69640 360252 69692
rect 84016 68960 84068 69012
rect 142436 68960 142488 69012
rect 143448 68960 143500 69012
rect 117228 68892 117280 68944
rect 139400 68892 139452 68944
rect 143448 68484 143500 68536
rect 229192 68484 229244 68536
rect 229744 68484 229796 68536
rect 368480 68484 368532 68536
rect 138480 68416 138532 68468
rect 290464 68416 290516 68468
rect 297088 68416 297140 68468
rect 404360 68416 404412 68468
rect 139400 68348 139452 68400
rect 302240 68348 302292 68400
rect 63224 68280 63276 68332
rect 361672 68280 361724 68332
rect 77944 66988 77996 67040
rect 255688 66988 255740 67040
rect 292120 66988 292172 67040
rect 396172 66988 396224 67040
rect 56508 66920 56560 66972
rect 356704 66920 356756 66972
rect 42064 66852 42116 66904
rect 348424 66852 348476 66904
rect 88340 66172 88392 66224
rect 143632 66172 143684 66224
rect 144828 66172 144880 66224
rect 295340 66172 295392 66224
rect 296628 66172 296680 66224
rect 356060 66172 356112 66224
rect 93860 66104 93912 66156
rect 142344 66104 142396 66156
rect 143448 66104 143500 66156
rect 96620 66036 96672 66088
rect 140780 66036 140832 66088
rect 141056 66036 141108 66088
rect 144828 65696 144880 65748
rect 232504 65696 232556 65748
rect 207664 65628 207716 65680
rect 295340 65628 295392 65680
rect 143448 65560 143500 65612
rect 236000 65560 236052 65612
rect 254032 65560 254084 65612
rect 280804 65560 280856 65612
rect 293960 65560 294012 65612
rect 398840 65560 398892 65612
rect 140780 65492 140832 65544
rect 237472 65492 237524 65544
rect 272248 65492 272300 65544
rect 381452 65492 381504 65544
rect 214288 64336 214340 64388
rect 366364 64336 366416 64388
rect 50344 64268 50396 64320
rect 353392 64268 353444 64320
rect 47584 64200 47636 64252
rect 351920 64200 351972 64252
rect 44824 64132 44876 64184
rect 350080 64132 350132 64184
rect 300768 63452 300820 63504
rect 360292 63452 360344 63504
rect 211160 62976 211212 63028
rect 300768 62976 300820 63028
rect 65524 62908 65576 62960
rect 322940 62908 322992 62960
rect 32404 62840 32456 62892
rect 341800 62840 341852 62892
rect 29644 62772 29696 62824
rect 340144 62772 340196 62824
rect 340236 62772 340288 62824
rect 392584 62772 392636 62824
rect 13084 62024 13136 62076
rect 57060 62024 57112 62076
rect 100760 62024 100812 62076
rect 140780 62024 140832 62076
rect 301412 62024 301464 62076
rect 371332 62024 371384 62076
rect 98368 61684 98420 61736
rect 239128 61684 239180 61736
rect 217600 61548 217652 61600
rect 301412 61548 301464 61600
rect 280528 61480 280580 61532
rect 395344 61480 395396 61532
rect 140780 61412 140832 61464
rect 141424 61412 141476 61464
rect 282092 61412 282144 61464
rect 282184 61412 282236 61464
rect 366640 61412 366692 61464
rect 220912 61344 220964 61396
rect 376024 61344 376076 61396
rect 294052 60664 294104 60716
rect 295248 60664 295300 60716
rect 353300 60664 353352 60716
rect 302332 60596 302384 60648
rect 357532 60596 357584 60648
rect 206008 60120 206060 60172
rect 294052 60120 294104 60172
rect 231124 60052 231176 60104
rect 364984 60052 365036 60104
rect 219440 59984 219492 60036
rect 374644 59984 374696 60036
rect 209320 59372 209372 59424
rect 302332 59372 302384 59424
rect 135260 58828 135312 58880
rect 204352 58828 204404 58880
rect 210424 58828 210476 58880
rect 234160 58828 234212 58880
rect 254584 58828 254636 58880
rect 288808 58828 288860 58880
rect 295432 58828 295484 58880
rect 402244 58828 402296 58880
rect 129740 58760 129792 58812
rect 307116 58760 307168 58812
rect 202880 58692 202932 58744
rect 414664 58692 414716 58744
rect 100024 58624 100076 58676
rect 343640 58624 343692 58676
rect 109040 57876 109092 57928
rect 142252 57876 142304 57928
rect 143448 57876 143500 57928
rect 311164 57876 311216 57928
rect 314016 57876 314068 57928
rect 318064 57876 318116 57928
rect 318984 57876 319036 57928
rect 319444 57876 319496 57928
rect 320640 57876 320692 57928
rect 328920 57876 328972 57928
rect 330484 57876 330536 57928
rect 114560 57808 114612 57860
rect 142160 57808 142212 57860
rect 143356 57808 143408 57860
rect 306380 57808 306432 57860
rect 312360 57808 312412 57860
rect 312544 57808 312596 57860
rect 315672 57808 315724 57860
rect 332232 57740 332284 57792
rect 334624 57740 334676 57792
rect 290464 57536 290516 57588
rect 307392 57604 307444 57656
rect 322940 57536 322992 57588
rect 363696 57536 363748 57588
rect 279240 57468 279292 57520
rect 340236 57468 340288 57520
rect 275928 57400 275980 57452
rect 351184 57400 351236 57452
rect 297364 57332 297416 57384
rect 383568 57332 383620 57384
rect 143448 57264 143500 57316
rect 287520 57264 287572 57316
rect 296076 57264 296128 57316
rect 385224 57264 385276 57316
rect 395160 57264 395212 57316
rect 418252 57264 418304 57316
rect 143356 57196 143408 57248
rect 290832 57196 290884 57248
rect 295984 57196 296036 57248
rect 388536 57196 388588 57248
rect 390192 57196 390244 57248
rect 422300 57196 422352 57248
rect 307116 56924 307168 56976
rect 310704 56924 310756 56976
rect 315304 56584 315356 56636
rect 317328 56584 317380 56636
rect 325608 56584 325660 56636
rect 327172 56584 327224 56636
rect 5172 56516 5224 56568
rect 57520 56516 57572 56568
rect 102140 55224 102192 55276
rect 196624 55224 196676 55276
rect 102140 53864 102192 53916
rect 103888 53864 103940 53916
rect 399484 53048 399536 53100
rect 580264 53048 580316 53100
rect 102140 52504 102192 52556
rect 196164 52504 196216 52556
rect 102232 52436 102284 52488
rect 103980 52436 104032 52488
rect 5080 52368 5132 52420
rect 57060 52368 57112 52420
rect 102876 52368 102928 52420
rect 195980 52368 196032 52420
rect 103152 52300 103204 52352
rect 196072 52300 196124 52352
rect 103060 51008 103112 51060
rect 195980 51008 196032 51060
rect 102140 49784 102192 49836
rect 104348 49784 104400 49836
rect 102784 49648 102836 49700
rect 195980 49648 196032 49700
rect 102600 49580 102652 49632
rect 196072 49580 196124 49632
rect 103888 48220 103940 48272
rect 195980 48220 196032 48272
rect 6184 46860 6236 46912
rect 57520 46860 57572 46912
rect 103980 46860 104032 46912
rect 195980 46860 196032 46912
rect 103244 45500 103296 45552
rect 195980 45500 196032 45552
rect 3332 44140 3384 44192
rect 60004 44140 60056 44192
rect 102876 44072 102928 44124
rect 196072 44072 196124 44124
rect 104348 44004 104400 44056
rect 195980 44004 196032 44056
rect 3516 42712 3568 42764
rect 57152 42712 57204 42764
rect 102600 42712 102652 42764
rect 196072 42712 196124 42764
rect 102968 42644 103020 42696
rect 195980 42644 196032 42696
rect 103520 41352 103572 41404
rect 195980 41352 196032 41404
rect 102140 40672 102192 40724
rect 196164 40672 196216 40724
rect 102324 39992 102376 40044
rect 196072 39992 196124 40044
rect 103612 39924 103664 39976
rect 195980 39924 196032 39976
rect 102232 38564 102284 38616
rect 195980 38564 196032 38616
rect 6276 37204 6328 37256
rect 57060 37204 57112 37256
rect 102140 37204 102192 37256
rect 195980 37204 196032 37256
rect 102784 35844 102836 35896
rect 195980 35844 196032 35896
rect 102600 35776 102652 35828
rect 196072 35776 196124 35828
rect 102692 34416 102744 34468
rect 196072 34416 196124 34468
rect 102876 34348 102928 34400
rect 195980 34348 196032 34400
rect 102140 33056 102192 33108
rect 195980 33056 196032 33108
rect 4896 31696 4948 31748
rect 57612 31696 57664 31748
rect 102140 31696 102192 31748
rect 196072 31696 196124 31748
rect 102324 31628 102376 31680
rect 195980 31628 196032 31680
rect 102140 30268 102192 30320
rect 196072 30268 196124 30320
rect 102232 30200 102284 30252
rect 195980 30200 196032 30252
rect 102140 28908 102192 28960
rect 195980 28908 196032 28960
rect 102140 28228 102192 28280
rect 195980 28228 196032 28280
rect 17224 27548 17276 27600
rect 57244 27548 57296 27600
rect 102140 27548 102192 27600
rect 195980 27548 196032 27600
rect 102784 26188 102836 26240
rect 195980 26188 196032 26240
rect 397184 24624 397236 24676
rect 399484 24624 399536 24676
rect 20628 24216 20680 24268
rect 356980 24216 357032 24268
rect 20076 24148 20128 24200
rect 360660 24148 360712 24200
rect 3424 24080 3476 24132
rect 371332 24080 371384 24132
rect 85488 23468 85540 23520
rect 266360 23468 266412 23520
rect 267372 23468 267424 23520
rect 60004 22244 60056 22296
rect 353760 22244 353812 22296
rect 3516 22176 3568 22228
rect 335820 22176 335872 22228
rect 3700 22108 3752 22160
rect 346584 22108 346636 22160
rect 62304 22040 62356 22092
rect 85488 22040 85540 22092
rect 200028 22040 200080 22092
rect 378876 22040 378928 22092
rect 386052 22040 386104 22092
rect 527824 22040 527876 22092
rect 19984 21972 20036 22024
rect 364524 21972 364576 22024
rect 3608 21904 3660 21956
rect 342996 21904 343048 21956
rect 199384 21836 199436 21888
rect 375288 21836 375340 21888
rect 199476 21768 199528 21820
rect 350172 21768 350224 21820
rect 184848 21428 184900 21480
rect 303528 21428 303580 21480
rect 151820 21360 151872 21412
rect 296352 21360 296404 21412
rect 132500 20068 132552 20120
rect 210240 20068 210292 20120
rect 142804 20000 142856 20052
rect 282000 20000 282052 20052
rect 167000 19932 167052 19984
rect 310704 19932 310756 19984
rect 175280 18708 175332 18760
rect 253296 18708 253348 18760
rect 135260 18640 135312 18692
rect 213828 18640 213880 18692
rect 160100 18572 160152 18624
rect 184848 18572 184900 18624
rect 184940 18572 184992 18624
rect 328644 18572 328696 18624
rect 171140 17348 171192 17400
rect 249708 17348 249760 17400
rect 131120 17280 131172 17332
rect 274824 17280 274876 17332
rect 71136 17212 71188 17264
rect 242900 17212 242952 17264
rect 168380 15988 168432 16040
rect 245660 15988 245712 16040
rect 135352 15920 135404 15972
rect 277400 15920 277452 15972
rect 74540 15852 74592 15904
rect 245936 15852 245988 15904
rect 164424 14560 164476 14612
rect 241520 14560 241572 14612
rect 178592 14492 178644 14544
rect 256700 14492 256752 14544
rect 173900 14424 173952 14476
rect 317420 14424 317472 14476
rect 139584 13200 139636 13252
rect 216680 13200 216732 13252
rect 217324 13200 217376 13252
rect 284300 13200 284352 13252
rect 161296 13132 161348 13184
rect 238760 13132 238812 13184
rect 176660 13064 176712 13116
rect 320180 13064 320232 13116
rect 150624 11908 150676 11960
rect 227720 11908 227772 11960
rect 125600 11840 125652 11892
rect 202880 11840 202932 11892
rect 186136 11772 186188 11824
rect 263600 11772 263652 11824
rect 145472 11704 145524 11756
rect 288440 11704 288492 11756
rect 147128 10480 147180 10532
rect 223580 10480 223632 10532
rect 188528 10412 188580 10464
rect 331220 10412 331272 10464
rect 149520 10344 149572 10396
rect 292580 10344 292632 10396
rect 3424 10276 3476 10328
rect 338120 10276 338172 10328
rect 170772 9052 170824 9104
rect 313280 9052 313332 9104
rect 163688 8984 163740 9036
rect 306380 8984 306432 9036
rect 84200 8916 84252 8968
rect 241704 8916 241756 8968
rect 157800 7692 157852 7744
rect 234620 7692 234672 7744
rect 128176 7624 128228 7676
rect 270500 7624 270552 7676
rect 88340 7556 88392 7608
rect 245200 7556 245252 7608
rect 143540 6332 143592 6384
rect 220820 6332 220872 6384
rect 181444 6264 181496 6316
rect 324320 6264 324372 6316
rect 92480 6196 92532 6248
rect 248788 6196 248840 6248
rect 78680 6128 78732 6180
rect 249984 6128 250036 6180
rect 182548 4972 182600 5024
rect 259460 4972 259512 5024
rect 154212 4904 154264 4956
rect 230480 4904 230532 4956
rect 129372 4836 129424 4888
rect 205640 4836 205692 4888
rect 96620 4768 96672 4820
rect 252376 4768 252428 4820
rect 138848 3952 138900 4004
rect 142804 3952 142856 4004
rect 135260 3544 135312 3596
rect 136456 3544 136508 3596
rect 142436 3544 142488 3596
rect 217324 3544 217376 3596
rect 151820 3476 151872 3528
rect 153016 3476 153068 3528
rect 156604 3476 156656 3528
rect 299480 3476 299532 3528
rect 66260 3408 66312 3460
rect 239312 3408 239364 3460
rect 266360 3408 266412 3460
rect 579804 3408 579856 3460
rect 176660 3340 176712 3392
rect 177856 3340 177908 3392
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 701010 8156 703520
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 20628 700392 20680 700398
rect 20628 700334 20680 700340
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 607209 2820 658135
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 2778 607200 2834 607209
rect 2778 607135 2834 607144
rect 3422 607200 3478 607209
rect 3422 607135 3478 607144
rect 3436 606121 3464 607135
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 2778 410544 2834 410553
rect 2778 410479 2834 410488
rect 2792 410106 2820 410479
rect 2780 410100 2832 410106
rect 2780 410042 2832 410048
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 2778 267200 2834 267209
rect 2778 267135 2834 267144
rect 2792 266422 2820 267135
rect 2780 266416 2832 266422
rect 2780 266358 2832 266364
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 2792 213994 2820 214911
rect 2780 213988 2832 213994
rect 2780 213930 2832 213936
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 2792 149530 2820 149767
rect 2780 149524 2832 149530
rect 2780 149466 2832 149472
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3054 71632 3110 71641
rect 3054 71567 3110 71576
rect 3068 70446 3096 71567
rect 3056 70440 3108 70446
rect 3056 70382 3108 70388
rect 3330 45520 3386 45529
rect 3330 45455 3386 45464
rect 3344 44198 3372 45455
rect 3332 44192 3384 44198
rect 3332 44134 3384 44140
rect 3436 24138 3464 606047
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 204105 3556 566879
rect 3620 332586 3648 619103
rect 20352 586084 20404 586090
rect 20352 586026 20404 586032
rect 19248 585948 19300 585954
rect 19248 585890 19300 585896
rect 17868 585880 17920 585886
rect 17868 585822 17920 585828
rect 17776 583364 17828 583370
rect 17776 583306 17828 583312
rect 17684 583228 17736 583234
rect 17684 583170 17736 583176
rect 15108 583092 15160 583098
rect 15108 583034 15160 583040
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3712 502489 3740 553823
rect 7564 514820 7616 514826
rect 7564 514762 7616 514768
rect 3698 502480 3754 502489
rect 3698 502415 3754 502424
rect 3712 501809 3740 502415
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3712 398886 3740 449511
rect 3700 398880 3752 398886
rect 3700 398822 3752 398828
rect 3712 397497 3740 398822
rect 3698 397488 3754 397497
rect 3698 397423 3754 397432
rect 3608 332580 3660 332586
rect 3608 332522 3660 332528
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3620 318850 3648 319223
rect 3608 318844 3660 318850
rect 3608 318786 3660 318792
rect 3514 204096 3570 204105
rect 3514 204031 3570 204040
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3528 42770 3556 188799
rect 3606 110664 3662 110673
rect 3606 110599 3662 110608
rect 3516 42764 3568 42770
rect 3516 42706 3568 42712
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3528 22234 3556 32399
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3620 21962 3648 110599
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 3712 22166 3740 84623
rect 4816 75857 4844 462538
rect 4988 410100 5040 410106
rect 4988 410042 5040 410048
rect 4896 292868 4948 292874
rect 4896 292810 4948 292816
rect 4802 75848 4858 75857
rect 4802 75783 4858 75792
rect 4908 31754 4936 292810
rect 5000 75721 5028 410042
rect 6184 266416 6236 266422
rect 6184 266358 6236 266364
rect 5080 240236 5132 240242
rect 5080 240178 5132 240184
rect 4986 75712 5042 75721
rect 4986 75647 5042 75656
rect 5092 52426 5120 240178
rect 5172 149524 5224 149530
rect 5172 149466 5224 149472
rect 5184 56574 5212 149466
rect 5172 56568 5224 56574
rect 5172 56510 5224 56516
rect 5080 52420 5132 52426
rect 5080 52362 5132 52368
rect 6196 46918 6224 266358
rect 6276 213988 6328 213994
rect 6276 213930 6328 213936
rect 6184 46912 6236 46918
rect 6184 46854 6236 46860
rect 6288 37262 6316 213930
rect 7576 204270 7604 514762
rect 15014 460184 15070 460193
rect 15014 460119 15070 460128
rect 15028 332926 15056 460119
rect 15120 458862 15148 583034
rect 16396 583024 16448 583030
rect 16396 582966 16448 582972
rect 15108 458856 15160 458862
rect 15108 458798 15160 458804
rect 16212 458856 16264 458862
rect 16212 458798 16264 458804
rect 16224 345014 16252 458798
rect 16408 455394 16436 582966
rect 17592 541884 17644 541890
rect 17592 541826 17644 541832
rect 16488 541680 16540 541686
rect 16488 541622 16540 541628
rect 16500 460970 16528 541622
rect 16488 460964 16540 460970
rect 17604 460934 17632 541826
rect 16488 460906 16540 460912
rect 17328 460906 17632 460934
rect 16396 455388 16448 455394
rect 16396 455330 16448 455336
rect 16224 344986 16436 345014
rect 16304 333260 16356 333266
rect 16304 333202 16356 333208
rect 15016 332920 15068 332926
rect 15016 332862 15068 332868
rect 16212 329656 16264 329662
rect 16212 329598 16264 329604
rect 7564 204264 7616 204270
rect 7564 204206 7616 204212
rect 16224 204202 16252 329598
rect 16212 204196 16264 204202
rect 16212 204138 16264 204144
rect 16120 203856 16172 203862
rect 16120 203798 16172 203804
rect 13084 136672 13136 136678
rect 13084 136614 13136 136620
rect 13096 62082 13124 136614
rect 16132 75478 16160 203798
rect 16224 75750 16252 204138
rect 16316 204066 16344 333202
rect 16408 332790 16436 344986
rect 16396 332784 16448 332790
rect 16396 332726 16448 332732
rect 16304 204060 16356 204066
rect 16304 204002 16356 204008
rect 16212 75744 16264 75750
rect 16212 75686 16264 75692
rect 16316 75682 16344 204002
rect 16408 203862 16436 332726
rect 16500 332654 16528 460906
rect 17328 459474 17356 460906
rect 17316 459468 17368 459474
rect 17316 459410 17368 459416
rect 16488 332648 16540 332654
rect 16488 332590 16540 332596
rect 16396 203856 16448 203862
rect 16396 203798 16448 203804
rect 16394 203552 16450 203561
rect 16394 203487 16450 203496
rect 16304 75676 16356 75682
rect 16304 75618 16356 75624
rect 16120 75472 16172 75478
rect 16120 75414 16172 75420
rect 16408 74458 16436 203487
rect 16500 199442 16528 332590
rect 17328 329662 17356 459410
rect 17696 459338 17724 583170
rect 17684 459332 17736 459338
rect 17684 459274 17736 459280
rect 17406 458280 17462 458289
rect 17406 458215 17462 458224
rect 17420 345014 17448 458215
rect 17592 454708 17644 454714
rect 17592 454650 17644 454656
rect 17420 344986 17540 345014
rect 17408 332716 17460 332722
rect 17408 332658 17460 332664
rect 17316 329656 17368 329662
rect 17316 329598 17368 329604
rect 17420 325694 17448 332658
rect 17512 330290 17540 344986
rect 17604 332722 17632 454650
rect 17696 332858 17724 459274
rect 17788 457434 17816 583306
rect 17880 457638 17908 585822
rect 19156 585812 19208 585818
rect 19156 585754 19208 585760
rect 19064 583296 19116 583302
rect 19064 583238 19116 583244
rect 18972 583160 19024 583166
rect 18972 583102 19024 583108
rect 18880 541816 18932 541822
rect 18880 541758 18932 541764
rect 18892 459513 18920 541758
rect 18878 459504 18934 459513
rect 18878 459439 18934 459448
rect 18892 458289 18920 459439
rect 18984 459406 19012 583102
rect 18972 459400 19024 459406
rect 18972 459342 19024 459348
rect 18878 458280 18934 458289
rect 18878 458215 18934 458224
rect 17868 457632 17920 457638
rect 17868 457574 17920 457580
rect 17776 457428 17828 457434
rect 17776 457370 17828 457376
rect 17880 456822 17908 457574
rect 18984 457178 19012 459342
rect 19076 459270 19104 583238
rect 19064 459264 19116 459270
rect 19064 459206 19116 459212
rect 19168 458017 19196 585754
rect 19260 458182 19288 585890
rect 20166 585848 20222 585857
rect 20166 585783 20222 585792
rect 19248 458176 19300 458182
rect 19248 458118 19300 458124
rect 19154 458008 19210 458017
rect 19154 457943 19210 457952
rect 19064 457564 19116 457570
rect 19064 457506 19116 457512
rect 18800 457150 19012 457178
rect 17868 456816 17920 456822
rect 17868 456758 17920 456764
rect 17868 455388 17920 455394
rect 17868 455330 17920 455336
rect 17880 454714 17908 455330
rect 17868 454708 17920 454714
rect 17868 454650 17920 454656
rect 18800 333266 18828 457150
rect 18880 456816 18932 456822
rect 18880 456758 18932 456764
rect 18972 456816 19024 456822
rect 18972 456758 19024 456764
rect 18788 333260 18840 333266
rect 18788 333202 18840 333208
rect 17776 332920 17828 332926
rect 17776 332862 17828 332868
rect 17684 332852 17736 332858
rect 17684 332794 17736 332800
rect 17592 332716 17644 332722
rect 17592 332658 17644 332664
rect 17512 330262 17632 330290
rect 17604 329798 17632 330262
rect 17592 329792 17644 329798
rect 17592 329734 17644 329740
rect 17420 325666 17540 325694
rect 17224 318844 17276 318850
rect 17224 318786 17276 318792
rect 16488 199436 16540 199442
rect 16488 199378 16540 199384
rect 16396 74452 16448 74458
rect 16396 74394 16448 74400
rect 13084 62076 13136 62082
rect 13084 62018 13136 62024
rect 6276 37256 6328 37262
rect 6276 37198 6328 37204
rect 4896 31748 4948 31754
rect 4896 31690 4948 31696
rect 17236 27606 17264 318786
rect 17512 200114 17540 325666
rect 17604 204241 17632 329734
rect 17590 204232 17646 204241
rect 17590 204167 17646 204176
rect 17696 203998 17724 332794
rect 17684 203992 17736 203998
rect 17684 203934 17736 203940
rect 17592 200116 17644 200122
rect 17512 200086 17592 200114
rect 17592 200058 17644 200064
rect 17604 75954 17632 200058
rect 17592 75948 17644 75954
rect 17592 75890 17644 75896
rect 17696 75614 17724 203934
rect 17788 203930 17816 332862
rect 18892 332450 18920 456758
rect 18880 332444 18932 332450
rect 18880 332386 18932 332392
rect 18892 209774 18920 332386
rect 18984 332314 19012 456758
rect 18972 332308 19024 332314
rect 18972 332250 19024 332256
rect 18800 209746 18920 209774
rect 18800 204377 18828 209746
rect 18984 204513 19012 332250
rect 19076 332246 19104 457506
rect 19168 332518 19196 457943
rect 19260 456822 19288 458118
rect 20180 457473 20208 585783
rect 20260 541748 20312 541754
rect 20260 541690 20312 541696
rect 20272 459202 20300 541690
rect 20364 459377 20392 586026
rect 20536 585200 20588 585206
rect 20536 585142 20588 585148
rect 20350 459368 20406 459377
rect 20350 459303 20406 459312
rect 20260 459196 20312 459202
rect 20260 459138 20312 459144
rect 20166 457464 20222 457473
rect 20166 457399 20222 457408
rect 19248 456816 19300 456822
rect 19248 456758 19300 456764
rect 19984 398880 20036 398886
rect 19984 398822 20036 398828
rect 19156 332512 19208 332518
rect 19156 332454 19208 332460
rect 19064 332240 19116 332246
rect 19064 332182 19116 332188
rect 18970 204504 19026 204513
rect 18970 204439 19026 204448
rect 18786 204368 18842 204377
rect 18786 204303 18842 204312
rect 17866 204232 17922 204241
rect 17866 204167 17922 204176
rect 17880 203969 17908 204167
rect 17866 203960 17922 203969
rect 17776 203924 17828 203930
rect 17866 203895 17922 203904
rect 17776 203866 17828 203872
rect 17684 75608 17736 75614
rect 17684 75550 17736 75556
rect 17788 75546 17816 203866
rect 17880 75818 17908 203895
rect 17868 75812 17920 75818
rect 17868 75754 17920 75760
rect 17776 75540 17828 75546
rect 17776 75482 17828 75488
rect 18800 74390 18828 204303
rect 18878 202872 18934 202881
rect 18878 202807 18934 202816
rect 18788 74384 18840 74390
rect 18788 74326 18840 74332
rect 18892 74254 18920 202807
rect 18984 75886 19012 204439
rect 19076 204406 19104 332182
rect 19064 204400 19116 204406
rect 19064 204342 19116 204348
rect 18972 75880 19024 75886
rect 18972 75822 19024 75828
rect 19076 74322 19104 204342
rect 19168 204338 19196 332454
rect 19248 331288 19300 331294
rect 19248 331230 19300 331236
rect 19156 204332 19208 204338
rect 19156 204274 19208 204280
rect 19168 74361 19196 204274
rect 19260 202881 19288 331230
rect 19246 202872 19302 202881
rect 19246 202807 19302 202816
rect 19154 74352 19210 74361
rect 19064 74316 19116 74322
rect 19154 74287 19210 74296
rect 19064 74258 19116 74264
rect 18880 74248 18932 74254
rect 18880 74190 18932 74196
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 19996 22030 20024 398822
rect 20076 345092 20128 345098
rect 20076 345034 20128 345040
rect 20088 24206 20116 345034
rect 20272 329798 20300 459138
rect 20364 332178 20392 459303
rect 20548 457502 20576 585142
rect 20640 462262 20668 700334
rect 24320 699718 24348 703520
rect 72988 701010 73016 703520
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 72988 700330 73016 700946
rect 89180 700398 89208 703520
rect 137848 700398 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 20720 699712 20772 699718
rect 20720 699654 20772 699660
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 20732 462670 20760 699654
rect 21974 587058 22002 587316
rect 24564 587302 24808 587330
rect 21974 587030 22048 587058
rect 22020 586498 22048 587030
rect 22008 586492 22060 586498
rect 22008 586434 22060 586440
rect 24780 586401 24808 587302
rect 26804 587302 27140 587330
rect 29380 587302 29716 587330
rect 31956 587302 32292 587330
rect 34532 587302 34868 587330
rect 37292 587302 37444 587330
rect 39684 587302 40020 587330
rect 42260 587302 42596 587330
rect 44836 587302 45172 587330
rect 47412 587302 47748 587330
rect 49988 587302 50324 587330
rect 52564 587302 52900 587330
rect 55232 587302 55476 587330
rect 57992 587302 58052 587330
rect 59372 587302 60628 587330
rect 62132 587302 63204 587330
rect 64892 587302 65780 587330
rect 68356 587302 68692 587330
rect 70932 587302 71084 587330
rect 24766 586392 24822 586401
rect 24766 586327 24822 586336
rect 21364 586016 21416 586022
rect 21364 585958 21416 585964
rect 20720 462664 20772 462670
rect 20720 462606 20772 462612
rect 20628 462256 20680 462262
rect 20628 462198 20680 462204
rect 21272 458108 21324 458114
rect 21272 458050 21324 458056
rect 21284 457502 21312 458050
rect 21376 457706 21404 585958
rect 21454 585712 21510 585721
rect 21454 585647 21510 585656
rect 21468 458153 21496 585647
rect 26804 585206 26832 587302
rect 29380 586090 29408 587302
rect 29368 586084 29420 586090
rect 29368 586026 29420 586032
rect 31956 586022 31984 587302
rect 31944 586016 31996 586022
rect 31944 585958 31996 585964
rect 34532 585954 34560 587302
rect 34520 585948 34572 585954
rect 34520 585890 34572 585896
rect 37292 585886 37320 587302
rect 37280 585880 37332 585886
rect 37280 585822 37332 585828
rect 39684 585818 39712 587302
rect 39672 585812 39724 585818
rect 39672 585754 39724 585760
rect 26792 585200 26844 585206
rect 26792 585142 26844 585148
rect 42260 583370 42288 587302
rect 42248 583364 42300 583370
rect 42248 583306 42300 583312
rect 44836 583302 44864 587302
rect 44824 583296 44876 583302
rect 44824 583238 44876 583244
rect 47412 583001 47440 587302
rect 49988 583234 50016 587302
rect 52564 585857 52592 587302
rect 52550 585848 52606 585857
rect 52550 585783 52606 585792
rect 55232 585721 55260 587302
rect 55218 585712 55274 585721
rect 55218 585647 55274 585656
rect 49976 583228 50028 583234
rect 49976 583170 50028 583176
rect 57992 583166 58020 587302
rect 57980 583160 58032 583166
rect 57980 583102 58032 583108
rect 47398 582992 47454 583001
rect 47398 582927 47454 582936
rect 59372 541890 59400 587302
rect 59360 541884 59412 541890
rect 59360 541826 59412 541832
rect 62132 541822 62160 587302
rect 62120 541816 62172 541822
rect 62120 541758 62172 541764
rect 64892 541754 64920 587302
rect 68664 586430 68692 587302
rect 71056 586430 71084 587302
rect 73172 587302 73508 587330
rect 75932 587302 76084 587330
rect 77312 587302 78660 587330
rect 80072 587302 81236 587330
rect 82832 587302 83812 587330
rect 85592 587302 86388 587330
rect 88352 587302 88964 587330
rect 91112 587302 91540 587330
rect 93872 587302 94116 587330
rect 96632 587302 96692 587330
rect 98012 587302 99268 587330
rect 100772 587302 101844 587330
rect 104420 587302 104756 587330
rect 106996 587302 107332 587330
rect 109572 587302 109908 587330
rect 112148 587302 112484 587330
rect 114724 587302 115060 587330
rect 68652 586424 68704 586430
rect 68652 586366 68704 586372
rect 71044 586424 71096 586430
rect 71044 586366 71096 586372
rect 71056 543046 71084 586366
rect 73172 583098 73200 587302
rect 73160 583092 73212 583098
rect 73160 583034 73212 583040
rect 75932 583030 75960 587302
rect 75920 583024 75972 583030
rect 75920 582966 75972 582972
rect 71044 543040 71096 543046
rect 71044 542982 71096 542988
rect 64880 541748 64932 541754
rect 64880 541690 64932 541696
rect 77312 541686 77340 587302
rect 80072 541754 80100 587302
rect 82832 541822 82860 587302
rect 85592 544406 85620 587302
rect 85580 544400 85632 544406
rect 85580 544342 85632 544348
rect 82820 541816 82872 541822
rect 88352 541793 88380 587302
rect 91112 541890 91140 587302
rect 93872 541958 93900 587302
rect 96632 542026 96660 587302
rect 96620 542020 96672 542026
rect 96620 541962 96672 541968
rect 93860 541952 93912 541958
rect 93860 541894 93912 541900
rect 91100 541884 91152 541890
rect 91100 541826 91152 541832
rect 82820 541758 82872 541764
rect 88338 541784 88394 541793
rect 80060 541748 80112 541754
rect 88338 541719 88394 541728
rect 80060 541690 80112 541696
rect 98012 541686 98040 587302
rect 100772 542094 100800 587302
rect 104728 583030 104756 587302
rect 107304 583098 107332 587302
rect 109880 583234 109908 587302
rect 109868 583228 109920 583234
rect 109868 583170 109920 583176
rect 112456 583166 112484 587302
rect 115032 583302 115060 587302
rect 117240 587302 117300 587330
rect 119876 587302 120028 587330
rect 122452 587302 122788 587330
rect 125028 587302 125364 587330
rect 127604 587302 127940 587330
rect 130180 587302 130516 587330
rect 132756 587302 133092 587330
rect 135332 587302 135668 587330
rect 117240 585857 117268 587302
rect 117226 585848 117282 585857
rect 120000 585818 120028 587302
rect 122760 585886 122788 587302
rect 125336 585954 125364 587302
rect 127912 586022 127940 587302
rect 130488 586090 130516 587302
rect 130476 586084 130528 586090
rect 130476 586026 130528 586032
rect 127900 586016 127952 586022
rect 127900 585958 127952 585964
rect 125324 585948 125376 585954
rect 125324 585890 125376 585896
rect 122748 585880 122800 585886
rect 122748 585822 122800 585828
rect 117226 585783 117282 585792
rect 119988 585812 120040 585818
rect 119988 585754 120040 585760
rect 133064 585721 133092 587302
rect 133050 585712 133106 585721
rect 133050 585647 133106 585656
rect 135640 585206 135668 587302
rect 136652 587302 137908 587330
rect 135628 585200 135680 585206
rect 135628 585142 135680 585148
rect 115020 583296 115072 583302
rect 115020 583238 115072 583244
rect 112444 583160 112496 583166
rect 112444 583102 112496 583108
rect 107292 583092 107344 583098
rect 107292 583034 107344 583040
rect 104716 583024 104768 583030
rect 104716 582966 104768 582972
rect 100760 542088 100812 542094
rect 100760 542030 100812 542036
rect 77300 541680 77352 541686
rect 77300 541622 77352 541628
rect 98000 541680 98052 541686
rect 136652 541657 136680 587302
rect 153212 586498 153240 702406
rect 198740 700392 198792 700398
rect 198740 700334 198792 700340
rect 198752 699854 198780 700334
rect 199384 700324 199436 700330
rect 199384 700266 199436 700272
rect 198740 699848 198792 699854
rect 198740 699790 198792 699796
rect 153200 586492 153252 586498
rect 153200 586434 153252 586440
rect 139492 586084 139544 586090
rect 139492 586026 139544 586032
rect 138664 586016 138716 586022
rect 138664 585958 138716 585964
rect 138572 585880 138624 585886
rect 138572 585822 138624 585828
rect 138388 585200 138440 585206
rect 138388 585142 138440 585148
rect 138296 583228 138348 583234
rect 138296 583170 138348 583176
rect 98000 541622 98052 541628
rect 136638 541648 136694 541657
rect 136638 541583 136694 541592
rect 21640 462664 21692 462670
rect 21692 462612 21988 462618
rect 21640 462606 21988 462612
rect 21652 462590 21988 462606
rect 24216 462256 24268 462262
rect 24268 462204 24564 462210
rect 24216 462198 24564 462204
rect 24228 462182 24564 462198
rect 26804 461230 27140 461258
rect 29380 461230 29716 461258
rect 31956 461230 32292 461258
rect 34532 461230 34868 461258
rect 37292 461230 37444 461258
rect 39684 461230 40020 461258
rect 42260 461230 42596 461258
rect 44836 461230 45172 461258
rect 47412 461230 47748 461258
rect 49988 461230 50324 461258
rect 52564 461230 52900 461258
rect 55232 461230 55476 461258
rect 57992 461230 58052 461258
rect 60292 461230 60628 461258
rect 62868 461230 63204 461258
rect 65444 461230 65780 461258
rect 68356 461230 68692 461258
rect 70932 461230 71084 461258
rect 23204 459264 23256 459270
rect 23204 459206 23256 459212
rect 23216 458289 23244 459206
rect 23202 458280 23258 458289
rect 23202 458215 23258 458224
rect 21454 458144 21510 458153
rect 26804 458114 26832 461230
rect 29380 459377 29408 461230
rect 29366 459368 29422 459377
rect 29366 459303 29422 459312
rect 21454 458079 21510 458088
rect 26792 458108 26844 458114
rect 21364 457700 21416 457706
rect 21364 457642 21416 457648
rect 21376 457570 21404 457642
rect 21364 457564 21416 457570
rect 21364 457506 21416 457512
rect 20536 457496 20588 457502
rect 20536 457438 20588 457444
rect 21272 457496 21324 457502
rect 21272 457438 21324 457444
rect 21362 457464 21418 457473
rect 20444 457428 20496 457434
rect 20444 457370 20496 457376
rect 20456 345014 20484 457370
rect 20456 344986 20576 345014
rect 20352 332172 20404 332178
rect 20352 332114 20404 332120
rect 20364 331294 20392 332114
rect 20548 332110 20576 344986
rect 21284 332382 21312 457438
rect 21362 457399 21418 457408
rect 21376 332489 21404 457399
rect 21362 332480 21418 332489
rect 21362 332415 21418 332424
rect 21272 332376 21324 332382
rect 21272 332318 21324 332324
rect 20536 332104 20588 332110
rect 20536 332046 20588 332052
rect 20352 331288 20404 331294
rect 20352 331230 20404 331236
rect 20260 329792 20312 329798
rect 20260 329734 20312 329740
rect 20548 202842 20576 332046
rect 21086 331392 21142 331401
rect 21086 331327 21142 331336
rect 20626 331256 20682 331265
rect 20626 331191 20682 331200
rect 20536 202836 20588 202842
rect 20536 202778 20588 202784
rect 20536 199436 20588 199442
rect 20536 199378 20588 199384
rect 20548 76022 20576 199378
rect 20536 76016 20588 76022
rect 20536 75958 20588 75964
rect 20640 24274 20668 331191
rect 20996 329792 21048 329798
rect 20994 329760 20996 329769
rect 21048 329760 21050 329769
rect 20994 329695 21050 329704
rect 21100 202881 21128 331327
rect 21178 331256 21234 331265
rect 21178 331191 21234 331200
rect 21192 209774 21220 331191
rect 21284 229094 21312 332318
rect 21376 331265 21404 332415
rect 21468 332217 21496 458079
rect 26792 458050 26844 458056
rect 31956 457706 31984 461230
rect 34532 458182 34560 461230
rect 37292 458266 37320 461230
rect 39120 459128 39172 459134
rect 39120 459070 39172 459076
rect 37200 458238 37320 458266
rect 34520 458176 34572 458182
rect 34520 458118 34572 458124
rect 31944 457700 31996 457706
rect 31944 457642 31996 457648
rect 37200 457570 37228 458238
rect 37188 457564 37240 457570
rect 37188 457506 37240 457512
rect 39132 457502 39160 459070
rect 39684 458017 39712 461230
rect 41418 460184 41474 460193
rect 41418 460119 41474 460128
rect 41432 459542 41460 460119
rect 41420 459536 41472 459542
rect 41420 459478 41472 459484
rect 42260 459134 42288 461230
rect 44836 459270 44864 461230
rect 47412 459542 47440 461230
rect 47400 459536 47452 459542
rect 47400 459478 47452 459484
rect 49988 459338 50016 461230
rect 49976 459332 50028 459338
rect 49976 459274 50028 459280
rect 44824 459264 44876 459270
rect 44824 459206 44876 459212
rect 42248 459128 42300 459134
rect 42248 459070 42300 459076
rect 39670 458008 39726 458017
rect 39670 457943 39726 457952
rect 39120 457496 39172 457502
rect 52564 457473 52592 461230
rect 55232 458153 55260 461230
rect 57992 459406 58020 461230
rect 60292 459474 60320 461230
rect 62868 459513 62896 461230
rect 62854 459504 62910 459513
rect 60280 459468 60332 459474
rect 62854 459439 62910 459448
rect 60280 459410 60332 459416
rect 57980 459400 58032 459406
rect 57980 459342 58032 459348
rect 65444 459202 65472 461230
rect 68664 459542 68692 461230
rect 71056 459542 71084 461230
rect 73172 461230 73508 461258
rect 75932 461230 76084 461258
rect 78324 461230 78660 461258
rect 81236 461230 81388 461258
rect 68652 459536 68704 459542
rect 68652 459478 68704 459484
rect 71044 459536 71096 459542
rect 71044 459478 71096 459484
rect 65432 459196 65484 459202
rect 65432 459138 65484 459144
rect 55218 458144 55274 458153
rect 55218 458079 55274 458088
rect 39120 457438 39172 457444
rect 52550 457464 52606 457473
rect 52550 457399 52606 457408
rect 71056 413302 71084 459478
rect 73172 458862 73200 461230
rect 73160 458856 73212 458862
rect 73160 458798 73212 458804
rect 75932 454714 75960 461230
rect 78324 460970 78352 461230
rect 81360 460970 81388 461230
rect 83798 461038 83826 461244
rect 86374 461106 86402 461244
rect 88964 461230 89300 461258
rect 91540 461230 91876 461258
rect 94116 461230 94452 461258
rect 96692 461230 97028 461258
rect 86362 461100 86414 461106
rect 86362 461042 86414 461048
rect 83786 461032 83838 461038
rect 83786 460974 83838 460980
rect 78312 460964 78364 460970
rect 78312 460906 78364 460912
rect 81348 460964 81400 460970
rect 81348 460906 81400 460912
rect 89272 458930 89300 461230
rect 91848 459338 91876 461230
rect 94424 459474 94452 461230
rect 94412 459468 94464 459474
rect 94412 459410 94464 459416
rect 91836 459332 91888 459338
rect 91836 459274 91888 459280
rect 97000 458998 97028 461230
rect 99254 461122 99282 461244
rect 101844 461230 102088 461258
rect 104420 461230 104756 461258
rect 106996 461230 107332 461258
rect 109572 461230 109908 461258
rect 112148 461230 112484 461258
rect 114724 461230 115060 461258
rect 99254 461094 99328 461122
rect 96988 458992 97040 458998
rect 96988 458934 97040 458940
rect 89260 458924 89312 458930
rect 89260 458866 89312 458872
rect 99300 458862 99328 461094
rect 102060 459406 102088 461230
rect 102048 459400 102100 459406
rect 102048 459342 102100 459348
rect 99288 458856 99340 458862
rect 99288 458798 99340 458804
rect 104728 458153 104756 461230
rect 107304 458182 107332 461230
rect 107292 458176 107344 458182
rect 104714 458144 104770 458153
rect 107292 458118 107344 458124
rect 104714 458079 104770 458088
rect 109880 458017 109908 461230
rect 112456 459066 112484 461230
rect 115032 461174 115060 461230
rect 117240 461230 117300 461258
rect 119876 461230 120028 461258
rect 122452 461230 122788 461258
rect 125028 461230 125364 461258
rect 127604 461230 127940 461258
rect 130180 461230 130516 461258
rect 132756 461230 133092 461258
rect 135332 461230 135668 461258
rect 115020 461168 115072 461174
rect 115020 461110 115072 461116
rect 112444 459060 112496 459066
rect 112444 459002 112496 459008
rect 117240 458114 117268 461230
rect 117228 458108 117280 458114
rect 117228 458050 117280 458056
rect 109866 458008 109922 458017
rect 109866 457943 109922 457952
rect 120000 457881 120028 461230
rect 122760 460873 122788 461230
rect 122746 460864 122802 460873
rect 122746 460799 122802 460808
rect 125336 458046 125364 461230
rect 127912 460737 127940 461230
rect 127898 460728 127954 460737
rect 127898 460663 127954 460672
rect 125324 458040 125376 458046
rect 125324 457982 125376 457988
rect 130488 457978 130516 461230
rect 133064 458833 133092 461230
rect 135640 459542 135668 461230
rect 137894 461122 137922 461244
rect 137894 461094 137968 461122
rect 135628 459536 135680 459542
rect 135628 459478 135680 459484
rect 135718 458960 135774 458969
rect 135718 458895 135720 458904
rect 135772 458895 135774 458904
rect 136546 458960 136602 458969
rect 136546 458895 136602 458904
rect 135720 458866 135772 458872
rect 133050 458824 133106 458833
rect 133050 458759 133106 458768
rect 130476 457972 130528 457978
rect 130476 457914 130528 457920
rect 119986 457872 120042 457881
rect 119986 457807 120042 457816
rect 75920 454708 75972 454714
rect 75920 454650 75972 454656
rect 136560 413953 136588 458895
rect 137940 458289 137968 461094
rect 137926 458280 137982 458289
rect 137926 458215 137982 458224
rect 138308 458017 138336 583170
rect 138400 459542 138428 585142
rect 138480 583024 138532 583030
rect 138480 582966 138532 582972
rect 138388 459536 138440 459542
rect 138388 459478 138440 459484
rect 138294 458008 138350 458017
rect 138294 457943 138350 457952
rect 136546 413944 136602 413953
rect 136546 413879 136602 413888
rect 71044 413296 71096 413302
rect 71044 413238 71096 413244
rect 24214 333976 24270 333985
rect 24270 333934 24564 333962
rect 24214 333911 24270 333920
rect 21652 333254 21988 333282
rect 26804 333254 27140 333282
rect 29380 333254 29716 333282
rect 31956 333254 32292 333282
rect 34532 333254 34868 333282
rect 37292 333254 37444 333282
rect 39684 333254 40020 333282
rect 42260 333254 42596 333282
rect 44836 333254 45172 333282
rect 47412 333254 47748 333282
rect 49988 333254 50324 333282
rect 52564 333254 52900 333282
rect 55324 333254 55476 333282
rect 57716 333266 58052 333282
rect 57704 333260 58052 333266
rect 21652 332586 21680 333254
rect 21640 332580 21692 332586
rect 21640 332522 21692 332528
rect 26804 332382 26832 333254
rect 26792 332376 26844 332382
rect 27528 332376 27580 332382
rect 26792 332318 26844 332324
rect 27526 332344 27528 332353
rect 27580 332344 27582 332353
rect 27526 332279 27582 332288
rect 21454 332208 21510 332217
rect 29380 332178 29408 333254
rect 31114 332480 31170 332489
rect 31114 332415 31170 332424
rect 31128 332217 31156 332415
rect 31956 332246 31984 333254
rect 34532 332314 34560 333254
rect 37292 332450 37320 333254
rect 39684 332518 39712 333254
rect 39672 332512 39724 332518
rect 39672 332454 39724 332460
rect 37280 332444 37332 332450
rect 37280 332386 37332 332392
rect 34520 332308 34572 332314
rect 34520 332250 34572 332256
rect 31944 332240 31996 332246
rect 31114 332208 31170 332217
rect 21454 332143 21510 332152
rect 29368 332172 29420 332178
rect 21468 331401 21496 332143
rect 31944 332182 31996 332188
rect 31114 332143 31170 332152
rect 29368 332114 29420 332120
rect 42260 332110 42288 333254
rect 44836 332382 44864 333254
rect 47412 332926 47440 333254
rect 47400 332920 47452 332926
rect 47400 332862 47452 332868
rect 49988 332858 50016 333254
rect 49976 332852 50028 332858
rect 49976 332794 50028 332800
rect 44824 332376 44876 332382
rect 52564 332353 52592 333254
rect 55324 332489 55352 333254
rect 57756 333254 58052 333260
rect 60292 333254 60628 333282
rect 62868 333254 63204 333282
rect 65444 333254 65780 333282
rect 68356 333254 68692 333282
rect 70932 333254 71084 333282
rect 57704 333202 57756 333208
rect 55310 332480 55366 332489
rect 55310 332415 55366 332424
rect 44824 332318 44876 332324
rect 52550 332344 52606 332353
rect 52550 332279 52606 332288
rect 42248 332104 42300 332110
rect 42248 332046 42300 332052
rect 21454 331392 21510 331401
rect 21454 331327 21510 331336
rect 21362 331256 21418 331265
rect 21362 331191 21418 331200
rect 60292 329662 60320 333254
rect 62868 329798 62896 333254
rect 62856 329792 62908 329798
rect 62856 329734 62908 329740
rect 65444 329730 65472 333254
rect 68664 332586 68692 333254
rect 71056 332586 71084 333254
rect 73172 333254 73508 333282
rect 75932 333254 76084 333282
rect 78324 333254 78660 333282
rect 81236 333254 81388 333282
rect 83812 333254 84056 333282
rect 86388 333254 86724 333282
rect 88964 333254 89300 333282
rect 91540 333254 91876 333282
rect 94116 333254 94452 333282
rect 96692 333254 97028 333282
rect 73172 332790 73200 333254
rect 73160 332784 73212 332790
rect 73160 332726 73212 332732
rect 75932 332722 75960 333254
rect 75920 332716 75972 332722
rect 75920 332658 75972 332664
rect 78324 332654 78352 333254
rect 78312 332648 78364 332654
rect 78312 332590 78364 332596
rect 68652 332580 68704 332586
rect 68652 332522 68704 332528
rect 71044 332580 71096 332586
rect 71044 332522 71096 332528
rect 65432 329724 65484 329730
rect 65432 329666 65484 329672
rect 60280 329656 60332 329662
rect 60280 329598 60332 329604
rect 71056 284986 71084 332522
rect 81360 329118 81388 333254
rect 84028 329798 84056 333254
rect 84016 329792 84068 329798
rect 84016 329734 84068 329740
rect 86696 329186 86724 333254
rect 89272 331294 89300 333254
rect 91848 332926 91876 333254
rect 91836 332920 91888 332926
rect 91836 332862 91888 332868
rect 94424 332586 94452 333254
rect 97000 333062 97028 333254
rect 99208 333254 99268 333282
rect 101844 333254 102088 333282
rect 104420 333254 104756 333282
rect 106996 333254 107332 333282
rect 109572 333254 109908 333282
rect 112148 333254 112484 333282
rect 114724 333254 115060 333282
rect 96988 333056 97040 333062
rect 96988 332998 97040 333004
rect 96526 332616 96582 332625
rect 94412 332580 94464 332586
rect 96526 332551 96528 332560
rect 94412 332522 94464 332528
rect 96580 332551 96582 332560
rect 96528 332522 96580 332528
rect 99208 331809 99236 333254
rect 99194 331800 99250 331809
rect 99194 331735 99250 331744
rect 89260 331288 89312 331294
rect 89260 331230 89312 331236
rect 91008 331288 91060 331294
rect 91008 331230 91060 331236
rect 102060 331242 102088 333254
rect 104728 332654 104756 333254
rect 107304 332790 107332 333254
rect 107292 332784 107344 332790
rect 107292 332726 107344 332732
rect 109880 332722 109908 333254
rect 112456 332858 112484 333254
rect 115032 332994 115060 333254
rect 117240 333254 117300 333282
rect 119876 333254 120028 333282
rect 122452 333254 122696 333282
rect 125028 333254 125364 333282
rect 127604 333254 127940 333282
rect 130180 333254 130516 333282
rect 132756 333254 133092 333282
rect 135332 333254 135668 333282
rect 115020 332988 115072 332994
rect 115020 332930 115072 332936
rect 112444 332852 112496 332858
rect 112444 332794 112496 332800
rect 109868 332716 109920 332722
rect 109868 332658 109920 332664
rect 104716 332648 104768 332654
rect 104716 332590 104768 332596
rect 117240 332178 117268 333254
rect 120000 332518 120028 333254
rect 119988 332512 120040 332518
rect 119988 332454 120040 332460
rect 122668 332450 122696 333254
rect 122656 332444 122708 332450
rect 122656 332386 122708 332392
rect 125336 332382 125364 333254
rect 125324 332376 125376 332382
rect 125324 332318 125376 332324
rect 127912 332314 127940 333254
rect 127900 332308 127952 332314
rect 127900 332250 127952 332256
rect 130488 332246 130516 333254
rect 130476 332240 130528 332246
rect 130476 332182 130528 332188
rect 117228 332172 117280 332178
rect 117228 332114 117280 332120
rect 133064 331945 133092 333254
rect 135640 332586 135668 333254
rect 136652 333254 137908 333282
rect 135628 332580 135680 332586
rect 135628 332522 135680 332528
rect 133050 331936 133106 331945
rect 133050 331871 133106 331880
rect 91020 329254 91048 331230
rect 102060 331214 102180 331242
rect 102152 329730 102180 331214
rect 102140 329724 102192 329730
rect 102140 329666 102192 329672
rect 91008 329248 91060 329254
rect 91008 329190 91060 329196
rect 86684 329180 86736 329186
rect 86684 329122 86736 329128
rect 81348 329112 81400 329118
rect 81348 329054 81400 329060
rect 136652 285054 136680 333254
rect 138296 332648 138348 332654
rect 138296 332590 138348 332596
rect 136640 285048 136692 285054
rect 136640 284990 136692 284996
rect 71044 284980 71096 284986
rect 71044 284922 71096 284928
rect 21284 229066 21496 229094
rect 21192 209746 21404 209774
rect 21086 202872 21142 202881
rect 21086 202807 21142 202816
rect 21100 200114 21128 202807
rect 21376 202745 21404 209746
rect 21468 204134 21496 229066
rect 21652 205278 21988 205306
rect 24228 205278 24564 205306
rect 26804 205278 27140 205306
rect 29380 205278 29716 205306
rect 31956 205278 32292 205306
rect 34532 205278 34868 205306
rect 37292 205278 37444 205306
rect 39684 205278 40020 205306
rect 42260 205278 42596 205306
rect 44836 205278 45172 205306
rect 47412 205278 47748 205306
rect 49988 205278 50324 205306
rect 52564 205278 52900 205306
rect 55324 205278 55476 205306
rect 57992 205278 58052 205306
rect 60292 205278 60628 205306
rect 62868 205278 63204 205306
rect 65444 205278 65780 205306
rect 68356 205278 68692 205306
rect 21652 204270 21680 205278
rect 21640 204264 21692 204270
rect 22008 204264 22060 204270
rect 21640 204206 21692 204212
rect 22006 204232 22008 204241
rect 22060 204232 22062 204241
rect 22006 204167 22062 204176
rect 21456 204128 21508 204134
rect 24228 204105 24256 205278
rect 26804 204134 26832 205278
rect 26792 204128 26844 204134
rect 21456 204070 21508 204076
rect 24214 204096 24270 204105
rect 21362 202736 21418 202745
rect 21362 202671 21418 202680
rect 21100 200086 21312 200114
rect 21284 74186 21312 200086
rect 21376 74497 21404 202671
rect 21468 74526 21496 204070
rect 26792 204070 26844 204076
rect 24214 204031 24270 204040
rect 23296 202836 23348 202842
rect 23296 202778 23348 202784
rect 23308 202337 23336 202778
rect 29380 202609 29408 205278
rect 31956 204406 31984 205278
rect 34532 204513 34560 205278
rect 34518 204504 34574 204513
rect 34518 204439 34574 204448
rect 31944 204400 31996 204406
rect 37292 204377 37320 205278
rect 31944 204342 31996 204348
rect 37278 204368 37334 204377
rect 39684 204338 39712 205278
rect 37278 204303 37334 204312
rect 39672 204332 39724 204338
rect 39672 204274 39724 204280
rect 30944 204202 31156 204218
rect 30932 204196 31168 204202
rect 30984 204190 31116 204196
rect 30932 204138 30984 204144
rect 31116 204138 31168 204144
rect 42260 202842 42288 205278
rect 44836 203969 44864 205278
rect 44822 203960 44878 203969
rect 47412 203930 47440 205278
rect 49988 203998 50016 205278
rect 49976 203992 50028 203998
rect 49976 203934 50028 203940
rect 44822 203895 44878 203904
rect 47400 203924 47452 203930
rect 47400 203866 47452 203872
rect 42248 202836 42300 202842
rect 42248 202778 42300 202784
rect 52564 202745 52592 205278
rect 55324 202881 55352 205278
rect 57992 204066 58020 205278
rect 60292 204202 60320 205278
rect 62868 204241 62896 205278
rect 62854 204232 62910 204241
rect 60280 204196 60332 204202
rect 62854 204167 62910 204176
rect 60280 204138 60332 204144
rect 65444 204134 65472 205278
rect 68664 204270 68692 205278
rect 70596 205278 70932 205306
rect 73172 205278 73508 205306
rect 75932 205278 76084 205306
rect 77312 205278 78660 205306
rect 81236 205278 81388 205306
rect 83812 205278 84056 205306
rect 86388 205278 86724 205306
rect 88964 205278 89300 205306
rect 91540 205278 91876 205306
rect 94116 205278 94452 205306
rect 96692 205278 97028 205306
rect 70596 204270 70624 205278
rect 68652 204264 68704 204270
rect 68652 204206 68704 204212
rect 70584 204264 70636 204270
rect 70584 204206 70636 204212
rect 71044 204264 71096 204270
rect 71044 204206 71096 204212
rect 65432 204128 65484 204134
rect 65432 204070 65484 204076
rect 57980 204060 58032 204066
rect 57980 204002 58032 204008
rect 55310 202872 55366 202881
rect 55310 202807 55366 202816
rect 52550 202736 52606 202745
rect 52550 202671 52606 202680
rect 29366 202600 29422 202609
rect 29366 202535 29422 202544
rect 23294 202328 23350 202337
rect 23294 202263 23350 202272
rect 71056 158030 71084 204206
rect 73172 203862 73200 205278
rect 73160 203856 73212 203862
rect 73160 203798 73212 203804
rect 75932 200122 75960 205278
rect 75920 200116 75972 200122
rect 75920 200058 75972 200064
rect 77312 199442 77340 205278
rect 81360 203930 81388 205278
rect 84028 204202 84056 205278
rect 86696 204678 86724 205278
rect 86684 204672 86736 204678
rect 86684 204614 86736 204620
rect 84016 204196 84068 204202
rect 84016 204138 84068 204144
rect 89272 204134 89300 205278
rect 89260 204128 89312 204134
rect 89260 204070 89312 204076
rect 91848 204066 91876 205278
rect 94424 204406 94452 205278
rect 97000 204474 97028 205278
rect 99208 205278 99268 205306
rect 101844 205278 102088 205306
rect 104420 205278 104756 205306
rect 106996 205278 107332 205306
rect 109572 205278 109908 205306
rect 112148 205278 112484 205306
rect 114724 205278 115060 205306
rect 96988 204468 97040 204474
rect 96988 204410 97040 204416
rect 94412 204400 94464 204406
rect 94412 204342 94464 204348
rect 91836 204060 91888 204066
rect 91836 204002 91888 204008
rect 81348 203924 81400 203930
rect 81348 203866 81400 203872
rect 99208 203658 99236 205278
rect 102060 204542 102088 205278
rect 102048 204536 102100 204542
rect 102048 204478 102100 204484
rect 99196 203652 99248 203658
rect 99196 203594 99248 203600
rect 104728 202881 104756 205278
rect 104714 202872 104770 202881
rect 107304 202842 107332 205278
rect 104714 202807 104770 202816
rect 107292 202836 107344 202842
rect 107292 202778 107344 202784
rect 109880 202745 109908 205278
rect 112456 203998 112484 205278
rect 115032 204610 115060 205278
rect 117240 205278 117300 205306
rect 119876 205278 120028 205306
rect 122452 205278 122604 205306
rect 125028 205278 125364 205306
rect 127604 205278 127940 205306
rect 130180 205278 130516 205306
rect 132756 205278 133092 205306
rect 135332 205278 135668 205306
rect 115020 204604 115072 204610
rect 115020 204546 115072 204552
rect 112444 203992 112496 203998
rect 112444 203934 112496 203940
rect 117240 203454 117268 205278
rect 120000 204377 120028 205278
rect 119986 204368 120042 204377
rect 119986 204303 120042 204312
rect 117228 203448 117280 203454
rect 117228 203390 117280 203396
rect 119988 203448 120040 203454
rect 119988 203390 120040 203396
rect 109866 202736 109922 202745
rect 109866 202671 109922 202680
rect 120000 202609 120028 203390
rect 122576 203386 122604 205278
rect 125336 203522 125364 205278
rect 127912 204270 127940 205278
rect 130488 204270 130516 205278
rect 127900 204264 127952 204270
rect 127900 204206 127952 204212
rect 130016 204264 130068 204270
rect 130016 204206 130068 204212
rect 130476 204264 130528 204270
rect 130476 204206 130528 204212
rect 130028 203561 130056 204206
rect 133064 203590 133092 205278
rect 133788 204264 133840 204270
rect 135640 204241 135668 205278
rect 136652 205278 137908 205306
rect 133788 204206 133840 204212
rect 135626 204232 135682 204241
rect 133800 204105 133828 204206
rect 135626 204167 135682 204176
rect 133786 204096 133842 204105
rect 133786 204031 133842 204040
rect 133052 203584 133104 203590
rect 130014 203552 130070 203561
rect 125324 203516 125376 203522
rect 125324 203458 125376 203464
rect 128268 203516 128320 203522
rect 133052 203526 133104 203532
rect 130014 203487 130070 203496
rect 128268 203458 128320 203464
rect 122564 203380 122616 203386
rect 122564 203322 122616 203328
rect 125508 203380 125560 203386
rect 125508 203322 125560 203328
rect 125520 202774 125548 203322
rect 125508 202768 125560 202774
rect 125508 202710 125560 202716
rect 119986 202600 120042 202609
rect 119986 202535 120042 202544
rect 128280 202162 128308 203458
rect 128268 202156 128320 202162
rect 128268 202098 128320 202104
rect 77300 199436 77352 199442
rect 77300 199378 77352 199384
rect 136652 158098 136680 205278
rect 138020 204332 138072 204338
rect 138020 204274 138072 204280
rect 138032 204134 138060 204274
rect 138020 204128 138072 204134
rect 138020 204070 138072 204076
rect 138308 202881 138336 332590
rect 138400 332586 138428 459478
rect 138492 458153 138520 582966
rect 138584 460934 138612 585822
rect 138676 480254 138704 585958
rect 139400 585948 139452 585954
rect 139400 585890 139452 585896
rect 138676 480226 138888 480254
rect 138584 460906 138796 460934
rect 138584 460873 138612 460906
rect 138570 460864 138626 460873
rect 138570 460799 138626 460808
rect 138478 458144 138534 458153
rect 138478 458079 138534 458088
rect 138492 451274 138520 458079
rect 138492 451246 138612 451274
rect 138584 332654 138612 451246
rect 138572 332648 138624 332654
rect 138572 332590 138624 332596
rect 138388 332580 138440 332586
rect 138388 332522 138440 332528
rect 138400 204241 138428 332522
rect 138768 332450 138796 460906
rect 138860 460737 138888 480226
rect 138846 460728 138902 460737
rect 138846 460663 138902 460672
rect 138756 332444 138808 332450
rect 138756 332386 138808 332392
rect 138768 331294 138796 332386
rect 138860 332314 138888 460663
rect 139412 458046 139440 585890
rect 139504 480254 139532 586026
rect 139674 585848 139730 585857
rect 139674 585783 139730 585792
rect 139860 585812 139912 585818
rect 139504 480226 139624 480254
rect 139400 458040 139452 458046
rect 139400 457982 139452 457988
rect 139412 456890 139440 457982
rect 139596 457978 139624 480226
rect 139688 458114 139716 585783
rect 139860 585754 139912 585760
rect 139768 583092 139820 583098
rect 139768 583034 139820 583040
rect 139780 458182 139808 583034
rect 139768 458176 139820 458182
rect 139768 458118 139820 458124
rect 139676 458108 139728 458114
rect 139676 458050 139728 458056
rect 139584 457972 139636 457978
rect 139584 457914 139636 457920
rect 139596 457042 139624 457914
rect 139688 457162 139716 458050
rect 139676 457156 139728 457162
rect 139676 457098 139728 457104
rect 139596 457014 139716 457042
rect 139400 456884 139452 456890
rect 139400 456826 139452 456832
rect 139584 456816 139636 456822
rect 139584 456758 139636 456764
rect 139596 335354 139624 456758
rect 139412 335326 139624 335354
rect 139308 332784 139360 332790
rect 139412 332738 139440 335326
rect 139360 332732 139440 332738
rect 139308 332726 139440 332732
rect 139320 332710 139440 332726
rect 138848 332308 138900 332314
rect 138848 332250 138900 332256
rect 138756 331288 138808 331294
rect 138756 331230 138808 331236
rect 138860 331106 138888 332250
rect 139412 331242 139440 332710
rect 139688 332246 139716 457014
rect 139780 456822 139808 458118
rect 139872 457881 139900 585754
rect 140780 583296 140832 583302
rect 140780 583238 140832 583244
rect 140792 461174 140820 583238
rect 142160 583160 142212 583166
rect 142160 583102 142212 583108
rect 140964 542088 141016 542094
rect 140964 542030 141016 542036
rect 140872 541884 140924 541890
rect 140872 541826 140924 541832
rect 140780 461168 140832 461174
rect 140780 461110 140832 461116
rect 139858 457872 139914 457881
rect 139858 457807 139914 457816
rect 139768 456816 139820 456822
rect 139768 456758 139820 456764
rect 139872 451274 139900 457807
rect 139952 457156 140004 457162
rect 139952 457098 140004 457104
rect 139780 451246 139900 451274
rect 139780 332518 139808 451246
rect 139768 332512 139820 332518
rect 139768 332454 139820 332460
rect 139676 332240 139728 332246
rect 139676 332182 139728 332188
rect 139492 331628 139544 331634
rect 139492 331570 139544 331576
rect 138584 331078 138888 331106
rect 139320 331214 139440 331242
rect 138584 316034 138612 331078
rect 138662 329760 138718 329769
rect 138662 329695 138718 329704
rect 138676 329254 138704 329695
rect 138664 329248 138716 329254
rect 138664 329190 138716 329196
rect 138492 316006 138612 316034
rect 138386 204232 138442 204241
rect 138386 204167 138442 204176
rect 138492 204082 138520 316006
rect 138676 204338 138704 329190
rect 138664 204332 138716 204338
rect 138664 204274 138716 204280
rect 138570 204232 138626 204241
rect 138570 204167 138626 204176
rect 138400 204054 138520 204082
rect 138400 203561 138428 204054
rect 138386 203552 138442 203561
rect 138386 203487 138442 203496
rect 138294 202872 138350 202881
rect 138020 202836 138072 202842
rect 138294 202807 138350 202816
rect 138020 202778 138072 202784
rect 138032 202706 138060 202778
rect 138020 202700 138072 202706
rect 138020 202642 138072 202648
rect 136640 158092 136692 158098
rect 136640 158034 136692 158040
rect 71044 158024 71096 158030
rect 71044 157966 71096 157972
rect 135628 78668 135680 78674
rect 135628 78610 135680 78616
rect 135640 78554 135668 78610
rect 135272 78526 135668 78554
rect 129752 77994 130516 78010
rect 129752 77988 130528 77994
rect 129752 77982 130476 77988
rect 68652 77376 68704 77382
rect 21652 77302 21988 77330
rect 24228 77302 24564 77330
rect 21652 75721 21680 77302
rect 24228 75857 24256 77302
rect 27126 77058 27154 77316
rect 29656 77302 29716 77330
rect 32292 77302 32444 77330
rect 27126 77030 27200 77058
rect 24214 75848 24270 75857
rect 24214 75783 24270 75792
rect 21638 75712 21694 75721
rect 21638 75647 21694 75656
rect 27172 74526 27200 77030
rect 21456 74520 21508 74526
rect 21362 74488 21418 74497
rect 21456 74462 21508 74468
rect 27160 74520 27212 74526
rect 27160 74462 27212 74468
rect 21362 74423 21418 74432
rect 21272 74180 21324 74186
rect 21272 74122 21324 74128
rect 27172 71058 27200 74462
rect 29656 74254 29684 77302
rect 32416 74322 32444 77302
rect 34532 77302 34868 77330
rect 34532 75886 34560 77302
rect 37430 77058 37458 77316
rect 39960 77302 40020 77330
rect 42076 77302 42596 77330
rect 44836 77302 45172 77330
rect 47596 77302 47748 77330
rect 37430 77030 37504 77058
rect 34520 75880 34572 75886
rect 34520 75822 34572 75828
rect 34532 75206 34560 75822
rect 34520 75200 34572 75206
rect 34520 75142 34572 75148
rect 37476 74390 37504 77030
rect 37464 74384 37516 74390
rect 39960 74361 39988 77302
rect 37464 74326 37516 74332
rect 39946 74352 40002 74361
rect 32404 74316 32456 74322
rect 32404 74258 32456 74264
rect 29644 74248 29696 74254
rect 29644 74190 29696 74196
rect 27160 71052 27212 71058
rect 27160 70994 27212 71000
rect 29656 62830 29684 74190
rect 32416 62898 32444 74258
rect 37476 71126 37504 74326
rect 39946 74287 40002 74296
rect 42076 74225 42104 77302
rect 44836 74458 44864 77302
rect 47596 75546 47624 77302
rect 50310 77058 50338 77316
rect 52900 77302 53052 77330
rect 55476 77302 55904 77330
rect 50310 77030 50384 77058
rect 50356 75614 50384 77030
rect 50344 75608 50396 75614
rect 50344 75550 50396 75556
rect 47584 75540 47636 75546
rect 47584 75482 47636 75488
rect 44824 74452 44876 74458
rect 44824 74394 44876 74400
rect 42062 74216 42118 74225
rect 42062 74151 42118 74160
rect 37464 71120 37516 71126
rect 37464 71062 37516 71068
rect 42076 66910 42104 74151
rect 42064 66904 42116 66910
rect 42064 66846 42116 66852
rect 44836 64190 44864 74394
rect 47596 64258 47624 75482
rect 50356 64326 50384 75550
rect 53024 74497 53052 77302
rect 53010 74488 53066 74497
rect 53010 74423 53066 74432
rect 53024 73953 53052 74423
rect 55876 74186 55904 77302
rect 57992 77302 58052 77330
rect 57992 75682 58020 77302
rect 60614 77058 60642 77316
rect 63190 77058 63218 77316
rect 65536 77302 65780 77330
rect 68356 77324 68652 77330
rect 68356 77318 68704 77324
rect 70584 77376 70636 77382
rect 70636 77324 71268 77330
rect 70584 77318 71268 77324
rect 68356 77302 68692 77318
rect 70596 77302 71268 77318
rect 60614 77030 60688 77058
rect 63190 77030 63264 77058
rect 60660 75750 60688 77030
rect 63236 75818 63264 77030
rect 63224 75812 63276 75818
rect 63224 75754 63276 75760
rect 60648 75744 60700 75750
rect 60648 75686 60700 75692
rect 57980 75676 58032 75682
rect 57980 75618 58032 75624
rect 57992 75410 58020 75618
rect 57980 75404 58032 75410
rect 57980 75346 58032 75352
rect 59268 75404 59320 75410
rect 59268 75346 59320 75352
rect 55864 74180 55916 74186
rect 55864 74122 55916 74128
rect 56508 74180 56560 74186
rect 56508 74122 56560 74128
rect 53010 73944 53066 73953
rect 53010 73879 53066 73888
rect 56520 66978 56548 74122
rect 59280 72486 59308 75346
rect 59268 72480 59320 72486
rect 59268 72422 59320 72428
rect 60660 69698 60688 75686
rect 60648 69692 60700 69698
rect 60648 69634 60700 69640
rect 63236 68338 63264 75754
rect 65536 75721 65564 77302
rect 65522 75712 65578 75721
rect 65522 75647 65578 75656
rect 63224 68332 63276 68338
rect 63224 68274 63276 68280
rect 56508 66972 56560 66978
rect 56508 66914 56560 66920
rect 50344 64320 50396 64326
rect 50344 64262 50396 64268
rect 47584 64252 47636 64258
rect 47584 64194 47636 64200
rect 44824 64184 44876 64190
rect 44824 64126 44876 64132
rect 65536 62966 65564 75647
rect 71240 75274 71268 77302
rect 73494 77058 73522 77316
rect 75932 77302 76084 77330
rect 73494 77030 73568 77058
rect 73540 75478 73568 77030
rect 75932 75954 75960 77302
rect 78646 77110 78674 77316
rect 81236 77302 81388 77330
rect 83812 77302 84056 77330
rect 86388 77302 86724 77330
rect 77300 77104 77352 77110
rect 77300 77046 77352 77052
rect 78634 77104 78686 77110
rect 78634 77046 78686 77052
rect 77312 76022 77340 77046
rect 77300 76016 77352 76022
rect 77300 75958 77352 75964
rect 75920 75948 75972 75954
rect 75920 75890 75972 75896
rect 73528 75472 73580 75478
rect 73528 75414 73580 75420
rect 71228 75268 71280 75274
rect 71228 75210 71280 75216
rect 73540 69902 73568 75414
rect 75932 72690 75960 75890
rect 75920 72684 75972 72690
rect 75920 72626 75972 72632
rect 73528 69896 73580 69902
rect 73528 69838 73580 69844
rect 77312 65521 77340 75958
rect 77944 75268 77996 75274
rect 77944 75210 77996 75216
rect 77956 67046 77984 75210
rect 81360 70378 81388 77302
rect 81348 70372 81400 70378
rect 81348 70314 81400 70320
rect 84028 69018 84056 77302
rect 86696 75177 86724 77302
rect 88352 77302 88964 77330
rect 91540 77302 91876 77330
rect 86682 75168 86738 75177
rect 86682 75103 86738 75112
rect 84016 69012 84068 69018
rect 84016 68954 84068 68960
rect 77944 67040 77996 67046
rect 77944 66982 77996 66988
rect 88352 66230 88380 77302
rect 91848 75886 91876 77302
rect 93872 77302 94116 77330
rect 96632 77302 96692 77330
rect 98380 77302 99268 77330
rect 100772 77302 101844 77330
rect 104420 77302 104664 77330
rect 106996 77302 107332 77330
rect 91836 75880 91888 75886
rect 91836 75822 91888 75828
rect 88340 66224 88392 66230
rect 88340 66166 88392 66172
rect 93872 66162 93900 77302
rect 93860 66156 93912 66162
rect 93860 66098 93912 66104
rect 96632 66094 96660 77302
rect 96620 66088 96672 66094
rect 96620 66030 96672 66036
rect 77298 65512 77354 65521
rect 77298 65447 77354 65456
rect 65524 62960 65576 62966
rect 65524 62902 65576 62908
rect 32404 62892 32456 62898
rect 32404 62834 32456 62840
rect 29644 62824 29696 62830
rect 29644 62766 29696 62772
rect 57060 62076 57112 62082
rect 57060 62018 57112 62024
rect 57072 61577 57100 62018
rect 98380 61742 98408 77302
rect 100024 75200 100076 75206
rect 100024 75142 100076 75148
rect 98368 61736 98420 61742
rect 98368 61678 98420 61684
rect 99286 61704 99342 61713
rect 99286 61639 99342 61648
rect 57058 61568 57114 61577
rect 57058 61503 57114 61512
rect 99300 60625 99328 61639
rect 99286 60616 99342 60625
rect 99286 60551 99342 60560
rect 100036 58682 100064 75142
rect 100772 62082 100800 77302
rect 104636 73166 104664 77302
rect 107304 75818 107332 77302
rect 109052 77302 109572 77330
rect 112148 77302 112484 77330
rect 107292 75812 107344 75818
rect 107292 75754 107344 75760
rect 104624 73160 104676 73166
rect 104624 73102 104676 73108
rect 100760 62076 100812 62082
rect 100760 62018 100812 62024
rect 102874 60752 102930 60761
rect 102874 60687 102930 60696
rect 100024 58676 100076 58682
rect 100024 58618 100076 58624
rect 102782 58032 102838 58041
rect 102782 57967 102838 57976
rect 102598 56672 102654 56681
rect 102598 56607 102654 56616
rect 57520 56568 57572 56574
rect 57520 56510 57572 56516
rect 57532 56409 57560 56510
rect 57518 56400 57574 56409
rect 57518 56335 57574 56344
rect 102138 55584 102194 55593
rect 102138 55519 102194 55528
rect 102152 55282 102180 55519
rect 102140 55276 102192 55282
rect 102140 55218 102192 55224
rect 102138 54360 102194 54369
rect 102138 54295 102194 54304
rect 102152 53922 102180 54295
rect 102140 53916 102192 53922
rect 102140 53858 102192 53864
rect 102230 53136 102286 53145
rect 102230 53071 102286 53080
rect 102138 52592 102194 52601
rect 102138 52527 102140 52536
rect 102192 52527 102194 52536
rect 102140 52498 102192 52504
rect 102244 52494 102272 53071
rect 102232 52488 102284 52494
rect 102232 52430 102284 52436
rect 57060 52420 57112 52426
rect 57060 52362 57112 52368
rect 57072 51785 57100 52362
rect 57058 51776 57114 51785
rect 57058 51711 57114 51720
rect 102138 50144 102194 50153
rect 102138 50079 102194 50088
rect 102152 49842 102180 50079
rect 102140 49836 102192 49842
rect 102140 49778 102192 49784
rect 102612 49638 102640 56607
rect 102796 49706 102824 57967
rect 102888 52426 102916 60687
rect 103150 59664 103206 59673
rect 103150 59599 103206 59608
rect 103058 58576 103114 58585
rect 103058 58511 103114 58520
rect 102876 52420 102928 52426
rect 102876 52362 102928 52368
rect 103072 51066 103100 58511
rect 103164 52358 103192 59599
rect 109052 57934 109080 77302
rect 112456 75750 112484 77302
rect 114572 77302 114724 77330
rect 117240 77302 117300 77330
rect 119876 77302 120028 77330
rect 122452 77302 122604 77330
rect 125028 77302 125364 77330
rect 127604 77302 127940 77330
rect 112444 75744 112496 75750
rect 112444 75686 112496 75692
rect 109040 57928 109092 57934
rect 109040 57870 109092 57876
rect 114572 57866 114600 77302
rect 117240 68950 117268 77302
rect 120000 75546 120028 77302
rect 122576 75682 122604 77302
rect 122564 75676 122616 75682
rect 122564 75618 122616 75624
rect 125336 75614 125364 77302
rect 125324 75608 125376 75614
rect 125324 75550 125376 75556
rect 119988 75540 120040 75546
rect 119988 75482 120040 75488
rect 127912 75478 127940 77302
rect 127900 75472 127952 75478
rect 127900 75414 127952 75420
rect 117228 68944 117280 68950
rect 117228 68886 117280 68892
rect 129752 58818 129780 77982
rect 130476 77930 130528 77936
rect 132756 77302 133092 77330
rect 131120 75540 131172 75546
rect 131120 75482 131172 75488
rect 131132 75177 131160 75482
rect 133064 75342 133092 77302
rect 133052 75336 133104 75342
rect 133052 75278 133104 75284
rect 131118 75168 131174 75177
rect 131118 75103 131174 75112
rect 135272 58886 135300 78526
rect 137894 77058 137922 77316
rect 137894 77030 137968 77058
rect 137940 71194 137968 77030
rect 138308 73166 138336 202807
rect 138400 75478 138428 203487
rect 138480 202836 138532 202842
rect 138480 202778 138532 202784
rect 138492 202162 138520 202778
rect 138480 202156 138532 202162
rect 138480 202098 138532 202104
rect 138492 75614 138520 202098
rect 138584 78674 138612 204167
rect 139320 202706 139348 331214
rect 139504 331106 139532 331570
rect 139584 331288 139636 331294
rect 139584 331230 139636 331236
rect 139412 331078 139532 331106
rect 139308 202700 139360 202706
rect 139308 202642 139360 202648
rect 139412 202609 139440 331078
rect 139492 331016 139544 331022
rect 139492 330958 139544 330964
rect 139504 202842 139532 330958
rect 139492 202836 139544 202842
rect 139492 202778 139544 202784
rect 139596 202774 139624 331230
rect 139688 209774 139716 332182
rect 139780 229094 139808 332454
rect 139964 332178 139992 457098
rect 140044 456884 140096 456890
rect 140044 456826 140096 456832
rect 140056 332382 140084 456826
rect 140792 332994 140820 461110
rect 140884 459338 140912 541826
rect 140976 459406 141004 542030
rect 141056 541748 141108 541754
rect 141056 541690 141108 541696
rect 141068 460970 141096 541690
rect 142066 461000 142122 461009
rect 141056 460964 141108 460970
rect 142066 460935 142068 460944
rect 141056 460906 141108 460912
rect 142120 460935 142122 460944
rect 142068 460906 142120 460912
rect 140964 459400 141016 459406
rect 140964 459342 141016 459348
rect 140872 459332 140924 459338
rect 140872 459274 140924 459280
rect 140884 459082 140912 459274
rect 140976 459218 141004 459342
rect 140976 459190 141280 459218
rect 140884 459054 141004 459082
rect 140872 458992 140924 458998
rect 140872 458934 140924 458940
rect 140884 458794 140912 458934
rect 140872 458788 140924 458794
rect 140872 458730 140924 458736
rect 140976 458674 141004 459054
rect 141148 459060 141200 459066
rect 141148 459002 141200 459008
rect 141056 458788 141108 458794
rect 141056 458730 141108 458736
rect 140884 458646 141004 458674
rect 140780 332988 140832 332994
rect 140780 332930 140832 332936
rect 140884 332926 140912 458646
rect 140964 458244 141016 458250
rect 140964 458186 141016 458192
rect 140872 332920 140924 332926
rect 140872 332862 140924 332868
rect 140044 332376 140096 332382
rect 140044 332318 140096 332324
rect 139952 332172 140004 332178
rect 139952 332114 140004 332120
rect 139964 331634 139992 332114
rect 139952 331628 140004 331634
rect 139952 331570 140004 331576
rect 140056 331022 140084 332318
rect 140044 331016 140096 331022
rect 140044 330958 140096 330964
rect 140780 329180 140832 329186
rect 140780 329122 140832 329128
rect 140792 327758 140820 329122
rect 140780 327752 140832 327758
rect 140780 327694 140832 327700
rect 140780 327616 140832 327622
rect 140780 327558 140832 327564
rect 139780 229066 139900 229094
rect 139688 209746 139808 209774
rect 139780 204105 139808 209746
rect 139872 204377 139900 229066
rect 140792 209774 140820 327558
rect 140884 229094 140912 332862
rect 140976 329730 141004 458186
rect 141068 333062 141096 458730
rect 141056 333056 141108 333062
rect 141056 332998 141108 333004
rect 140964 329724 141016 329730
rect 140964 329666 141016 329672
rect 141068 229094 141096 332998
rect 141160 332858 141188 459002
rect 141252 458250 141280 459190
rect 142172 459066 142200 583102
rect 142436 544400 142488 544406
rect 142436 544342 142488 544348
rect 142252 542020 142304 542026
rect 142252 541962 142304 541968
rect 142160 459060 142212 459066
rect 142160 459002 142212 459008
rect 142264 458794 142292 541962
rect 142344 541952 142396 541958
rect 142344 541894 142396 541900
rect 142356 459474 142384 541894
rect 142448 461106 142476 544342
rect 142528 541816 142580 541822
rect 142528 541758 142580 541764
rect 142436 461100 142488 461106
rect 142436 461042 142488 461048
rect 142540 461038 142568 541758
rect 143540 461100 143592 461106
rect 143540 461042 143592 461048
rect 142528 461032 142580 461038
rect 142528 460974 142580 460980
rect 142344 459468 142396 459474
rect 142344 459410 142396 459416
rect 142252 458788 142304 458794
rect 142252 458730 142304 458736
rect 141240 458244 141292 458250
rect 141240 458186 141292 458192
rect 142250 458008 142306 458017
rect 142250 457943 142306 457952
rect 142160 332988 142212 332994
rect 142160 332930 142212 332936
rect 141148 332852 141200 332858
rect 141148 332794 141200 332800
rect 141160 327622 141188 332794
rect 141514 329760 141570 329769
rect 141514 329695 141570 329704
rect 141528 329118 141556 329695
rect 141516 329112 141568 329118
rect 141516 329054 141568 329060
rect 141148 327616 141200 327622
rect 141148 327558 141200 327564
rect 140884 229066 141004 229094
rect 141068 229066 141188 229094
rect 140976 209774 141004 229066
rect 140792 209746 140912 209774
rect 140976 209746 141096 209774
rect 140780 206372 140832 206378
rect 140780 206314 140832 206320
rect 140792 204678 140820 206314
rect 140780 204672 140832 204678
rect 140780 204614 140832 204620
rect 139858 204368 139914 204377
rect 139858 204303 139914 204312
rect 139766 204096 139822 204105
rect 139766 204031 139822 204040
rect 139584 202768 139636 202774
rect 139584 202710 139636 202716
rect 139398 202600 139454 202609
rect 139398 202535 139454 202544
rect 138572 78668 138624 78674
rect 138572 78610 138624 78616
rect 138480 75608 138532 75614
rect 138480 75550 138532 75556
rect 138388 75472 138440 75478
rect 138388 75414 138440 75420
rect 138400 73846 138428 75414
rect 138388 73840 138440 73846
rect 138388 73782 138440 73788
rect 138296 73160 138348 73166
rect 138296 73102 138348 73108
rect 138308 72758 138336 73102
rect 138296 72752 138348 72758
rect 138296 72694 138348 72700
rect 137928 71188 137980 71194
rect 137928 71130 137980 71136
rect 138492 68474 138520 75550
rect 139412 68950 139440 202535
rect 139492 75812 139544 75818
rect 139492 75754 139544 75760
rect 139504 75206 139532 75754
rect 139596 75682 139624 202710
rect 139676 202700 139728 202706
rect 139676 202642 139728 202648
rect 139688 75818 139716 202642
rect 139780 77994 139808 204031
rect 139768 77988 139820 77994
rect 139768 77930 139820 77936
rect 139676 75812 139728 75818
rect 139676 75754 139728 75760
rect 139584 75676 139636 75682
rect 139584 75618 139636 75624
rect 139492 75200 139544 75206
rect 139492 75142 139544 75148
rect 139596 72554 139624 75618
rect 139872 75177 139900 204303
rect 140884 203998 140912 209746
rect 141068 204066 141096 209746
rect 141160 204474 141188 229066
rect 141240 205624 141292 205630
rect 141240 205566 141292 205572
rect 141252 204542 141280 205566
rect 141240 204536 141292 204542
rect 141240 204478 141292 204484
rect 141148 204468 141200 204474
rect 141148 204410 141200 204416
rect 141056 204060 141108 204066
rect 141056 204002 141108 204008
rect 140872 203992 140924 203998
rect 140872 203934 140924 203940
rect 140884 200114 140912 203934
rect 140884 200086 141004 200114
rect 140976 84194 141004 200086
rect 140884 84166 141004 84194
rect 140780 75880 140832 75886
rect 140780 75822 140832 75828
rect 140792 75410 140820 75822
rect 140884 75750 140912 84166
rect 141068 75886 141096 204002
rect 141056 75880 141108 75886
rect 141056 75822 141108 75828
rect 140872 75744 140924 75750
rect 140872 75686 140924 75692
rect 140780 75404 140832 75410
rect 140780 75346 140832 75352
rect 140884 75274 140912 75686
rect 140872 75268 140924 75274
rect 140872 75210 140924 75216
rect 139858 75168 139914 75177
rect 139858 75103 139914 75112
rect 139584 72548 139636 72554
rect 139584 72490 139636 72496
rect 139872 69766 139900 75103
rect 141160 74534 141188 204410
rect 141252 203402 141280 204478
rect 141528 203930 141556 329054
rect 142068 327752 142120 327758
rect 142068 327694 142120 327700
rect 142080 206378 142108 327694
rect 142068 206372 142120 206378
rect 142068 206314 142120 206320
rect 142172 204610 142200 332930
rect 142264 332722 142292 457943
rect 142252 332716 142304 332722
rect 142252 332658 142304 332664
rect 142160 204604 142212 204610
rect 142160 204546 142212 204552
rect 141516 203924 141568 203930
rect 141516 203866 141568 203872
rect 141252 203374 141464 203402
rect 141240 203312 141292 203318
rect 141240 203254 141292 203260
rect 141068 74506 141188 74534
rect 139860 69760 139912 69766
rect 139860 69702 139912 69708
rect 139400 68944 139452 68950
rect 139400 68886 139452 68892
rect 138480 68468 138532 68474
rect 138480 68410 138532 68416
rect 139412 68406 139440 68886
rect 139400 68400 139452 68406
rect 139400 68342 139452 68348
rect 141068 66094 141096 74506
rect 141252 71618 141280 203254
rect 141160 71590 141280 71618
rect 141160 70378 141188 71590
rect 141148 70372 141200 70378
rect 141148 70314 141200 70320
rect 141160 69970 141188 70314
rect 141148 69964 141200 69970
rect 141148 69906 141200 69912
rect 140780 66088 140832 66094
rect 140780 66030 140832 66036
rect 141056 66088 141108 66094
rect 141056 66030 141108 66036
rect 140792 65550 140820 66030
rect 140780 65544 140832 65550
rect 140780 65486 140832 65492
rect 140780 62076 140832 62082
rect 140780 62018 140832 62024
rect 140792 61470 140820 62018
rect 141436 61470 141464 203374
rect 141528 203318 141556 203866
rect 141516 203312 141568 203318
rect 141516 203254 141568 203260
rect 140780 61464 140832 61470
rect 140780 61406 140832 61412
rect 141424 61464 141476 61470
rect 141424 61406 141476 61412
rect 135260 58880 135312 58886
rect 135260 58822 135312 58828
rect 129740 58812 129792 58818
rect 129740 58754 129792 58760
rect 142172 57866 142200 204546
rect 142264 202745 142292 332658
rect 142356 332625 142384 459410
rect 142540 335354 142568 460974
rect 142448 335326 142568 335354
rect 142342 332616 142398 332625
rect 142342 332551 142398 332560
rect 142356 204406 142384 332551
rect 142448 329798 142476 335326
rect 142436 329792 142488 329798
rect 142436 329734 142488 329740
rect 142344 204400 142396 204406
rect 142344 204342 142396 204348
rect 142250 202736 142306 202745
rect 142250 202671 142306 202680
rect 142264 57934 142292 202671
rect 142356 66162 142384 204342
rect 142448 204202 142476 329734
rect 142528 329724 142580 329730
rect 142528 329666 142580 329672
rect 142540 205630 142568 329666
rect 143552 327758 143580 461042
rect 143540 327752 143592 327758
rect 143540 327694 143592 327700
rect 143540 206372 143592 206378
rect 143540 206314 143592 206320
rect 142528 205624 142580 205630
rect 142528 205566 142580 205572
rect 142436 204196 142488 204202
rect 142436 204138 142488 204144
rect 142448 69018 142476 204138
rect 142436 69012 142488 69018
rect 142436 68954 142488 68960
rect 143448 69012 143500 69018
rect 143448 68954 143500 68960
rect 143460 68542 143488 68954
rect 143448 68536 143500 68542
rect 143448 68478 143500 68484
rect 142344 66156 142396 66162
rect 142344 66098 142396 66104
rect 143448 66156 143500 66162
rect 143448 66098 143500 66104
rect 143460 65618 143488 66098
rect 143448 65612 143500 65618
rect 143448 65554 143500 65560
rect 143552 60625 143580 206314
rect 143632 204332 143684 204338
rect 143632 204274 143684 204280
rect 143644 66230 143672 204274
rect 143632 66224 143684 66230
rect 143632 66166 143684 66172
rect 144828 66224 144880 66230
rect 144828 66166 144880 66172
rect 144840 65754 144868 66166
rect 144828 65748 144880 65754
rect 144828 65690 144880 65696
rect 143538 60616 143594 60625
rect 143538 60551 143594 60560
rect 144826 60616 144882 60625
rect 144826 60551 144882 60560
rect 144840 59945 144868 60551
rect 144826 59936 144882 59945
rect 144826 59871 144882 59880
rect 142252 57928 142304 57934
rect 142252 57870 142304 57876
rect 143448 57928 143500 57934
rect 143448 57870 143500 57876
rect 114560 57860 114612 57866
rect 114560 57802 114612 57808
rect 142160 57860 142212 57866
rect 142160 57802 142212 57808
rect 143356 57860 143408 57866
rect 143356 57802 143408 57808
rect 143368 57254 143396 57802
rect 143460 57322 143488 57870
rect 143448 57316 143500 57322
rect 143448 57258 143500 57264
rect 143356 57248 143408 57254
rect 143356 57190 143408 57196
rect 196624 55276 196676 55282
rect 196624 55218 196676 55224
rect 103888 53916 103940 53922
rect 103888 53858 103940 53864
rect 103152 52352 103204 52358
rect 103152 52294 103204 52300
rect 103242 51096 103298 51105
rect 103060 51060 103112 51066
rect 103242 51031 103298 51040
rect 103060 51002 103112 51008
rect 102784 49700 102836 49706
rect 102784 49642 102836 49648
rect 102600 49632 102652 49638
rect 102600 49574 102652 49580
rect 102874 48784 102930 48793
rect 102874 48719 102930 48728
rect 102598 47016 102654 47025
rect 102598 46951 102654 46960
rect 57520 46912 57572 46918
rect 57518 46880 57520 46889
rect 57572 46880 57574 46889
rect 57518 46815 57574 46824
rect 60004 44192 60056 44198
rect 60004 44134 60056 44140
rect 57152 42764 57204 42770
rect 57152 42706 57204 42712
rect 57164 42129 57192 42706
rect 57150 42120 57206 42129
rect 57150 42055 57206 42064
rect 57060 37256 57112 37262
rect 57060 37198 57112 37204
rect 57072 36961 57100 37198
rect 57058 36952 57114 36961
rect 57058 36887 57114 36896
rect 57612 31748 57664 31754
rect 57612 31690 57664 31696
rect 57624 31657 57652 31690
rect 57610 31648 57666 31657
rect 57610 31583 57666 31592
rect 57244 27600 57296 27606
rect 57244 27542 57296 27548
rect 57256 27169 57284 27542
rect 57242 27160 57298 27169
rect 57242 27095 57298 27104
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 60016 22302 60044 44134
rect 102322 43344 102378 43353
rect 102322 43279 102378 43288
rect 102138 42936 102194 42945
rect 102138 42871 102194 42880
rect 102152 40730 102180 42871
rect 102230 41440 102286 41449
rect 102230 41375 102286 41384
rect 102140 40724 102192 40730
rect 102140 40666 102192 40672
rect 102138 40080 102194 40089
rect 102138 40015 102194 40024
rect 102152 37262 102180 40015
rect 102244 38622 102272 41375
rect 102336 40050 102364 43279
rect 102612 42770 102640 46951
rect 102888 44130 102916 48719
rect 102966 47696 103022 47705
rect 102966 47631 103022 47640
rect 102876 44124 102928 44130
rect 102876 44066 102928 44072
rect 102600 42764 102652 42770
rect 102600 42706 102652 42712
rect 102980 42702 103008 47631
rect 103256 45558 103284 51031
rect 103900 48278 103928 53858
rect 196164 52556 196216 52562
rect 196164 52498 196216 52504
rect 103980 52488 104032 52494
rect 103980 52430 104032 52436
rect 103888 48272 103940 48278
rect 103888 48214 103940 48220
rect 103992 46918 104020 52430
rect 195980 52420 196032 52426
rect 195980 52362 196032 52368
rect 195992 52329 196020 52362
rect 196072 52352 196124 52358
rect 195978 52320 196034 52329
rect 196072 52294 196124 52300
rect 195978 52255 196034 52264
rect 196084 51785 196112 52294
rect 196070 51776 196126 51785
rect 196070 51711 196126 51720
rect 195980 51060 196032 51066
rect 195980 51002 196032 51008
rect 195992 50969 196020 51002
rect 195978 50960 196034 50969
rect 195978 50895 196034 50904
rect 104348 49836 104400 49842
rect 104348 49778 104400 49784
rect 103980 46912 104032 46918
rect 103980 46854 104032 46860
rect 103426 45656 103482 45665
rect 103482 45614 103560 45642
rect 103426 45591 103482 45600
rect 103244 45552 103296 45558
rect 103244 45494 103296 45500
rect 102968 42696 103020 42702
rect 102968 42638 103020 42644
rect 103532 41410 103560 45614
rect 103610 44432 103666 44441
rect 103610 44367 103666 44376
rect 103520 41404 103572 41410
rect 103520 41346 103572 41352
rect 102324 40044 102376 40050
rect 102324 39986 102376 39992
rect 103624 39982 103652 44367
rect 104360 44062 104388 49778
rect 195980 49700 196032 49706
rect 195980 49642 196032 49648
rect 195992 49609 196020 49642
rect 196072 49632 196124 49638
rect 195978 49600 196034 49609
rect 196072 49574 196124 49580
rect 195978 49535 196034 49544
rect 196084 49201 196112 49574
rect 196070 49192 196126 49201
rect 196070 49127 196126 49136
rect 195980 48272 196032 48278
rect 195980 48214 196032 48220
rect 195992 47841 196020 48214
rect 195978 47832 196034 47841
rect 195978 47767 196034 47776
rect 195980 46912 196032 46918
rect 195978 46880 195980 46889
rect 196032 46880 196034 46889
rect 195978 46815 196034 46824
rect 196176 46209 196204 52498
rect 196636 48249 196664 55218
rect 196622 48240 196678 48249
rect 196622 48175 196678 48184
rect 196162 46200 196218 46209
rect 196162 46135 196218 46144
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 195992 45257 196020 45494
rect 195978 45248 196034 45257
rect 195978 45183 196034 45192
rect 196072 44124 196124 44130
rect 196072 44066 196124 44072
rect 104348 44056 104400 44062
rect 195980 44056 196032 44062
rect 104348 43998 104400 44004
rect 195978 44024 195980 44033
rect 196032 44024 196034 44033
rect 195978 43959 196034 43968
rect 196084 43625 196112 44066
rect 196070 43616 196126 43625
rect 196070 43551 196126 43560
rect 196072 42764 196124 42770
rect 196072 42706 196124 42712
rect 195980 42696 196032 42702
rect 195980 42638 196032 42644
rect 195992 42537 196020 42638
rect 195978 42528 196034 42537
rect 195978 42463 196034 42472
rect 196084 42129 196112 42706
rect 196070 42120 196126 42129
rect 196070 42055 196126 42064
rect 195980 41404 196032 41410
rect 195980 41346 196032 41352
rect 195992 41177 196020 41346
rect 195978 41168 196034 41177
rect 195978 41103 196034 41112
rect 196164 40724 196216 40730
rect 196164 40666 196216 40672
rect 196072 40044 196124 40050
rect 196072 39986 196124 39992
rect 103612 39976 103664 39982
rect 195980 39976 196032 39982
rect 103612 39918 103664 39924
rect 195978 39944 195980 39953
rect 196032 39944 196034 39953
rect 195978 39879 196034 39888
rect 196084 39545 196112 39986
rect 196070 39536 196126 39545
rect 196070 39471 196126 39480
rect 102782 38992 102838 39001
rect 102782 38927 102838 38936
rect 102232 38616 102284 38622
rect 102232 38558 102284 38564
rect 102598 37904 102654 37913
rect 102598 37839 102654 37848
rect 102140 37256 102192 37262
rect 102140 37198 102192 37204
rect 102612 35834 102640 37839
rect 102690 36136 102746 36145
rect 102690 36071 102746 36080
rect 102600 35828 102652 35834
rect 102600 35770 102652 35776
rect 102138 34640 102194 34649
rect 102138 34575 102194 34584
rect 102152 33114 102180 34575
rect 102704 34474 102732 36071
rect 102796 35902 102824 38927
rect 195980 38616 196032 38622
rect 196176 38593 196204 40666
rect 195980 38558 196032 38564
rect 196162 38584 196218 38593
rect 195992 38049 196020 38558
rect 196162 38519 196218 38528
rect 195978 38040 196034 38049
rect 195978 37975 196034 37984
rect 102874 37360 102930 37369
rect 102874 37295 102930 37304
rect 102784 35896 102836 35902
rect 102784 35838 102836 35844
rect 102692 34468 102744 34474
rect 102692 34410 102744 34416
rect 102888 34406 102916 37295
rect 195980 37256 196032 37262
rect 195980 37198 196032 37204
rect 195992 37097 196020 37198
rect 195978 37088 196034 37097
rect 195978 37023 196034 37032
rect 195980 35896 196032 35902
rect 195978 35864 195980 35873
rect 196032 35864 196034 35873
rect 195978 35799 196034 35808
rect 196072 35828 196124 35834
rect 196072 35770 196124 35776
rect 196084 35465 196112 35770
rect 196070 35456 196126 35465
rect 196070 35391 196126 35400
rect 196072 34468 196124 34474
rect 196072 34410 196124 34416
rect 102876 34400 102928 34406
rect 195980 34400 196032 34406
rect 102876 34342 102928 34348
rect 195978 34368 195980 34377
rect 196032 34368 196034 34377
rect 195978 34303 196034 34312
rect 196084 33969 196112 34410
rect 196070 33960 196126 33969
rect 196070 33895 196126 33904
rect 102322 33552 102378 33561
rect 102322 33487 102378 33496
rect 102140 33108 102192 33114
rect 102140 33050 102192 33056
rect 102138 32464 102194 32473
rect 102138 32399 102194 32408
rect 102152 31754 102180 32399
rect 102230 31784 102286 31793
rect 102140 31748 102192 31754
rect 102230 31719 102286 31728
rect 102140 31690 102192 31696
rect 102138 30560 102194 30569
rect 102138 30495 102194 30504
rect 102152 30326 102180 30495
rect 102140 30320 102192 30326
rect 102140 30262 102192 30268
rect 102244 30258 102272 31719
rect 102336 31686 102364 33487
rect 195980 33108 196032 33114
rect 195980 33050 196032 33056
rect 195992 33017 196020 33050
rect 195978 33008 196034 33017
rect 195978 32943 196034 32952
rect 196072 31748 196124 31754
rect 196072 31690 196124 31696
rect 102324 31680 102376 31686
rect 195980 31680 196032 31686
rect 102324 31622 102376 31628
rect 195978 31648 195980 31657
rect 196032 31648 196034 31657
rect 195978 31583 196034 31592
rect 196084 31521 196112 31690
rect 196070 31512 196126 31521
rect 196070 31447 196126 31456
rect 196072 30320 196124 30326
rect 196072 30262 196124 30268
rect 102232 30252 102284 30258
rect 102232 30194 102284 30200
rect 195980 30252 196032 30258
rect 195980 30194 196032 30200
rect 195992 30161 196020 30194
rect 195978 30152 196034 30161
rect 195978 30087 196034 30096
rect 196084 29753 196112 30262
rect 196070 29744 196126 29753
rect 196070 29679 196126 29688
rect 102138 29336 102194 29345
rect 102138 29271 102194 29280
rect 102152 28966 102180 29271
rect 102140 28960 102192 28966
rect 195980 28960 196032 28966
rect 102140 28902 102192 28908
rect 195978 28928 195980 28937
rect 196032 28928 196034 28937
rect 195978 28863 196034 28872
rect 102138 28520 102194 28529
rect 102138 28455 102194 28464
rect 102152 28286 102180 28455
rect 102140 28280 102192 28286
rect 102140 28222 102192 28228
rect 195980 28280 196032 28286
rect 195980 28222 196032 28228
rect 195992 28121 196020 28222
rect 195978 28112 196034 28121
rect 195978 28047 196034 28056
rect 102138 27704 102194 27713
rect 102138 27639 102194 27648
rect 102152 27606 102180 27639
rect 102140 27600 102192 27606
rect 102140 27542 102192 27548
rect 195980 27600 196032 27606
rect 195980 27542 196032 27548
rect 195992 27305 196020 27542
rect 195978 27296 196034 27305
rect 195978 27231 196034 27240
rect 102782 26344 102838 26353
rect 102782 26279 102838 26288
rect 102796 26246 102824 26279
rect 102784 26240 102836 26246
rect 195980 26240 196032 26246
rect 102784 26182 102836 26188
rect 195978 26208 195980 26217
rect 196032 26208 196034 26217
rect 195978 26143 196034 26152
rect 60004 22296 60056 22302
rect 60004 22238 60056 22244
rect 62316 22098 62344 24140
rect 66272 24126 66746 24154
rect 62304 22092 62356 22098
rect 62304 22034 62356 22040
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3424 10328 3476 10334
rect 3424 10270 3476 10276
rect 3436 6497 3464 10270
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 66272 3466 66300 24126
rect 71148 17270 71176 24140
rect 74552 24126 75578 24154
rect 78692 24126 79994 24154
rect 84212 24126 84410 24154
rect 88352 24126 88826 24154
rect 92492 24126 93242 24154
rect 96632 24126 97658 24154
rect 71136 17264 71188 17270
rect 71136 17206 71188 17212
rect 74552 15910 74580 24126
rect 74540 15904 74592 15910
rect 74540 15846 74592 15852
rect 78692 6186 78720 24126
rect 84212 8974 84240 24126
rect 85488 23520 85540 23526
rect 85488 23462 85540 23468
rect 85500 22098 85528 23462
rect 85488 22092 85540 22098
rect 85488 22034 85540 22040
rect 84200 8968 84252 8974
rect 84200 8910 84252 8916
rect 88352 7614 88380 24126
rect 88340 7608 88392 7614
rect 88340 7550 88392 7556
rect 92492 6254 92520 24126
rect 92480 6248 92532 6254
rect 92480 6190 92532 6196
rect 78680 6180 78732 6186
rect 78680 6122 78732 6128
rect 96632 4826 96660 24126
rect 199396 21894 199424 700266
rect 202800 699854 202828 703520
rect 200028 699848 200080 699854
rect 200028 699790 200080 699796
rect 202788 699848 202840 699854
rect 202788 699790 202840 699796
rect 199476 70440 199528 70446
rect 199476 70382 199528 70388
rect 199384 21888 199436 21894
rect 199384 21830 199436 21836
rect 199488 21826 199516 70382
rect 200040 22098 200068 699790
rect 218072 586401 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 412652 667214 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 462332 701010 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 418160 701004 418212 701010
rect 418160 700946 418212 700952
rect 462320 701004 462372 701010
rect 462320 700946 462372 700952
rect 418172 699825 418200 700946
rect 418158 699816 418214 699825
rect 418158 699751 418214 699760
rect 300860 667208 300912 667214
rect 300860 667150 300912 667156
rect 412640 667208 412692 667214
rect 412640 667150 412692 667156
rect 300872 596174 300900 667150
rect 300872 596146 301452 596174
rect 301424 588690 301452 596146
rect 301424 588662 301990 588690
rect 304552 586566 304580 587316
rect 304540 586560 304592 586566
rect 304540 586502 304592 586508
rect 218058 586392 218114 586401
rect 218058 586327 218114 586336
rect 300768 586152 300820 586158
rect 300768 586094 300820 586100
rect 300584 586084 300636 586090
rect 300584 586026 300636 586032
rect 299388 585948 299440 585954
rect 299388 585890 299440 585896
rect 299112 585880 299164 585886
rect 298006 585848 298062 585857
rect 299112 585822 299164 585828
rect 298006 585783 298062 585792
rect 297916 583228 297968 583234
rect 297916 583170 297968 583176
rect 296628 583160 296680 583166
rect 296628 583102 296680 583108
rect 296536 583092 296588 583098
rect 296536 583034 296588 583040
rect 247040 544400 247092 544406
rect 247040 544342 247092 544348
rect 245660 541680 245712 541686
rect 245660 541622 245712 541628
rect 244280 458856 244332 458862
rect 244280 458798 244332 458804
rect 229742 331936 229798 331945
rect 229742 331871 229798 331880
rect 210424 75404 210476 75410
rect 210424 75346 210476 75352
rect 207664 65680 207716 65686
rect 207664 65622 207716 65628
rect 206008 60172 206060 60178
rect 206008 60114 206060 60120
rect 204352 58880 204404 58886
rect 204352 58822 204404 58828
rect 202880 58744 202932 58750
rect 202880 58686 202932 58692
rect 202892 54754 202920 58686
rect 204364 54754 204392 58822
rect 206020 54754 206048 60114
rect 207676 54754 207704 65622
rect 209320 59424 209372 59430
rect 209320 59366 209372 59372
rect 209332 54754 209360 59366
rect 210436 58886 210464 75346
rect 224224 72684 224276 72690
rect 224224 72626 224276 72632
rect 212632 72616 212684 72622
rect 212632 72558 212684 72564
rect 211160 63028 211212 63034
rect 211160 62970 211212 62976
rect 210424 58880 210476 58886
rect 210424 58822 210476 58828
rect 211172 54754 211200 62970
rect 212644 54754 212672 72558
rect 222568 69896 222620 69902
rect 222568 69838 222620 69844
rect 215944 69828 215996 69834
rect 215944 69770 215996 69776
rect 214288 64388 214340 64394
rect 214288 64330 214340 64336
rect 214300 54754 214328 64330
rect 215956 54754 215984 69770
rect 217600 61600 217652 61606
rect 217600 61542 217652 61548
rect 217612 54754 217640 61542
rect 220912 61396 220964 61402
rect 220912 61338 220964 61344
rect 219440 60036 219492 60042
rect 219440 59978 219492 59984
rect 219452 54754 219480 59978
rect 220924 54754 220952 61338
rect 222580 54754 222608 69838
rect 224236 54754 224264 72626
rect 227720 69964 227772 69970
rect 227720 69906 227772 69912
rect 226246 57352 226302 57361
rect 226246 57287 226302 57296
rect 202892 54726 203090 54754
rect 204364 54726 204746 54754
rect 206020 54726 206402 54754
rect 207676 54726 208058 54754
rect 209332 54726 209714 54754
rect 211172 54726 211370 54754
rect 212644 54726 213026 54754
rect 214300 54726 214682 54754
rect 215956 54726 216338 54754
rect 217612 54726 217994 54754
rect 219452 54726 219650 54754
rect 220924 54726 221306 54754
rect 222580 54726 222962 54754
rect 224236 54726 224618 54754
rect 226260 54740 226288 57287
rect 227732 54754 227760 69906
rect 229756 68542 229784 331871
rect 241518 331800 241574 331809
rect 241518 331735 241574 331744
rect 240140 203652 240192 203658
rect 240140 203594 240192 203600
rect 231124 75336 231176 75342
rect 231124 75278 231176 75284
rect 229192 68536 229244 68542
rect 229192 68478 229244 68484
rect 229744 68536 229796 68542
rect 229744 68478 229796 68484
rect 229204 54754 229232 68478
rect 231136 60110 231164 75278
rect 240152 74534 240180 203594
rect 241532 74534 241560 331735
rect 240152 74506 240824 74534
rect 241532 74506 242480 74534
rect 232504 65748 232556 65754
rect 232504 65690 232556 65696
rect 231124 60104 231176 60110
rect 231124 60046 231176 60052
rect 230846 59936 230902 59945
rect 230846 59871 230902 59880
rect 230860 54754 230888 59871
rect 232516 54754 232544 65690
rect 236000 65612 236052 65618
rect 236000 65554 236052 65560
rect 234160 58880 234212 58886
rect 234160 58822 234212 58828
rect 234172 54754 234200 58822
rect 236012 54754 236040 65554
rect 237472 65544 237524 65550
rect 237472 65486 237524 65492
rect 237484 54754 237512 65486
rect 239128 61736 239180 61742
rect 239128 61678 239180 61684
rect 239140 54754 239168 61678
rect 240796 54754 240824 74506
rect 242452 54754 242480 74506
rect 244292 54754 244320 458798
rect 245672 74534 245700 541622
rect 247052 74534 247080 544342
rect 262220 543040 262272 543046
rect 262220 542982 262272 542988
rect 248420 416084 248472 416090
rect 248420 416026 248472 416032
rect 248432 74534 248460 416026
rect 260840 413296 260892 413302
rect 260840 413238 260892 413244
rect 249800 287700 249852 287706
rect 249800 287642 249852 287648
rect 249812 74534 249840 287642
rect 258080 284980 258132 284986
rect 258080 284922 258132 284928
rect 252560 164892 252612 164898
rect 252560 164834 252612 164840
rect 245672 74506 245792 74534
rect 247052 74506 247448 74534
rect 248432 74506 249104 74534
rect 249812 74506 250760 74534
rect 245764 54754 245792 74506
rect 247420 54754 247448 74506
rect 249076 54754 249104 74506
rect 250732 54754 250760 74506
rect 252572 54754 252600 164834
rect 256700 158024 256752 158030
rect 256700 157966 256752 157972
rect 254584 75268 254636 75274
rect 254584 75210 254636 75216
rect 254032 65612 254084 65618
rect 254032 65554 254084 65560
rect 254044 54754 254072 65554
rect 254596 58886 254624 75210
rect 256712 74534 256740 157966
rect 258092 74534 258120 284922
rect 256712 74506 257384 74534
rect 258092 74506 259040 74534
rect 255688 67040 255740 67046
rect 255688 66982 255740 66988
rect 254584 58880 254636 58886
rect 254584 58822 254636 58828
rect 255700 54754 255728 66982
rect 257356 54754 257384 74506
rect 259012 54754 259040 74506
rect 260852 54754 260880 413238
rect 262232 74534 262260 542982
rect 263600 541680 263652 541686
rect 263600 541622 263652 541628
rect 295982 541648 296038 541657
rect 263612 74534 263640 541622
rect 295982 541583 296038 541592
rect 264980 458856 265032 458862
rect 264980 458798 265032 458804
rect 269762 458824 269818 458833
rect 264992 74534 265020 458798
rect 269762 458759 269818 458768
rect 266360 331900 266412 331906
rect 266360 331842 266412 331848
rect 266372 74534 266400 331842
rect 269120 158024 269172 158030
rect 269120 157966 269172 157972
rect 262232 74506 262352 74534
rect 263612 74506 264008 74534
rect 264992 74506 265664 74534
rect 266372 74506 267320 74534
rect 262324 54754 262352 74506
rect 263980 54754 264008 74506
rect 265636 54754 265664 74506
rect 267292 54754 267320 74506
rect 269132 54754 269160 157966
rect 269776 77994 269804 458759
rect 295248 204332 295300 204338
rect 295248 204274 295300 204280
rect 282184 203584 282236 203590
rect 282184 203526 282236 203532
rect 269764 77988 269816 77994
rect 269764 77930 269816 77936
rect 280804 75404 280856 75410
rect 280804 75346 280856 75352
rect 273260 75336 273312 75342
rect 273260 75278 273312 75284
rect 273272 74534 273300 75278
rect 277400 75268 277452 75274
rect 277400 75210 277452 75216
rect 273272 74506 273944 74534
rect 270592 71256 270644 71262
rect 270592 71198 270644 71204
rect 270604 54754 270632 71198
rect 272248 65544 272300 65550
rect 272248 65486 272300 65492
rect 272260 54754 272288 65486
rect 273916 54754 273944 74506
rect 275928 57452 275980 57458
rect 275928 57394 275980 57400
rect 227732 54726 227930 54754
rect 229204 54726 229586 54754
rect 230860 54726 231242 54754
rect 232516 54726 232898 54754
rect 234172 54726 234554 54754
rect 236012 54726 236210 54754
rect 237484 54726 237866 54754
rect 239140 54726 239522 54754
rect 240796 54726 241178 54754
rect 242452 54726 242834 54754
rect 244292 54726 244490 54754
rect 245764 54726 246146 54754
rect 247420 54726 247802 54754
rect 249076 54726 249458 54754
rect 250732 54726 251114 54754
rect 252572 54726 252770 54754
rect 254044 54726 254426 54754
rect 255700 54726 256082 54754
rect 257356 54726 257738 54754
rect 259012 54726 259394 54754
rect 260852 54726 261050 54754
rect 262324 54726 262706 54754
rect 263980 54726 264362 54754
rect 265636 54726 266018 54754
rect 267292 54726 267674 54754
rect 269132 54726 269330 54754
rect 270604 54726 270986 54754
rect 272260 54726 272642 54754
rect 273916 54726 274298 54754
rect 275940 54740 275968 57394
rect 277412 54754 277440 75210
rect 280816 65618 280844 75346
rect 280804 65612 280856 65618
rect 280804 65554 280856 65560
rect 280528 61532 280580 61538
rect 280528 61474 280580 61480
rect 279240 57520 279292 57526
rect 279240 57462 279292 57468
rect 277412 54726 277610 54754
rect 279252 54740 279280 57462
rect 280540 54754 280568 61474
rect 282196 61470 282224 203526
rect 285680 75200 285732 75206
rect 285680 75142 285732 75148
rect 283840 72752 283892 72758
rect 283840 72694 283892 72700
rect 282092 61464 282144 61470
rect 282092 61406 282144 61412
rect 282184 61464 282236 61470
rect 282184 61406 282236 61412
rect 282104 55214 282132 61406
rect 282104 55186 282224 55214
rect 282196 54754 282224 55186
rect 283852 54754 283880 72694
rect 285692 54754 285720 75142
rect 290464 68468 290516 68474
rect 290464 68410 290516 68416
rect 288808 58880 288860 58886
rect 288808 58822 288860 58828
rect 287520 57316 287572 57322
rect 287520 57258 287572 57264
rect 280540 54726 280922 54754
rect 282196 54726 282578 54754
rect 283852 54726 284234 54754
rect 285692 54726 285890 54754
rect 287532 54740 287560 57258
rect 288820 54754 288848 58822
rect 290476 57594 290504 68410
rect 292120 67040 292172 67046
rect 292120 66982 292172 66988
rect 290464 57588 290516 57594
rect 290464 57530 290516 57536
rect 290832 57248 290884 57254
rect 290832 57190 290884 57196
rect 288820 54726 289202 54754
rect 290844 54740 290872 57190
rect 292132 54754 292160 66982
rect 293960 65612 294012 65618
rect 293960 65554 294012 65560
rect 293972 54754 294000 65554
rect 295260 60722 295288 204274
rect 295340 66224 295392 66230
rect 295340 66166 295392 66172
rect 295352 65686 295380 66166
rect 295340 65680 295392 65686
rect 295340 65622 295392 65628
rect 294052 60716 294104 60722
rect 294052 60658 294104 60664
rect 295248 60716 295300 60722
rect 295248 60658 295300 60664
rect 294064 60178 294092 60658
rect 294052 60172 294104 60178
rect 294052 60114 294104 60120
rect 295432 58880 295484 58886
rect 295432 58822 295484 58828
rect 295444 54754 295472 58822
rect 295996 57254 296024 541583
rect 296548 458930 296576 583034
rect 296640 458998 296668 583102
rect 297732 583024 297784 583030
rect 297732 582966 297784 582972
rect 296628 458992 296680 458998
rect 296628 458934 296680 458940
rect 296536 458924 296588 458930
rect 296536 458866 296588 458872
rect 297548 458924 297600 458930
rect 297548 458866 297600 458872
rect 297560 306374 297588 458866
rect 297640 458244 297692 458250
rect 297640 458186 297692 458192
rect 297652 332654 297680 458186
rect 297744 456686 297772 582966
rect 297824 541748 297876 541754
rect 297824 541690 297876 541696
rect 297836 459950 297864 541690
rect 297824 459944 297876 459950
rect 297824 459886 297876 459892
rect 297928 459542 297956 583170
rect 298020 460902 298048 585783
rect 298928 462664 298980 462670
rect 298928 462606 298980 462612
rect 298008 460896 298060 460902
rect 298008 460838 298060 460844
rect 298836 460216 298888 460222
rect 298836 460158 298888 460164
rect 298848 459950 298876 460158
rect 298836 459944 298888 459950
rect 298836 459886 298888 459892
rect 297916 459536 297968 459542
rect 297916 459478 297968 459484
rect 297928 459082 297956 459478
rect 297928 459054 298048 459082
rect 297916 458992 297968 458998
rect 297916 458934 297968 458940
rect 297732 456680 297784 456686
rect 297732 456622 297784 456628
rect 297640 332648 297692 332654
rect 297640 332590 297692 332596
rect 297560 306346 297680 306374
rect 296628 287088 296680 287094
rect 296628 287030 296680 287036
rect 296076 285048 296128 285054
rect 296076 284990 296128 284996
rect 296088 57322 296116 284990
rect 296640 201414 296668 287030
rect 297652 285569 297680 306346
rect 297744 288318 297772 456622
rect 297732 288312 297784 288318
rect 297732 288254 297784 288260
rect 297744 287094 297772 288254
rect 297732 287088 297784 287094
rect 297928 287054 297956 458934
rect 297732 287030 297784 287036
rect 297836 287026 297956 287054
rect 297836 285666 297864 287026
rect 297824 285660 297876 285666
rect 297824 285602 297876 285608
rect 297638 285560 297694 285569
rect 297638 285495 297694 285504
rect 297548 204876 297600 204882
rect 297548 204818 297600 204824
rect 296628 201408 296680 201414
rect 296628 201350 296680 201356
rect 296640 66230 296668 201350
rect 297364 158092 297416 158098
rect 297364 158034 297416 158040
rect 297088 68468 297140 68474
rect 297088 68410 297140 68416
rect 296628 66224 296680 66230
rect 296628 66166 296680 66172
rect 296076 57316 296128 57322
rect 296076 57258 296128 57264
rect 295984 57248 296036 57254
rect 295984 57190 296036 57196
rect 297100 54754 297128 68410
rect 297376 57390 297404 158034
rect 297560 78130 297588 204818
rect 297652 204338 297680 285495
rect 297732 284368 297784 284374
rect 297732 284310 297784 284316
rect 297640 204332 297692 204338
rect 297640 204274 297692 204280
rect 297744 158574 297772 284310
rect 297836 158642 297864 285602
rect 298020 285598 298048 459054
rect 298848 330546 298876 459886
rect 298940 331809 298968 462606
rect 299124 462330 299152 585822
rect 299296 583432 299348 583438
rect 299296 583374 299348 583380
rect 299204 583364 299256 583370
rect 299204 583306 299256 583312
rect 299112 462324 299164 462330
rect 299112 462266 299164 462272
rect 299216 460934 299244 583306
rect 299124 460906 299244 460934
rect 299124 459406 299152 460906
rect 299112 459400 299164 459406
rect 299112 459342 299164 459348
rect 299020 456816 299072 456822
rect 299020 456758 299072 456764
rect 299032 332858 299060 456758
rect 299020 332852 299072 332858
rect 299020 332794 299072 332800
rect 299124 332790 299152 459342
rect 299308 458182 299336 583374
rect 299296 458176 299348 458182
rect 299296 458118 299348 458124
rect 299308 456822 299336 458118
rect 299400 458114 299428 585890
rect 300400 585200 300452 585206
rect 300400 585142 300452 585148
rect 300412 470594 300440 585142
rect 300492 583296 300544 583302
rect 300492 583238 300544 583244
rect 300320 470566 300440 470594
rect 300320 459241 300348 470566
rect 300400 462324 300452 462330
rect 300400 462266 300452 462272
rect 300412 461038 300440 462266
rect 300400 461032 300452 461038
rect 300400 460974 300452 460980
rect 300306 459232 300362 459241
rect 300412 459202 300440 460974
rect 300504 459474 300532 583238
rect 300492 459468 300544 459474
rect 300492 459410 300544 459416
rect 300306 459167 300362 459176
rect 300400 459196 300452 459202
rect 299388 458108 299440 458114
rect 299388 458050 299440 458056
rect 299296 456816 299348 456822
rect 299296 456758 299348 456764
rect 299400 451274 299428 458050
rect 299216 451246 299428 451274
rect 299216 345014 299244 451246
rect 299216 344986 299336 345014
rect 299112 332784 299164 332790
rect 299112 332726 299164 332732
rect 298926 331800 298982 331809
rect 298926 331735 298982 331744
rect 298940 331265 298968 331735
rect 298926 331256 298982 331265
rect 298926 331191 298982 331200
rect 299308 331158 299336 344986
rect 300320 332586 300348 459167
rect 300400 459138 300452 459144
rect 300400 459060 300452 459066
rect 300400 459002 300452 459008
rect 300412 458289 300440 459002
rect 300398 458280 300454 458289
rect 300504 458250 300532 459410
rect 300398 458215 300454 458224
rect 300492 458244 300544 458250
rect 300412 332722 300440 458215
rect 300492 458186 300544 458192
rect 300596 457706 300624 586026
rect 300676 459196 300728 459202
rect 300676 459138 300728 459144
rect 300584 457700 300636 457706
rect 300584 457642 300636 457648
rect 300490 456920 300546 456929
rect 300490 456855 300546 456864
rect 300504 345014 300532 456855
rect 300504 344986 300624 345014
rect 300400 332716 300452 332722
rect 300400 332658 300452 332664
rect 300308 332580 300360 332586
rect 300308 332522 300360 332528
rect 300216 331288 300268 331294
rect 299386 331256 299442 331265
rect 300216 331230 300268 331236
rect 299386 331191 299442 331200
rect 299296 331152 299348 331158
rect 299296 331094 299348 331100
rect 298836 330540 298888 330546
rect 298836 330482 298888 330488
rect 298008 285592 298060 285598
rect 298008 285534 298060 285540
rect 297916 285116 297968 285122
rect 297916 285058 297968 285064
rect 297928 204814 297956 285058
rect 298020 284374 298048 285534
rect 299204 285184 299256 285190
rect 299204 285126 299256 285132
rect 299020 285048 299072 285054
rect 299020 284990 299072 284996
rect 298008 284368 298060 284374
rect 298008 284310 298060 284316
rect 298928 204944 298980 204950
rect 298928 204886 298980 204892
rect 297916 204808 297968 204814
rect 297916 204750 297968 204756
rect 298008 204740 298060 204746
rect 298008 204682 298060 204688
rect 297824 158636 297876 158642
rect 297824 158578 297876 158584
rect 297732 158568 297784 158574
rect 297732 158510 297784 158516
rect 297548 78124 297600 78130
rect 297548 78066 297600 78072
rect 297744 75478 297772 158510
rect 297732 75472 297784 75478
rect 297732 75414 297784 75420
rect 297836 75206 297864 158578
rect 298020 75546 298048 204682
rect 298008 75540 298060 75546
rect 298008 75482 298060 75488
rect 297824 75200 297876 75206
rect 297824 75142 297876 75148
rect 298940 74458 298968 204886
rect 299032 204882 299060 284990
rect 299112 284980 299164 284986
rect 299112 284922 299164 284928
rect 299020 204876 299072 204882
rect 299020 204818 299072 204824
rect 299032 204474 299060 204818
rect 299124 204746 299152 284922
rect 299112 204740 299164 204746
rect 299112 204682 299164 204688
rect 299020 204468 299072 204474
rect 299020 204410 299072 204416
rect 299124 204406 299152 204682
rect 299112 204400 299164 204406
rect 299112 204342 299164 204348
rect 299112 204196 299164 204202
rect 299112 204138 299164 204144
rect 299124 203862 299152 204138
rect 299112 203856 299164 203862
rect 299112 203798 299164 203804
rect 299020 200660 299072 200666
rect 299020 200602 299072 200608
rect 299032 76566 299060 200602
rect 299020 76560 299072 76566
rect 299020 76502 299072 76508
rect 298928 74452 298980 74458
rect 298928 74394 298980 74400
rect 299124 74322 299152 203798
rect 299216 203561 299244 285126
rect 299308 204066 299336 331094
rect 299400 204202 299428 331191
rect 300228 325694 300256 331230
rect 300320 330834 300348 332522
rect 300596 332178 300624 344986
rect 300688 332926 300716 459138
rect 300780 458153 300808 586094
rect 301228 586016 301280 586022
rect 301228 585958 301280 585964
rect 301240 462670 301268 585958
rect 301412 585812 301464 585818
rect 301412 585754 301464 585760
rect 301318 585712 301374 585721
rect 301318 585647 301374 585656
rect 301228 462664 301280 462670
rect 301228 462606 301280 462612
rect 301332 461009 301360 585647
rect 301318 461000 301374 461009
rect 301424 460970 301452 585754
rect 307128 585206 307156 587316
rect 309704 586158 309732 587316
rect 309692 586152 309744 586158
rect 309692 586094 309744 586100
rect 312280 586090 312308 587316
rect 312268 586084 312320 586090
rect 312268 586026 312320 586032
rect 314856 586022 314884 587316
rect 314844 586016 314896 586022
rect 314844 585958 314896 585964
rect 317432 585954 317460 587316
rect 317420 585948 317472 585954
rect 317420 585890 317472 585896
rect 320008 585886 320036 587316
rect 319996 585880 320048 585886
rect 319996 585822 320048 585828
rect 307116 585200 307168 585206
rect 307116 585142 307168 585148
rect 322584 583438 322612 587316
rect 322572 583432 322624 583438
rect 322572 583374 322624 583380
rect 325160 583370 325188 587316
rect 325148 583364 325200 583370
rect 325148 583306 325200 583312
rect 327736 583001 327764 587316
rect 330312 583302 330340 587316
rect 332888 585818 332916 587316
rect 332876 585812 332928 585818
rect 332876 585754 332928 585760
rect 335464 585721 335492 587316
rect 338040 585993 338068 587316
rect 338026 585984 338082 585993
rect 338026 585919 338082 585928
rect 335450 585712 335506 585721
rect 335450 585647 335506 585656
rect 330300 583296 330352 583302
rect 330300 583238 330352 583244
rect 340616 583234 340644 587316
rect 340604 583228 340656 583234
rect 340604 583170 340656 583176
rect 343192 583166 343220 587316
rect 345032 587302 345782 587330
rect 348358 587302 348464 587330
rect 343180 583160 343232 583166
rect 343180 583102 343232 583108
rect 327722 582992 327778 583001
rect 327722 582927 327778 582936
rect 345032 541754 345060 587302
rect 348436 586498 348464 587302
rect 350920 586498 350948 587316
rect 348424 586492 348476 586498
rect 348424 586434 348476 586440
rect 350908 586492 350960 586498
rect 350908 586434 350960 586440
rect 345020 541748 345072 541754
rect 345020 541690 345072 541696
rect 348436 541686 348464 586434
rect 353496 583098 353524 587316
rect 353484 583092 353536 583098
rect 353484 583034 353536 583040
rect 356072 583030 356100 587316
rect 358648 585857 358676 587316
rect 358634 585848 358690 585857
rect 358634 585783 358690 585792
rect 356060 583024 356112 583030
rect 356060 582966 356112 582972
rect 361224 580281 361252 587316
rect 363800 583030 363828 587316
rect 366376 583098 366404 587316
rect 368952 583166 368980 587316
rect 371252 587302 371542 587330
rect 374012 587302 374118 587330
rect 375392 587302 376694 587330
rect 378152 587302 379270 587330
rect 380912 587302 381846 587330
rect 368940 583160 368992 583166
rect 368940 583102 368992 583108
rect 366364 583092 366416 583098
rect 366364 583034 366416 583040
rect 363788 583024 363840 583030
rect 363788 582966 363840 582972
rect 361210 580272 361266 580281
rect 361210 580207 361266 580216
rect 371252 541686 371280 587302
rect 374012 541754 374040 587302
rect 375392 541822 375420 587302
rect 378152 544406 378180 587302
rect 378140 544400 378192 544406
rect 378140 544342 378192 544348
rect 380912 541890 380940 587302
rect 384408 585721 384436 587316
rect 384394 585712 384450 585721
rect 384394 585647 384450 585656
rect 386984 583234 387012 587316
rect 389560 583302 389588 587316
rect 392136 583370 392164 587316
rect 394712 583438 394740 587316
rect 397288 585818 397316 587316
rect 399864 585886 399892 587316
rect 402440 585954 402468 587316
rect 405016 586022 405044 587316
rect 407592 586090 407620 587316
rect 410168 586158 410196 587316
rect 410156 586152 410208 586158
rect 410156 586094 410208 586100
rect 407580 586084 407632 586090
rect 407580 586026 407632 586032
rect 405004 586016 405056 586022
rect 405004 585958 405056 585964
rect 402428 585948 402480 585954
rect 402428 585890 402480 585896
rect 399852 585880 399904 585886
rect 412744 585857 412772 587316
rect 415320 586022 415348 587316
rect 415308 586016 415360 586022
rect 415308 585958 415360 585964
rect 415124 585948 415176 585954
rect 415124 585890 415176 585896
rect 399852 585822 399904 585828
rect 412730 585848 412786 585857
rect 397276 585812 397328 585818
rect 412730 585783 412786 585792
rect 397276 585754 397328 585760
rect 415136 585750 415164 585890
rect 415124 585744 415176 585750
rect 415124 585686 415176 585692
rect 417896 585177 417924 587316
rect 477512 586566 477540 702406
rect 527192 697610 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 697604 527232 697610
rect 527180 697546 527232 697552
rect 527824 697604 527876 697610
rect 527824 697546 527876 697552
rect 477500 586560 477552 586566
rect 477500 586502 477552 586508
rect 418804 586152 418856 586158
rect 418804 586094 418856 586100
rect 418436 585948 418488 585954
rect 418436 585890 418488 585896
rect 418344 585880 418396 585886
rect 418344 585822 418396 585828
rect 418250 585712 418306 585721
rect 418250 585647 418306 585656
rect 417882 585168 417938 585177
rect 417882 585103 417938 585112
rect 394700 583432 394752 583438
rect 394700 583374 394752 583380
rect 392124 583364 392176 583370
rect 392124 583306 392176 583312
rect 389548 583296 389600 583302
rect 389548 583238 389600 583244
rect 386972 583228 387024 583234
rect 386972 583170 387024 583176
rect 380900 541884 380952 541890
rect 380900 541826 380952 541832
rect 375380 541816 375432 541822
rect 375380 541758 375432 541764
rect 374000 541748 374052 541754
rect 374000 541690 374052 541696
rect 348424 541680 348476 541686
rect 348424 541622 348476 541628
rect 371240 541680 371292 541686
rect 371240 541622 371292 541628
rect 314660 462664 314712 462670
rect 382096 462664 382148 462670
rect 314712 462612 314870 462618
rect 314660 462606 314870 462612
rect 314672 462590 314870 462606
rect 381846 462612 382096 462618
rect 381846 462606 382148 462612
rect 385500 462664 385552 462670
rect 385500 462606 385552 462612
rect 381846 462590 382136 462606
rect 348608 461304 348660 461310
rect 348358 461252 348608 461258
rect 348358 461246 348660 461252
rect 350540 461304 350592 461310
rect 350592 461252 350934 461258
rect 350540 461246 350934 461252
rect 348358 461244 348648 461246
rect 301318 460935 301374 460944
rect 301412 460964 301464 460970
rect 300766 458144 300822 458153
rect 300766 458079 300822 458088
rect 300780 456929 300808 458079
rect 301228 457700 301280 457706
rect 301228 457642 301280 457648
rect 301240 457502 301268 457642
rect 301228 457496 301280 457502
rect 301228 457438 301280 457444
rect 300766 456920 300822 456929
rect 300766 456855 300822 456864
rect 300860 456748 300912 456754
rect 300860 456690 300912 456696
rect 300872 456634 300900 456690
rect 300780 456606 300900 456634
rect 300676 332920 300728 332926
rect 300676 332862 300728 332868
rect 300584 332172 300636 332178
rect 300584 332114 300636 332120
rect 300596 331106 300624 332114
rect 300596 331078 300716 331106
rect 300320 330806 300624 330834
rect 300228 325666 300532 325694
rect 300400 285252 300452 285258
rect 300400 285194 300452 285200
rect 300412 204950 300440 285194
rect 300400 204944 300452 204950
rect 300400 204886 300452 204892
rect 300308 204808 300360 204814
rect 300308 204750 300360 204756
rect 300320 204542 300348 204750
rect 300308 204536 300360 204542
rect 300308 204478 300360 204484
rect 299388 204196 299440 204202
rect 299388 204138 299440 204144
rect 299296 204060 299348 204066
rect 299296 204002 299348 204008
rect 299202 203552 299258 203561
rect 299202 203487 299258 203496
rect 299112 74316 299164 74322
rect 299112 74258 299164 74264
rect 299216 74186 299244 203487
rect 299308 74390 299336 204002
rect 300320 75614 300348 204478
rect 300504 204134 300532 325666
rect 300596 204202 300624 330806
rect 300584 204196 300636 204202
rect 300584 204138 300636 204144
rect 300492 204128 300544 204134
rect 300492 204070 300544 204076
rect 300504 200114 300532 204070
rect 300412 200086 300532 200114
rect 300412 78062 300440 200086
rect 300596 78674 300624 204138
rect 300688 203930 300716 331078
rect 300780 288386 300808 456606
rect 301240 335354 301268 457438
rect 301056 335326 301268 335354
rect 301056 332382 301084 335326
rect 301332 332450 301360 460935
rect 301412 460906 301464 460912
rect 301320 332444 301372 332450
rect 301320 332386 301372 332392
rect 301044 332376 301096 332382
rect 301044 332318 301096 332324
rect 300768 288380 300820 288386
rect 300768 288322 300820 288328
rect 300676 203924 300728 203930
rect 300676 203866 300728 203872
rect 300584 78668 300636 78674
rect 300584 78610 300636 78616
rect 300400 78056 300452 78062
rect 300400 77998 300452 78004
rect 300308 75608 300360 75614
rect 300308 75550 300360 75556
rect 300688 74526 300716 203866
rect 300780 201482 300808 288322
rect 300952 206644 301004 206650
rect 300952 206586 301004 206592
rect 300768 201476 300820 201482
rect 300768 201418 300820 201424
rect 300676 74520 300728 74526
rect 300676 74462 300728 74468
rect 299296 74384 299348 74390
rect 299296 74326 299348 74332
rect 299204 74180 299256 74186
rect 299204 74122 299256 74128
rect 300400 72684 300452 72690
rect 300400 72626 300452 72632
rect 298744 69896 298796 69902
rect 298744 69838 298796 69844
rect 297364 57384 297416 57390
rect 297364 57326 297416 57332
rect 298756 54754 298784 69838
rect 300412 54754 300440 72626
rect 300780 63510 300808 201418
rect 300964 201346 300992 206586
rect 301056 206514 301084 332318
rect 301228 330540 301280 330546
rect 301228 330482 301280 330488
rect 301240 215294 301268 330482
rect 301148 215266 301268 215294
rect 301148 206650 301176 215266
rect 301136 206644 301188 206650
rect 301136 206586 301188 206592
rect 301044 206508 301096 206514
rect 301044 206450 301096 206456
rect 301332 204898 301360 332386
rect 301424 332314 301452 460906
rect 301976 459377 302004 461244
rect 302700 460896 302752 460902
rect 302700 460838 302752 460844
rect 302712 459649 302740 460838
rect 302698 459640 302754 459649
rect 302698 459575 302754 459584
rect 304552 459513 304580 461244
rect 304538 459504 304594 459513
rect 304538 459439 304594 459448
rect 301962 459368 302018 459377
rect 301962 459303 302018 459312
rect 307128 459241 307156 461244
rect 307114 459232 307170 459241
rect 307114 459167 307170 459176
rect 309704 458153 309732 461244
rect 309690 458144 309746 458153
rect 309690 458079 309746 458088
rect 312280 457502 312308 461244
rect 317432 458114 317460 461244
rect 320008 461038 320036 461244
rect 319996 461032 320048 461038
rect 319996 460974 320048 460980
rect 322584 458182 322612 461244
rect 325160 459406 325188 461244
rect 325148 459400 325200 459406
rect 325148 459342 325200 459348
rect 327736 459066 327764 461244
rect 330312 459474 330340 461244
rect 332888 460970 332916 461244
rect 335464 461009 335492 461244
rect 338040 461145 338068 461244
rect 338026 461136 338082 461145
rect 338026 461071 338082 461080
rect 335450 461000 335506 461009
rect 332876 460964 332928 460970
rect 335450 460935 335506 460944
rect 332876 460906 332928 460912
rect 340616 459542 340644 461244
rect 340604 459536 340656 459542
rect 340604 459478 340656 459484
rect 330300 459468 330352 459474
rect 330300 459410 330352 459416
rect 327724 459060 327776 459066
rect 327724 459002 327776 459008
rect 343192 458998 343220 461244
rect 345768 460222 345796 461244
rect 348344 461230 348648 461244
rect 350552 461230 350934 461246
rect 345756 460216 345808 460222
rect 345756 460158 345808 460164
rect 343180 458992 343232 458998
rect 343180 458934 343232 458940
rect 348344 458862 348372 461230
rect 353496 458930 353524 461244
rect 353484 458924 353536 458930
rect 353484 458866 353536 458872
rect 348332 458856 348384 458862
rect 348332 458798 348384 458804
rect 322572 458176 322624 458182
rect 322572 458118 322624 458124
rect 317420 458108 317472 458114
rect 317420 458050 317472 458056
rect 312268 457496 312320 457502
rect 312268 457438 312320 457444
rect 301502 456784 301558 456793
rect 301502 456719 301504 456728
rect 301556 456719 301558 456728
rect 301504 456690 301556 456696
rect 356072 456686 356100 461244
rect 358648 460902 358676 461244
rect 358636 460896 358688 460902
rect 358636 460838 358688 460844
rect 361224 456754 361252 461244
rect 363800 459338 363828 461244
rect 363788 459332 363840 459338
rect 363788 459274 363840 459280
rect 366376 458930 366404 461244
rect 366364 458924 366416 458930
rect 366364 458866 366416 458872
rect 368952 458862 368980 461244
rect 371528 461038 371556 461244
rect 371516 461032 371568 461038
rect 371516 460974 371568 460980
rect 374104 460970 374132 461244
rect 376680 461106 376708 461244
rect 378152 461230 379270 461258
rect 376668 461100 376720 461106
rect 376668 461042 376720 461048
rect 374092 460964 374144 460970
rect 374092 460906 374144 460912
rect 368940 458856 368992 458862
rect 368940 458798 368992 458804
rect 361212 456748 361264 456754
rect 361212 456690 361264 456696
rect 356060 456680 356112 456686
rect 356060 456622 356112 456628
rect 378152 416090 378180 461230
rect 383568 461100 383620 461106
rect 383568 461042 383620 461048
rect 383580 460834 383608 461042
rect 383568 460828 383620 460834
rect 383568 460770 383620 460776
rect 384408 458182 384436 461244
rect 385512 461038 385540 462606
rect 418160 462256 418212 462262
rect 418160 462198 418212 462204
rect 418068 462188 418120 462194
rect 418068 462130 418120 462136
rect 385500 461032 385552 461038
rect 386984 461009 387012 461244
rect 389560 461145 389588 461244
rect 389546 461136 389602 461145
rect 389546 461071 389602 461080
rect 385500 460974 385552 460980
rect 386970 461000 387026 461009
rect 386970 460935 387026 460944
rect 392136 459474 392164 461244
rect 392124 459468 392176 459474
rect 392124 459410 392176 459416
rect 394712 458998 394740 461244
rect 397288 459542 397316 461244
rect 397276 459536 397328 459542
rect 397276 459478 397328 459484
rect 399864 459066 399892 461244
rect 402440 459542 402468 461244
rect 405016 460970 405044 461244
rect 405004 460964 405056 460970
rect 405004 460906 405056 460912
rect 407026 459640 407082 459649
rect 407026 459575 407082 459584
rect 407040 459542 407068 459575
rect 407592 459542 407620 461244
rect 402428 459536 402480 459542
rect 402428 459478 402480 459484
rect 407028 459536 407080 459542
rect 407028 459478 407080 459484
rect 407580 459536 407632 459542
rect 407580 459478 407632 459484
rect 410168 459406 410196 461244
rect 410156 459400 410208 459406
rect 410156 459342 410208 459348
rect 399852 459060 399904 459066
rect 399852 459002 399904 459008
rect 409880 459060 409932 459066
rect 409880 459002 409932 459008
rect 394700 458992 394752 458998
rect 394700 458934 394752 458940
rect 384396 458176 384448 458182
rect 384396 458118 384448 458124
rect 409892 458114 409920 459002
rect 412744 458289 412772 461244
rect 415216 459672 415268 459678
rect 415216 459614 415268 459620
rect 415228 459542 415256 459614
rect 415320 459542 415348 461244
rect 415216 459536 415268 459542
rect 415216 459478 415268 459484
rect 415308 459536 415360 459542
rect 415308 459478 415360 459484
rect 417896 459270 417924 461244
rect 418080 459542 418108 462130
rect 418172 459649 418200 462198
rect 418158 459640 418214 459649
rect 418158 459575 418214 459584
rect 418068 459536 418120 459542
rect 418068 459478 418120 459484
rect 417884 459264 417936 459270
rect 417884 459206 417936 459212
rect 418160 458924 418212 458930
rect 418160 458866 418212 458872
rect 412730 458280 412786 458289
rect 412730 458215 412786 458224
rect 418172 458182 418200 458866
rect 418068 458176 418120 458182
rect 418068 458118 418120 458124
rect 418160 458176 418212 458182
rect 418160 458118 418212 458124
rect 409880 458108 409932 458114
rect 409880 458050 409932 458056
rect 418080 457994 418108 458118
rect 418264 457994 418292 585647
rect 418356 458114 418384 585822
rect 418448 480254 418476 585890
rect 418448 480226 418568 480254
rect 418436 461780 418488 461786
rect 418436 461722 418488 461728
rect 418448 459610 418476 461722
rect 418540 460970 418568 480226
rect 418816 462330 418844 586094
rect 419540 586084 419592 586090
rect 419540 586026 419592 586032
rect 418804 462324 418856 462330
rect 418804 462266 418856 462272
rect 418528 460964 418580 460970
rect 418528 460906 418580 460912
rect 419552 459678 419580 586026
rect 419632 586016 419684 586022
rect 419632 585958 419684 585964
rect 419644 462466 419672 585958
rect 419816 585812 419868 585818
rect 419816 585754 419868 585760
rect 419724 585744 419776 585750
rect 419724 585686 419776 585692
rect 419632 462460 419684 462466
rect 419632 462402 419684 462408
rect 419632 462324 419684 462330
rect 419632 462266 419684 462272
rect 419644 460934 419672 462266
rect 419736 462262 419764 585686
rect 419724 462256 419776 462262
rect 419724 462198 419776 462204
rect 419828 461786 419856 585754
rect 422298 585168 422354 585177
rect 422298 585103 422354 585112
rect 420920 583432 420972 583438
rect 420920 583374 420972 583380
rect 420828 470620 420880 470626
rect 420828 470562 420880 470568
rect 419816 461780 419868 461786
rect 419816 461722 419868 461728
rect 419644 460906 419764 460934
rect 419540 459672 419592 459678
rect 418710 459640 418766 459649
rect 418436 459604 418488 459610
rect 419540 459614 419592 459620
rect 418710 459575 418766 459584
rect 418436 459546 418488 459552
rect 418344 458108 418396 458114
rect 418344 458050 418396 458056
rect 418080 457966 418292 457994
rect 418264 456822 418292 457966
rect 418252 456816 418304 456822
rect 418252 456758 418304 456764
rect 418356 451274 418384 458050
rect 418448 457314 418476 459546
rect 418448 457286 418660 457314
rect 418528 456816 418580 456822
rect 418528 456758 418580 456764
rect 418356 451246 418476 451274
rect 378140 416084 378192 416090
rect 378140 416026 378192 416032
rect 301976 332489 302004 333268
rect 303528 332512 303580 332518
rect 301962 332480 302018 332489
rect 303528 332454 303580 332460
rect 301962 332415 302018 332424
rect 303540 332353 303568 332454
rect 304552 332353 304580 333268
rect 307128 332586 307156 333268
rect 307116 332580 307168 332586
rect 307116 332522 307168 332528
rect 303526 332344 303582 332353
rect 301412 332308 301464 332314
rect 303526 332279 303582 332288
rect 304538 332344 304594 332353
rect 304538 332279 304594 332288
rect 301412 332250 301464 332256
rect 301424 331294 301452 332250
rect 309704 332178 309732 333268
rect 310980 332512 311032 332518
rect 311032 332460 311204 332466
rect 310980 332454 311204 332460
rect 310992 332450 311204 332454
rect 310992 332444 311216 332450
rect 310992 332438 311164 332444
rect 311164 332386 311216 332392
rect 312280 332382 312308 333268
rect 312268 332376 312320 332382
rect 312268 332318 312320 332324
rect 309692 332172 309744 332178
rect 309692 332114 309744 332120
rect 314856 331974 314884 333268
rect 306748 331968 306800 331974
rect 306748 331910 306800 331916
rect 314844 331968 314896 331974
rect 314844 331910 314896 331916
rect 306760 331809 306788 331910
rect 306746 331800 306802 331809
rect 306746 331735 306802 331744
rect 317432 331294 317460 333268
rect 320008 332926 320036 333268
rect 318800 332920 318852 332926
rect 318800 332862 318852 332868
rect 319996 332920 320048 332926
rect 319996 332862 320048 332868
rect 301412 331288 301464 331294
rect 301412 331230 301464 331236
rect 311900 331288 311952 331294
rect 311900 331230 311952 331236
rect 317420 331288 317472 331294
rect 317420 331230 317472 331236
rect 303528 331220 303580 331226
rect 303528 331162 303580 331168
rect 303540 331129 303568 331162
rect 311912 331158 311940 331230
rect 311900 331152 311952 331158
rect 303526 331120 303582 331129
rect 311900 331094 311952 331100
rect 303526 331055 303582 331064
rect 318812 285258 318840 332862
rect 322584 332858 322612 333268
rect 321560 332852 321612 332858
rect 321560 332794 321612 332800
rect 322572 332852 322624 332858
rect 322572 332794 322624 332800
rect 318800 285252 318852 285258
rect 318800 285194 318852 285200
rect 321572 285190 321600 332794
rect 325160 332790 325188 333268
rect 327276 333254 327750 333282
rect 329852 333254 330326 333282
rect 327276 332858 327304 333254
rect 327264 332852 327316 332858
rect 327264 332794 327316 332800
rect 324320 332784 324372 332790
rect 324320 332726 324372 332732
rect 325148 332784 325200 332790
rect 325148 332726 325200 332732
rect 321560 285184 321612 285190
rect 321560 285126 321612 285132
rect 324332 285122 324360 332726
rect 327276 316034 327304 332794
rect 329852 332654 329880 333254
rect 329840 332648 329892 332654
rect 329840 332590 329892 332596
rect 327092 316006 327304 316034
rect 324320 285116 324372 285122
rect 324320 285058 324372 285064
rect 327092 285054 327120 316006
rect 327080 285048 327132 285054
rect 327080 284990 327132 284996
rect 329852 284986 329880 332590
rect 332888 332450 332916 333268
rect 335464 332586 335492 333268
rect 335452 332580 335504 332586
rect 335452 332522 335504 332528
rect 338040 332518 338068 333268
rect 339512 333254 340630 333282
rect 342272 333254 343206 333282
rect 338028 332512 338080 332518
rect 338028 332454 338080 332460
rect 332876 332444 332928 332450
rect 332876 332386 332928 332392
rect 339512 285598 339540 333254
rect 342272 285666 342300 333254
rect 345768 330546 345796 333268
rect 348344 332586 348372 333268
rect 350920 332586 350948 333268
rect 353312 333254 353510 333282
rect 348332 332580 348384 332586
rect 348332 332522 348384 332528
rect 350908 332580 350960 332586
rect 350908 332522 350960 332528
rect 348344 331906 348372 332522
rect 348332 331900 348384 331906
rect 348332 331842 348384 331848
rect 350540 331900 350592 331906
rect 350540 331842 350592 331848
rect 350552 331226 350580 331842
rect 350540 331220 350592 331226
rect 350540 331162 350592 331168
rect 345756 330540 345808 330546
rect 345756 330482 345808 330488
rect 342260 285660 342312 285666
rect 342260 285602 342312 285608
rect 339500 285592 339552 285598
rect 353312 285569 353340 333254
rect 356072 288318 356100 333268
rect 358648 331906 358676 333268
rect 360212 333254 361238 333282
rect 358636 331900 358688 331906
rect 358636 331842 358688 331848
rect 360212 288386 360240 333254
rect 363800 331226 363828 333268
rect 366376 332586 366404 333268
rect 366364 332580 366416 332586
rect 366364 332522 366416 332528
rect 368952 331294 368980 333268
rect 371528 332722 371556 333268
rect 371516 332716 371568 332722
rect 371516 332658 371568 332664
rect 374104 331294 374132 333268
rect 376680 331430 376708 333268
rect 378152 333254 379270 333282
rect 376668 331424 376720 331430
rect 376668 331366 376720 331372
rect 368940 331288 368992 331294
rect 368940 331230 368992 331236
rect 373264 331288 373316 331294
rect 373264 331230 373316 331236
rect 374092 331288 374144 331294
rect 374092 331230 374144 331236
rect 363788 331220 363840 331226
rect 363788 331162 363840 331168
rect 373276 329118 373304 331230
rect 373264 329112 373316 329118
rect 373264 329054 373316 329060
rect 360200 288380 360252 288386
rect 360200 288322 360252 288328
rect 356060 288312 356112 288318
rect 356060 288254 356112 288260
rect 378152 287706 378180 333254
rect 381832 331294 381860 333268
rect 384408 332722 384436 333268
rect 386524 333254 386998 333282
rect 386524 332790 386552 333254
rect 386512 332784 386564 332790
rect 386512 332726 386564 332732
rect 383660 332716 383712 332722
rect 383660 332658 383712 332664
rect 384396 332716 384448 332722
rect 384396 332658 384448 332664
rect 382464 331424 382516 331430
rect 382464 331366 382516 331372
rect 379428 331288 379480 331294
rect 379428 331230 379480 331236
rect 381820 331288 381872 331294
rect 381820 331230 381872 331236
rect 379440 329769 379468 331230
rect 382476 329798 382504 331366
rect 382464 329792 382516 329798
rect 379426 329760 379482 329769
rect 382464 329734 382516 329740
rect 379426 329695 379482 329704
rect 378140 287700 378192 287706
rect 378140 287642 378192 287648
rect 339500 285534 339552 285540
rect 353298 285560 353354 285569
rect 353298 285495 353354 285504
rect 379440 284986 379468 329695
rect 383672 285122 383700 332658
rect 386328 331288 386380 331294
rect 386328 331230 386380 331236
rect 386340 329730 386368 331230
rect 386328 329724 386380 329730
rect 386328 329666 386380 329672
rect 386524 316034 386552 332726
rect 389560 329594 389588 333268
rect 392136 329662 392164 333268
rect 392124 329656 392176 329662
rect 392124 329598 392176 329604
rect 393228 329656 393280 329662
rect 393228 329598 393280 329604
rect 393320 329656 393372 329662
rect 393372 329604 393544 329610
rect 393320 329598 393544 329604
rect 389548 329588 389600 329594
rect 389548 329530 389600 329536
rect 390468 329588 390520 329594
rect 390468 329530 390520 329536
rect 386432 316006 386552 316034
rect 383660 285116 383712 285122
rect 383660 285058 383712 285064
rect 386432 285054 386460 316006
rect 390480 285190 390508 329530
rect 393240 285258 393268 329598
rect 393332 329594 393544 329598
rect 393332 329588 393556 329594
rect 393332 329582 393504 329588
rect 393504 329530 393556 329536
rect 394712 329458 394740 333268
rect 397288 332246 397316 333268
rect 399864 332518 399892 333268
rect 399852 332512 399904 332518
rect 399852 332454 399904 332460
rect 402440 332450 402468 333268
rect 402428 332444 402480 332450
rect 402428 332386 402480 332392
rect 397276 332240 397328 332246
rect 397276 332182 397328 332188
rect 405016 331906 405044 333268
rect 407592 332382 407620 333268
rect 407580 332376 407632 332382
rect 407580 332318 407632 332324
rect 410168 332314 410196 333268
rect 410156 332308 410208 332314
rect 410156 332250 410208 332256
rect 405004 331900 405056 331906
rect 405004 331842 405056 331848
rect 394700 329452 394752 329458
rect 394700 329394 394752 329400
rect 395988 329452 396040 329458
rect 395988 329394 396040 329400
rect 396000 285326 396028 329394
rect 412744 329186 412772 333268
rect 415320 332586 415348 333268
rect 416688 332852 416740 332858
rect 416688 332794 416740 332800
rect 415308 332580 415360 332586
rect 415308 332522 415360 332528
rect 412732 329180 412784 329186
rect 412732 329122 412784 329128
rect 395988 285320 396040 285326
rect 395988 285262 396040 285268
rect 393228 285252 393280 285258
rect 393228 285194 393280 285200
rect 390468 285184 390520 285190
rect 390468 285126 390520 285132
rect 386420 285048 386472 285054
rect 386420 284990 386472 284996
rect 329840 284980 329892 284986
rect 329840 284922 329892 284928
rect 379428 284980 379480 284986
rect 379428 284922 379480 284928
rect 416700 284374 416728 332794
rect 417896 331265 417924 333268
rect 418448 332518 418476 451246
rect 418540 332722 418568 456758
rect 418528 332716 418580 332722
rect 418528 332658 418580 332664
rect 418436 332512 418488 332518
rect 418436 332454 418488 332460
rect 418448 331294 418476 332454
rect 418632 332246 418660 457286
rect 418724 332450 418752 459575
rect 418804 458176 418856 458182
rect 418804 458118 418856 458124
rect 418816 332858 418844 458118
rect 419552 457178 419580 459614
rect 419736 459406 419764 460906
rect 419724 459400 419776 459406
rect 419724 459342 419776 459348
rect 419552 457150 419672 457178
rect 419540 457088 419592 457094
rect 419540 457030 419592 457036
rect 418804 332852 418856 332858
rect 418804 332794 418856 332800
rect 418712 332444 418764 332450
rect 418712 332386 418764 332392
rect 418620 332240 418672 332246
rect 418620 332182 418672 332188
rect 418632 331362 418660 332182
rect 418620 331356 418672 331362
rect 418620 331298 418672 331304
rect 418436 331288 418488 331294
rect 417882 331256 417938 331265
rect 418436 331230 418488 331236
rect 417882 331191 417938 331200
rect 417424 329792 417476 329798
rect 417424 329734 417476 329740
rect 417436 329526 417464 329734
rect 417424 329520 417476 329526
rect 417424 329462 417476 329468
rect 418724 316034 418752 332386
rect 419448 331900 419500 331906
rect 419448 331842 419500 331848
rect 418804 331152 418856 331158
rect 418804 331094 418856 331100
rect 418356 316006 418752 316034
rect 418252 285116 418304 285122
rect 418252 285058 418304 285064
rect 416688 284368 416740 284374
rect 416688 284310 416740 284316
rect 301412 206508 301464 206514
rect 301412 206450 301464 206456
rect 301148 204870 301360 204898
rect 301148 204105 301176 204870
rect 301424 204796 301452 206450
rect 371608 206304 371660 206310
rect 371608 206246 371660 206252
rect 371620 205306 371648 206246
rect 301332 204768 301452 204796
rect 301134 204096 301190 204105
rect 301134 204031 301190 204040
rect 300952 201340 301004 201346
rect 300952 201282 301004 201288
rect 300964 200666 300992 201282
rect 300952 200660 301004 200666
rect 300952 200602 301004 200608
rect 301148 76634 301176 204031
rect 301332 203998 301360 204768
rect 301412 204604 301464 204610
rect 301412 204546 301464 204552
rect 301320 203992 301372 203998
rect 301320 203934 301372 203940
rect 301136 76628 301188 76634
rect 301136 76570 301188 76576
rect 301332 74254 301360 203934
rect 301320 74248 301372 74254
rect 301320 74190 301372 74196
rect 300768 63504 300820 63510
rect 300768 63446 300820 63452
rect 300780 63034 300808 63446
rect 300768 63028 300820 63034
rect 300768 62970 300820 62976
rect 301424 62082 301452 204546
rect 301976 204241 302004 205292
rect 304552 204377 304580 205292
rect 304538 204368 304594 204377
rect 304538 204303 304594 204312
rect 307128 204270 307156 205292
rect 309048 204944 309100 204950
rect 309048 204886 309100 204892
rect 309060 204270 309088 204886
rect 307116 204264 307168 204270
rect 301962 204232 302018 204241
rect 307116 204206 307168 204212
rect 309048 204264 309100 204270
rect 309048 204206 309100 204212
rect 301962 204167 302018 204176
rect 302792 204060 302844 204066
rect 302792 204002 302844 204008
rect 302804 203862 302832 204002
rect 309704 203930 309732 205292
rect 312280 203998 312308 205292
rect 314856 204066 314884 205292
rect 317432 204134 317460 205292
rect 320008 204270 320036 205292
rect 319996 204264 320048 204270
rect 319996 204206 320048 204212
rect 317420 204128 317472 204134
rect 317420 204070 317472 204076
rect 314844 204060 314896 204066
rect 314844 204002 314896 204008
rect 322584 203998 322612 205292
rect 325160 204542 325188 205292
rect 325148 204536 325200 204542
rect 325148 204478 325200 204484
rect 327736 204474 327764 205292
rect 327724 204468 327776 204474
rect 327724 204410 327776 204416
rect 330312 204406 330340 205292
rect 330300 204400 330352 204406
rect 330300 204342 330352 204348
rect 332888 204202 332916 205292
rect 332876 204196 332928 204202
rect 332876 204138 332928 204144
rect 335464 204105 335492 205292
rect 335450 204096 335506 204105
rect 335450 204031 335506 204040
rect 312268 203992 312320 203998
rect 312268 203934 312320 203940
rect 319352 203992 319404 203998
rect 319352 203934 319404 203940
rect 322572 203992 322624 203998
rect 322572 203934 322624 203940
rect 309692 203924 309744 203930
rect 309692 203866 309744 203872
rect 302792 203856 302844 203862
rect 303528 203856 303580 203862
rect 302792 203798 302844 203804
rect 303526 203824 303528 203833
rect 303580 203824 303582 203833
rect 303526 203759 303582 203768
rect 319364 203561 319392 203934
rect 338040 203862 338068 205292
rect 339512 205278 340630 205306
rect 342272 205278 343206 205306
rect 371542 205292 371648 205306
rect 338028 203856 338080 203862
rect 338028 203798 338080 203804
rect 319350 203552 319406 203561
rect 319350 203487 319406 203496
rect 303528 158704 303580 158710
rect 303526 158672 303528 158681
rect 303580 158672 303582 158681
rect 303526 158607 303582 158616
rect 339512 158574 339540 205278
rect 342272 158642 342300 205278
rect 345768 201346 345796 205292
rect 348344 204270 348372 205292
rect 350920 204270 350948 205292
rect 353496 204338 353524 205292
rect 353484 204332 353536 204338
rect 353484 204274 353536 204280
rect 348332 204264 348384 204270
rect 348332 204206 348384 204212
rect 350908 204264 350960 204270
rect 350908 204206 350960 204212
rect 345756 201340 345808 201346
rect 345756 201282 345808 201288
rect 348344 200114 348372 204206
rect 352564 203584 352616 203590
rect 352564 203526 352616 203532
rect 348344 200086 348464 200114
rect 342260 158636 342312 158642
rect 342260 158578 342312 158584
rect 339500 158568 339552 158574
rect 339500 158510 339552 158516
rect 348436 158030 348464 200086
rect 352576 158710 352604 203526
rect 356072 201414 356100 205292
rect 358648 203590 358676 205292
rect 358636 203584 358688 203590
rect 358636 203526 358688 203532
rect 361224 201482 361252 205292
rect 363800 201482 363828 205292
rect 365628 204604 365680 204610
rect 365628 204546 365680 204552
rect 365640 204202 365668 204546
rect 365628 204196 365680 204202
rect 365628 204138 365680 204144
rect 366376 203114 366404 205292
rect 368952 204270 368980 205292
rect 371528 205278 371648 205292
rect 368940 204264 368992 204270
rect 368940 204206 368992 204212
rect 371528 204202 371556 205278
rect 372620 204740 372672 204746
rect 372620 204682 372672 204688
rect 372632 204270 372660 204682
rect 374104 204338 374132 205292
rect 374092 204332 374144 204338
rect 374092 204274 374144 204280
rect 372620 204264 372672 204270
rect 372620 204206 372672 204212
rect 371516 204196 371568 204202
rect 371516 204138 371568 204144
rect 376680 203182 376708 205292
rect 378152 205278 379270 205306
rect 376668 203176 376720 203182
rect 376668 203118 376720 203124
rect 366364 203108 366416 203114
rect 366364 203050 366416 203056
rect 370136 203108 370188 203114
rect 370136 203050 370188 203056
rect 361212 201476 361264 201482
rect 361212 201418 361264 201424
rect 363788 201476 363840 201482
rect 363788 201418 363840 201424
rect 370148 201414 370176 203050
rect 356060 201408 356112 201414
rect 356060 201350 356112 201356
rect 370136 201408 370188 201414
rect 370136 201350 370188 201356
rect 378152 164898 378180 205278
rect 381832 202978 381860 205292
rect 384408 204406 384436 205292
rect 386984 204474 387012 205292
rect 389560 204542 389588 205292
rect 392136 204610 392164 205292
rect 394712 204678 394740 205292
rect 394700 204672 394752 204678
rect 394700 204614 394752 204620
rect 392124 204604 392176 204610
rect 392124 204546 392176 204552
rect 389548 204536 389600 204542
rect 389548 204478 389600 204484
rect 386972 204468 387024 204474
rect 386972 204410 387024 204416
rect 384396 204400 384448 204406
rect 384396 204342 384448 204348
rect 397288 204270 397316 205292
rect 397276 204264 397328 204270
rect 397276 204206 397328 204212
rect 399864 203930 399892 205292
rect 402440 204202 402468 205292
rect 402428 204196 402480 204202
rect 402428 204138 402480 204144
rect 405016 204066 405044 205292
rect 405004 204060 405056 204066
rect 405004 204002 405056 204008
rect 407592 203998 407620 205292
rect 410168 204134 410196 205292
rect 411260 204264 411312 204270
rect 411260 204206 411312 204212
rect 410156 204128 410208 204134
rect 410156 204070 410208 204076
rect 407580 203992 407632 203998
rect 407580 203934 407632 203940
rect 399852 203924 399904 203930
rect 399852 203866 399904 203872
rect 411272 203561 411300 204206
rect 411258 203552 411314 203561
rect 411258 203487 411314 203496
rect 382648 203176 382700 203182
rect 382648 203118 382700 203124
rect 381820 202972 381872 202978
rect 381820 202914 381872 202920
rect 382660 201346 382688 203118
rect 385408 202972 385460 202978
rect 385408 202914 385460 202920
rect 382648 201340 382700 201346
rect 382648 201282 382700 201288
rect 385420 201278 385448 202914
rect 412744 202910 412772 205292
rect 415320 204270 415348 205292
rect 417910 205278 418108 205306
rect 415308 204264 415360 204270
rect 415308 204206 415360 204212
rect 416780 204264 416832 204270
rect 416780 204206 416832 204212
rect 416792 204105 416820 204206
rect 416778 204096 416834 204105
rect 416778 204031 416834 204040
rect 418080 202994 418108 205278
rect 418264 204746 418292 285058
rect 418252 204740 418304 204746
rect 418252 204682 418304 204688
rect 418356 204202 418384 316006
rect 418528 284368 418580 284374
rect 418528 284310 418580 284316
rect 418436 204740 418488 204746
rect 418436 204682 418488 204688
rect 418448 204406 418476 204682
rect 418436 204400 418488 204406
rect 418436 204342 418488 204348
rect 418344 204196 418396 204202
rect 418344 204138 418396 204144
rect 418080 202966 418292 202994
rect 412732 202904 412784 202910
rect 412732 202846 412784 202852
rect 385408 201272 385460 201278
rect 385408 201214 385460 201220
rect 378140 164892 378192 164898
rect 378140 164834 378192 164840
rect 352564 158704 352616 158710
rect 352564 158646 352616 158652
rect 348424 158024 348476 158030
rect 348424 157966 348476 157972
rect 306656 78668 306708 78674
rect 306656 78610 306708 78616
rect 302054 78568 302110 78577
rect 301990 78526 302054 78554
rect 302054 78503 302110 78512
rect 306668 77330 306696 78610
rect 410432 78328 410484 78334
rect 407132 78266 407896 78282
rect 409892 78276 410432 78282
rect 409892 78270 410484 78276
rect 407132 78260 407908 78266
rect 407132 78254 407856 78260
rect 405280 78192 405332 78198
rect 327368 78130 327750 78146
rect 399878 78130 400168 78146
rect 404372 78140 405280 78146
rect 404372 78134 405332 78140
rect 327172 78124 327224 78130
rect 327172 78066 327224 78072
rect 327356 78124 327750 78130
rect 327408 78118 327750 78124
rect 398840 78124 398892 78130
rect 327356 78066 327408 78072
rect 399878 78124 400180 78130
rect 399878 78118 400128 78124
rect 398840 78066 398892 78072
rect 400128 78066 400180 78072
rect 404372 78118 405320 78134
rect 304552 75954 304580 77316
rect 306668 77302 307142 77330
rect 304540 75948 304592 75954
rect 304540 75890 304592 75896
rect 305368 72548 305420 72554
rect 305368 72490 305420 72496
rect 303712 69760 303764 69766
rect 303712 69702 303764 69708
rect 302240 68400 302292 68406
rect 302240 68342 302292 68348
rect 301412 62076 301464 62082
rect 301412 62018 301464 62024
rect 301424 61606 301452 62018
rect 301412 61600 301464 61606
rect 301412 61542 301464 61548
rect 302252 54754 302280 68342
rect 302332 60648 302384 60654
rect 302330 60616 302332 60625
rect 302384 60616 302386 60625
rect 302330 60551 302386 60560
rect 302344 59430 302372 60551
rect 302332 59424 302384 59430
rect 302332 59366 302384 59372
rect 303724 54754 303752 69702
rect 305380 54754 305408 72490
rect 306668 64874 306696 77302
rect 309704 74526 309732 77316
rect 312294 77302 312584 77330
rect 314870 77302 315344 77330
rect 317446 77302 318104 77330
rect 309692 74520 309744 74526
rect 309692 74462 309744 74468
rect 308680 73840 308732 73846
rect 308680 73782 308732 73788
rect 306392 64846 306696 64874
rect 306392 57866 306420 64846
rect 307116 58812 307168 58818
rect 307116 58754 307168 58760
rect 306380 57860 306432 57866
rect 306380 57802 306432 57808
rect 307128 56982 307156 58754
rect 307392 57656 307444 57662
rect 307392 57598 307444 57604
rect 307116 56976 307168 56982
rect 307116 56918 307168 56924
rect 292132 54726 292514 54754
rect 293972 54726 294170 54754
rect 295444 54726 295826 54754
rect 297100 54726 297482 54754
rect 298756 54726 299138 54754
rect 300412 54726 300794 54754
rect 302252 54726 302450 54754
rect 303724 54726 304106 54754
rect 305380 54726 305762 54754
rect 307404 54740 307432 57598
rect 308692 54754 308720 73782
rect 309704 73234 309732 74462
rect 312556 74254 312584 77302
rect 315316 74322 315344 77302
rect 318076 74390 318104 77302
rect 319456 77302 320022 77330
rect 319456 74458 319484 77302
rect 319444 74452 319496 74458
rect 319444 74394 319496 74400
rect 318064 74384 318116 74390
rect 318064 74326 318116 74332
rect 315304 74316 315356 74322
rect 315304 74258 315356 74264
rect 312544 74248 312596 74254
rect 312544 74190 312596 74196
rect 309692 73228 309744 73234
rect 309692 73170 309744 73176
rect 311164 73228 311216 73234
rect 311164 73170 311216 73176
rect 311176 57934 311204 73170
rect 311164 57928 311216 57934
rect 311164 57870 311216 57876
rect 312556 57866 312584 74190
rect 314016 57928 314068 57934
rect 314016 57870 314068 57876
rect 312360 57860 312412 57866
rect 312360 57802 312412 57808
rect 312544 57860 312596 57866
rect 312544 57802 312596 57808
rect 310704 56976 310756 56982
rect 310704 56918 310756 56924
rect 308692 54726 309074 54754
rect 310716 54740 310744 56918
rect 312372 54740 312400 57802
rect 314028 54740 314056 57870
rect 315316 56642 315344 74258
rect 318076 57934 318104 74326
rect 319456 57934 319484 74394
rect 322584 74186 322612 77316
rect 325160 75818 325188 77316
rect 322940 75812 322992 75818
rect 322940 75754 322992 75760
rect 325148 75812 325200 75818
rect 325148 75754 325200 75760
rect 327080 75812 327132 75818
rect 327080 75754 327132 75760
rect 322952 75614 322980 75754
rect 322940 75608 322992 75614
rect 322940 75550 322992 75556
rect 322952 74534 322980 75550
rect 327092 75546 327120 75754
rect 327080 75540 327132 75546
rect 327080 75482 327132 75488
rect 322952 74506 323624 74534
rect 322572 74180 322624 74186
rect 322572 74122 322624 74128
rect 322584 73234 322612 74122
rect 321928 73228 321980 73234
rect 321928 73170 321980 73176
rect 322572 73228 322624 73234
rect 322572 73170 322624 73176
rect 318064 57928 318116 57934
rect 318064 57870 318116 57876
rect 318984 57928 319036 57934
rect 318984 57870 319036 57876
rect 319444 57928 319496 57934
rect 319444 57870 319496 57876
rect 320640 57928 320692 57934
rect 320640 57870 320692 57876
rect 315672 57860 315724 57866
rect 315672 57802 315724 57808
rect 315304 56636 315356 56642
rect 315304 56578 315356 56584
rect 315684 54740 315712 57802
rect 317328 56636 317380 56642
rect 317328 56578 317380 56584
rect 317340 54740 317368 56578
rect 318996 54740 319024 57870
rect 320652 54740 320680 57870
rect 321940 54754 321968 73170
rect 322940 62960 322992 62966
rect 322940 62902 322992 62908
rect 322952 57594 322980 62902
rect 322940 57588 322992 57594
rect 322940 57530 322992 57536
rect 323596 54754 323624 74506
rect 325608 56636 325660 56642
rect 325608 56578 325660 56584
rect 321940 54726 322322 54754
rect 323596 54726 323978 54754
rect 325620 54740 325648 56578
rect 327092 54754 327120 75482
rect 327184 56642 327212 78066
rect 330484 78056 330536 78062
rect 330484 77998 330536 78004
rect 332600 78056 332652 78062
rect 396172 78056 396224 78062
rect 332652 78004 332902 78010
rect 332600 77998 332902 78004
rect 397368 78056 397420 78062
rect 396172 77998 396224 78004
rect 397302 78004 397368 78010
rect 397302 77998 397420 78004
rect 329932 76628 329984 76634
rect 329932 76570 329984 76576
rect 329944 75750 329972 76570
rect 330312 75818 330340 77316
rect 330300 75812 330352 75818
rect 330300 75754 330352 75760
rect 329932 75744 329984 75750
rect 329932 75686 329984 75692
rect 329944 74534 329972 75686
rect 329944 74506 330248 74534
rect 328920 57928 328972 57934
rect 328920 57870 328972 57876
rect 327172 56636 327224 56642
rect 327172 56578 327224 56584
rect 327092 54726 327290 54754
rect 328932 54740 328960 57870
rect 330220 54754 330248 74506
rect 330496 57934 330524 77998
rect 332612 77982 332902 77998
rect 369860 77988 369912 77994
rect 369860 77930 369912 77936
rect 393320 77988 393372 77994
rect 393320 77930 393372 77936
rect 348608 77376 348660 77382
rect 348358 77324 348608 77330
rect 348358 77318 348660 77324
rect 350540 77376 350592 77382
rect 350592 77324 350934 77330
rect 350540 77318 350934 77324
rect 348358 77316 348648 77318
rect 333978 76664 334034 76673
rect 333978 76599 334034 76608
rect 333992 75886 334020 76599
rect 333980 75880 334032 75886
rect 333980 75822 334032 75828
rect 334624 75880 334676 75886
rect 334624 75822 334676 75828
rect 332600 75472 332652 75478
rect 332600 75414 332652 75420
rect 332612 74534 332640 75414
rect 332612 74506 333560 74534
rect 330484 57928 330536 57934
rect 330484 57870 330536 57876
rect 332232 57792 332284 57798
rect 332232 57734 332284 57740
rect 330220 54726 330602 54754
rect 332244 54740 332272 57734
rect 333532 54754 333560 74506
rect 334636 57798 334664 75822
rect 335464 75750 335492 77316
rect 336740 76560 336792 76566
rect 336740 76502 336792 76508
rect 336752 75818 336780 76502
rect 338040 75886 338068 77316
rect 338028 75880 338080 75886
rect 338028 75822 338080 75828
rect 336740 75812 336792 75818
rect 336740 75754 336792 75760
rect 335452 75744 335504 75750
rect 335452 75686 335504 75692
rect 335360 75200 335412 75206
rect 335360 75142 335412 75148
rect 334624 57792 334676 57798
rect 334624 57734 334676 57740
rect 335372 54754 335400 75142
rect 336752 74534 336780 75754
rect 340616 75478 340644 77316
rect 340604 75472 340656 75478
rect 340604 75414 340656 75420
rect 343192 75206 343220 77316
rect 345768 75886 345796 77316
rect 348344 77302 348648 77316
rect 350552 77302 350934 77318
rect 353312 77302 353510 77330
rect 345756 75880 345808 75886
rect 345756 75822 345808 75828
rect 343180 75200 343232 75206
rect 343180 75142 343232 75148
rect 336752 74506 336872 74534
rect 336844 54754 336872 74506
rect 346766 73808 346822 73817
rect 346766 73743 346822 73752
rect 345112 71120 345164 71126
rect 345112 71062 345164 71068
rect 338488 71052 338540 71058
rect 338488 70994 338540 71000
rect 338500 54754 338528 70994
rect 341800 62892 341852 62898
rect 341800 62834 341852 62840
rect 340144 62824 340196 62830
rect 340144 62766 340196 62772
rect 340236 62824 340288 62830
rect 340236 62766 340288 62772
rect 340156 54754 340184 62766
rect 340248 57526 340276 62766
rect 340236 57520 340288 57526
rect 340236 57462 340288 57468
rect 341812 54754 341840 62834
rect 343640 58676 343692 58682
rect 343640 58618 343692 58624
rect 343652 54754 343680 58618
rect 345124 54754 345152 71062
rect 346780 54754 346808 73743
rect 348344 71262 348372 77302
rect 351184 75200 351236 75206
rect 351184 75142 351236 75148
rect 348332 71256 348384 71262
rect 348332 71198 348384 71204
rect 348424 66904 348476 66910
rect 348424 66846 348476 66852
rect 348436 54754 348464 66846
rect 350080 64184 350132 64190
rect 350080 64126 350132 64132
rect 350092 54754 350120 64126
rect 351196 57458 351224 75142
rect 351920 64252 351972 64258
rect 351920 64194 351972 64200
rect 351184 57452 351236 57458
rect 351184 57394 351236 57400
rect 351932 54754 351960 64194
rect 353312 60722 353340 77302
rect 355046 73944 355102 73953
rect 355046 73879 355102 73888
rect 353392 64320 353444 64326
rect 353392 64262 353444 64268
rect 353300 60716 353352 60722
rect 353300 60658 353352 60664
rect 353404 54754 353432 64262
rect 355060 54754 355088 73879
rect 356072 66230 356100 77316
rect 357544 77302 358662 77330
rect 360304 77302 361238 77330
rect 357440 72480 357492 72486
rect 357440 72422 357492 72428
rect 356704 66972 356756 66978
rect 356704 66914 356756 66920
rect 356060 66224 356112 66230
rect 356060 66166 356112 66172
rect 356716 54754 356744 66914
rect 357452 55214 357480 72422
rect 357544 60654 357572 77302
rect 360200 69692 360252 69698
rect 360200 69634 360252 69640
rect 357532 60648 357584 60654
rect 357532 60590 357584 60596
rect 357452 55186 358400 55214
rect 358372 54754 358400 55186
rect 360212 54754 360240 69634
rect 360304 63510 360332 77302
rect 363800 75886 363828 77316
rect 363788 75880 363840 75886
rect 363788 75822 363840 75828
rect 363800 72622 363828 75822
rect 366376 74497 366404 77316
rect 368952 74526 368980 77316
rect 369872 74534 369900 77930
rect 371146 77888 371202 77897
rect 371202 77846 371280 77874
rect 371146 77823 371202 77832
rect 368940 74520 368992 74526
rect 366362 74488 366418 74497
rect 369872 74506 369992 74534
rect 368940 74462 368992 74468
rect 366362 74423 366418 74432
rect 363788 72616 363840 72622
rect 363788 72558 363840 72564
rect 361672 68332 361724 68338
rect 361672 68274 361724 68280
rect 360292 63504 360344 63510
rect 360292 63446 360344 63452
rect 361684 54754 361712 68274
rect 366376 64394 366404 74423
rect 368952 69834 368980 74462
rect 368940 69828 368992 69834
rect 368940 69770 368992 69776
rect 368480 68536 368532 68542
rect 368480 68478 368532 68484
rect 366364 64388 366416 64394
rect 366364 64330 366416 64336
rect 366640 61464 366692 61470
rect 366640 61406 366692 61412
rect 364984 60104 365036 60110
rect 364984 60046 365036 60052
rect 363696 57588 363748 57594
rect 363696 57530 363748 57536
rect 333532 54726 333914 54754
rect 335372 54726 335570 54754
rect 336844 54726 337226 54754
rect 338500 54726 338882 54754
rect 340156 54726 340538 54754
rect 341812 54726 342194 54754
rect 343652 54726 343850 54754
rect 345124 54726 345506 54754
rect 346780 54726 347162 54754
rect 348436 54726 348818 54754
rect 350092 54726 350474 54754
rect 351932 54726 352130 54754
rect 353404 54726 353786 54754
rect 355060 54726 355442 54754
rect 356716 54726 357098 54754
rect 358372 54726 358754 54754
rect 360212 54726 360410 54754
rect 361684 54726 362066 54754
rect 363708 54740 363736 57530
rect 364996 54754 365024 60046
rect 366652 54754 366680 61406
rect 368492 54754 368520 68478
rect 369964 54754 369992 74506
rect 371252 55214 371280 77846
rect 371344 77302 371542 77330
rect 371344 62082 371372 77302
rect 373998 76800 374054 76809
rect 373998 76735 374054 76744
rect 372618 76664 372674 76673
rect 372618 76599 372674 76608
rect 372632 74534 372660 76599
rect 372632 74506 373304 74534
rect 371332 62076 371384 62082
rect 371332 62018 371384 62024
rect 371252 55186 371648 55214
rect 371620 54754 371648 55186
rect 373276 54754 373304 74506
rect 374012 55214 374040 76735
rect 374104 74361 374132 77316
rect 376680 74458 376708 77316
rect 378232 76628 378284 76634
rect 378232 76570 378284 76576
rect 376760 76560 376812 76566
rect 376760 76502 376812 76508
rect 376668 74452 376720 74458
rect 376668 74394 376720 74400
rect 374090 74352 374146 74361
rect 374090 74287 374146 74296
rect 374642 74352 374698 74361
rect 374642 74287 374698 74296
rect 374656 60042 374684 74287
rect 376680 73234 376708 74394
rect 376024 73228 376076 73234
rect 376024 73170 376076 73176
rect 376668 73228 376720 73234
rect 376668 73170 376720 73176
rect 376036 61402 376064 73170
rect 376024 61396 376076 61402
rect 376024 61338 376076 61344
rect 374644 60036 374696 60042
rect 374644 59978 374696 59984
rect 374012 55186 374960 55214
rect 374932 54754 374960 55186
rect 376772 54754 376800 76502
rect 378244 54754 378272 76570
rect 379256 75410 379284 77316
rect 381556 77302 381846 77330
rect 379244 75404 379296 75410
rect 379244 75346 379296 75352
rect 379520 75404 379572 75410
rect 379520 75346 379572 75352
rect 379532 74534 379560 75346
rect 381556 74534 381584 77302
rect 384408 75342 384436 77316
rect 386510 76528 386566 76537
rect 386510 76463 386566 76472
rect 384948 75744 385000 75750
rect 384948 75686 385000 75692
rect 384960 75342 384988 75686
rect 384396 75336 384448 75342
rect 384396 75278 384448 75284
rect 384948 75336 385000 75342
rect 384948 75278 385000 75284
rect 379532 74506 379928 74534
rect 379900 54754 379928 74506
rect 381464 74506 381584 74534
rect 381464 74390 381492 74506
rect 381452 74384 381504 74390
rect 381452 74326 381504 74332
rect 381464 65550 381492 74326
rect 381544 71188 381596 71194
rect 381544 71130 381596 71136
rect 381452 65544 381504 65550
rect 381452 65486 381504 65492
rect 381556 54754 381584 71130
rect 383568 57384 383620 57390
rect 383568 57326 383620 57332
rect 364996 54726 365378 54754
rect 366652 54726 367034 54754
rect 368492 54726 368690 54754
rect 369964 54726 370346 54754
rect 371620 54726 372002 54754
rect 373276 54726 373658 54754
rect 374932 54726 375314 54754
rect 376772 54726 376970 54754
rect 378244 54726 378626 54754
rect 379900 54726 380282 54754
rect 381556 54726 381938 54754
rect 383580 54740 383608 57326
rect 385224 57316 385276 57322
rect 385224 57258 385276 57264
rect 385236 54740 385264 57258
rect 386524 54754 386552 76463
rect 386984 75818 387012 77316
rect 386972 75812 387024 75818
rect 386972 75754 387024 75760
rect 386984 75206 387012 75754
rect 389560 75682 389588 77316
rect 392150 77302 392532 77330
rect 390560 76696 390612 76702
rect 390560 76638 390612 76644
rect 389548 75676 389600 75682
rect 389548 75618 389600 75624
rect 389560 75274 389588 75618
rect 389548 75268 389600 75274
rect 389548 75210 389600 75216
rect 386972 75200 387024 75206
rect 386972 75142 387024 75148
rect 390572 74534 390600 76638
rect 392504 74534 392532 77302
rect 390572 74506 391520 74534
rect 392504 74506 392624 74534
rect 388536 57248 388588 57254
rect 388536 57190 388588 57196
rect 390192 57248 390244 57254
rect 390192 57190 390244 57196
rect 386524 54726 386906 54754
rect 388548 54740 388576 57190
rect 390204 54740 390232 57190
rect 391492 54754 391520 74506
rect 392596 74322 392624 74506
rect 392584 74316 392636 74322
rect 392584 74258 392636 74264
rect 392596 62830 392624 74258
rect 392584 62824 392636 62830
rect 392584 62766 392636 62772
rect 393332 54754 393360 77930
rect 394712 74254 394740 77316
rect 396080 75200 396132 75206
rect 396080 75142 396132 75148
rect 394700 74248 394752 74254
rect 394700 74190 394752 74196
rect 394712 73574 394740 74190
rect 394700 73568 394752 73574
rect 394700 73510 394752 73516
rect 395344 73568 395396 73574
rect 395344 73510 395396 73516
rect 395356 61538 395384 73510
rect 396092 64874 396120 75142
rect 396184 67046 396212 77998
rect 397302 77982 397408 77998
rect 396172 67040 396224 67046
rect 396172 66982 396224 66988
rect 398852 65618 398880 78066
rect 402256 77302 402454 77330
rect 402256 74186 402284 77302
rect 402244 74180 402296 74186
rect 402244 74122 402296 74128
rect 398840 65612 398892 65618
rect 398840 65554 398892 65560
rect 396092 64846 396488 64874
rect 395344 61532 395396 61538
rect 395344 61474 395396 61480
rect 395160 57316 395212 57322
rect 395160 57258 395212 57264
rect 391492 54726 391874 54754
rect 393332 54726 393530 54754
rect 395172 54740 395200 57258
rect 396460 54754 396488 64846
rect 402256 58886 402284 74122
rect 404372 68474 404400 78118
rect 407132 69902 407160 78254
rect 407856 78202 407908 78208
rect 409892 78254 410472 78270
rect 409892 72690 409920 78254
rect 412744 75410 412772 77316
rect 412732 75404 412784 75410
rect 412732 75346 412784 75352
rect 415320 74118 415348 77316
rect 417896 75206 417924 77316
rect 417884 75200 417936 75206
rect 417884 75142 417936 75148
rect 415308 74112 415360 74118
rect 415308 74054 415360 74060
rect 415320 73234 415348 74054
rect 414664 73228 414716 73234
rect 414664 73170 414716 73176
rect 415308 73228 415360 73234
rect 415308 73170 415360 73176
rect 409880 72684 409932 72690
rect 409880 72626 409932 72632
rect 407120 69896 407172 69902
rect 407120 69838 407172 69844
rect 404360 68468 404412 68474
rect 404360 68410 404412 68416
rect 402244 58880 402296 58886
rect 402244 58822 402296 58828
rect 414676 58750 414704 73170
rect 414664 58744 414716 58750
rect 414664 58686 414716 58692
rect 418264 57322 418292 202966
rect 418356 74186 418384 204138
rect 418448 75750 418476 204342
rect 418540 201414 418568 284310
rect 418816 203998 418844 331094
rect 419460 331022 419488 331842
rect 419448 331016 419500 331022
rect 419448 330958 419500 330964
rect 419460 204202 419488 330958
rect 419552 329458 419580 457030
rect 419644 332382 419672 457150
rect 419736 345014 419764 459342
rect 419816 458992 419868 458998
rect 419816 458934 419868 458940
rect 419828 457094 419856 458934
rect 419816 457088 419868 457094
rect 419816 457030 419868 457036
rect 419736 344986 419948 345014
rect 419632 332376 419684 332382
rect 419632 332318 419684 332324
rect 419644 331158 419672 332318
rect 419920 332314 419948 344986
rect 419908 332308 419960 332314
rect 419908 332250 419960 332256
rect 419632 331152 419684 331158
rect 419632 331094 419684 331100
rect 419816 329792 419868 329798
rect 419816 329734 419868 329740
rect 419540 329452 419592 329458
rect 419540 329394 419592 329400
rect 419828 329118 419856 329734
rect 419816 329112 419868 329118
rect 419816 329054 419868 329060
rect 419828 209774 419856 329054
rect 419552 209746 419856 209774
rect 419552 205086 419580 209746
rect 419540 205080 419592 205086
rect 419540 205022 419592 205028
rect 419448 204196 419500 204202
rect 419448 204138 419500 204144
rect 418804 203992 418856 203998
rect 418804 203934 418856 203940
rect 418528 201408 418580 201414
rect 418528 201350 418580 201356
rect 418436 75744 418488 75750
rect 418436 75686 418488 75692
rect 418540 74497 418568 201350
rect 418816 200114 418844 203934
rect 418632 200086 418844 200114
rect 418632 78266 418660 200086
rect 418620 78260 418672 78266
rect 418620 78202 418672 78208
rect 419552 74526 419580 205022
rect 419920 204626 419948 332250
rect 420840 331401 420868 470562
rect 420932 458998 420960 583374
rect 421380 583296 421432 583302
rect 421380 583238 421432 583244
rect 421196 583228 421248 583234
rect 421196 583170 421248 583176
rect 421104 541884 421156 541890
rect 421104 541826 421156 541832
rect 421116 463078 421144 541826
rect 421208 465458 421236 583170
rect 421288 541680 421340 541686
rect 421288 541622 421340 541628
rect 421196 465452 421248 465458
rect 421196 465394 421248 465400
rect 421300 465338 421328 541622
rect 421208 465310 421328 465338
rect 421104 463072 421156 463078
rect 421104 463014 421156 463020
rect 421208 463010 421236 465310
rect 421288 465248 421340 465254
rect 421288 465190 421340 465196
rect 421196 463004 421248 463010
rect 421196 462946 421248 462952
rect 421208 462398 421236 462946
rect 421196 462392 421248 462398
rect 421196 462334 421248 462340
rect 421104 462324 421156 462330
rect 421104 462266 421156 462272
rect 421012 460964 421064 460970
rect 421012 460906 421064 460912
rect 420920 458992 420972 458998
rect 420920 458934 420972 458940
rect 420920 458856 420972 458862
rect 420920 458798 420972 458804
rect 420932 458114 420960 458798
rect 420920 458108 420972 458114
rect 420920 458050 420972 458056
rect 420826 331392 420882 331401
rect 420092 331356 420144 331362
rect 420826 331327 420882 331336
rect 420092 331298 420144 331304
rect 420000 331288 420052 331294
rect 420000 331230 420052 331236
rect 419644 204598 419948 204626
rect 419644 204270 419672 204598
rect 420012 204490 420040 331230
rect 419736 204462 420040 204490
rect 419632 204264 419684 204270
rect 419632 204206 419684 204212
rect 419644 78334 419672 204206
rect 419736 203930 419764 204462
rect 420104 204354 420132 331298
rect 421024 331022 421052 460906
rect 421116 332586 421144 462266
rect 421300 462210 421328 465190
rect 421208 462182 421328 462210
rect 421208 460986 421236 462182
rect 421392 461145 421420 583238
rect 421378 461136 421434 461145
rect 421378 461071 421434 461080
rect 421286 461000 421342 461009
rect 421208 460958 421286 460986
rect 421208 332790 421236 460958
rect 421286 460935 421342 460944
rect 421472 459264 421524 459270
rect 421472 459206 421524 459212
rect 421196 332784 421248 332790
rect 421196 332726 421248 332732
rect 421104 332580 421156 332586
rect 421104 332522 421156 332528
rect 421012 331016 421064 331022
rect 421012 330958 421064 330964
rect 421012 285184 421064 285190
rect 421012 285126 421064 285132
rect 421024 209774 421052 285126
rect 420932 209746 421052 209774
rect 420932 205426 420960 209746
rect 420920 205420 420972 205426
rect 420920 205362 420972 205368
rect 420932 204542 420960 205362
rect 420920 204536 420972 204542
rect 420920 204478 420972 204484
rect 419828 204326 420132 204354
rect 419724 203924 419776 203930
rect 419724 203866 419776 203872
rect 419632 78328 419684 78334
rect 419632 78270 419684 78276
rect 419736 78130 419764 203866
rect 419828 203561 419856 204326
rect 419908 204196 419960 204202
rect 419908 204138 419960 204144
rect 419814 203552 419870 203561
rect 419814 203487 419870 203496
rect 419724 78124 419776 78130
rect 419724 78066 419776 78072
rect 419828 78062 419856 203487
rect 419920 78198 419948 204138
rect 421116 204105 421144 332522
rect 421196 285048 421248 285054
rect 421196 284990 421248 284996
rect 421208 204474 421236 284990
rect 421196 204468 421248 204474
rect 421196 204410 421248 204416
rect 421102 204096 421158 204105
rect 421102 204031 421158 204040
rect 419908 78192 419960 78198
rect 419908 78134 419960 78140
rect 419816 78056 419868 78062
rect 419816 77998 419868 78004
rect 419540 74520 419592 74526
rect 418526 74488 418582 74497
rect 419540 74462 419592 74468
rect 418526 74423 418582 74432
rect 418344 74180 418396 74186
rect 418344 74122 418396 74128
rect 421116 74118 421144 204031
rect 421208 75818 421236 204410
rect 421380 204332 421432 204338
rect 421380 204274 421432 204280
rect 421288 202904 421340 202910
rect 421288 202846 421340 202852
rect 421300 76634 421328 202846
rect 421288 76628 421340 76634
rect 421288 76570 421340 76576
rect 421196 75812 421248 75818
rect 421196 75754 421248 75760
rect 421392 74361 421420 204274
rect 421484 76702 421512 459206
rect 421564 458108 421616 458114
rect 421564 458050 421616 458056
rect 421576 329798 421604 458050
rect 421564 329792 421616 329798
rect 421564 329734 421616 329740
rect 421564 204944 421616 204950
rect 421564 204886 421616 204892
rect 421576 204338 421604 204886
rect 421564 204332 421616 204338
rect 421564 204274 421616 204280
rect 421472 76696 421524 76702
rect 421472 76638 421524 76644
rect 421378 74352 421434 74361
rect 421378 74287 421434 74296
rect 421104 74112 421156 74118
rect 421104 74054 421156 74060
rect 418252 57316 418304 57322
rect 418252 57258 418304 57264
rect 422312 57254 422340 585103
rect 422576 583364 422628 583370
rect 422576 583306 422628 583312
rect 422392 541816 422444 541822
rect 422392 541758 422444 541764
rect 422404 460834 422432 541758
rect 422484 541748 422536 541754
rect 422484 541690 422536 541696
rect 422496 460902 422524 541690
rect 422484 460896 422536 460902
rect 422484 460838 422536 460844
rect 422392 460828 422444 460834
rect 422392 460770 422444 460776
rect 422404 459610 422432 460770
rect 422392 459604 422444 459610
rect 422392 459546 422444 459552
rect 422390 331256 422446 331265
rect 422390 331191 422446 331200
rect 422404 77994 422432 331191
rect 422496 329769 422524 460838
rect 422588 459474 422616 583306
rect 423680 583160 423732 583166
rect 423680 583102 423732 583108
rect 422666 461000 422722 461009
rect 422666 460935 422722 460944
rect 422576 459468 422628 459474
rect 422576 459410 422628 459416
rect 422482 329760 422538 329769
rect 422482 329695 422538 329704
rect 422588 329594 422616 459410
rect 422680 329662 422708 460935
rect 423692 458114 423720 583102
rect 425152 583092 425204 583098
rect 425152 583034 425204 583040
rect 423864 583024 423916 583030
rect 423864 582966 423916 582972
rect 423772 462392 423824 462398
rect 423772 462334 423824 462340
rect 423680 458108 423732 458114
rect 423680 458050 423732 458056
rect 423784 332654 423812 462334
rect 423876 459338 423904 582966
rect 425060 463072 425112 463078
rect 425060 463014 425112 463020
rect 423956 459604 424008 459610
rect 423956 459546 424008 459552
rect 423864 459332 423916 459338
rect 423864 459274 423916 459280
rect 423772 332648 423824 332654
rect 423772 332590 423824 332596
rect 423876 331106 423904 459274
rect 423784 331090 423904 331106
rect 423772 331084 423904 331090
rect 423824 331078 423904 331084
rect 423772 331026 423824 331032
rect 422668 329656 422720 329662
rect 422668 329598 422720 329604
rect 422576 329588 422628 329594
rect 422576 329530 422628 329536
rect 423680 329520 423732 329526
rect 423680 329462 423732 329468
rect 422484 329180 422536 329186
rect 422484 329122 422536 329128
rect 422392 77988 422444 77994
rect 422392 77930 422444 77936
rect 422496 76566 422524 329122
rect 422576 285252 422628 285258
rect 422576 285194 422628 285200
rect 422588 204610 422616 285194
rect 422668 205420 422720 205426
rect 422668 205362 422720 205368
rect 422576 204604 422628 204610
rect 422576 204546 422628 204552
rect 422484 76560 422536 76566
rect 422484 76502 422536 76508
rect 422680 75682 422708 205362
rect 423692 201346 423720 329462
rect 423784 209774 423812 331026
rect 423968 329526 423996 459546
rect 424048 332648 424100 332654
rect 424048 332590 424100 332596
rect 423956 329520 424008 329526
rect 423956 329462 424008 329468
rect 423956 285320 424008 285326
rect 423956 285262 424008 285268
rect 423784 209746 423904 209774
rect 423876 201482 423904 209746
rect 423968 205018 423996 285262
rect 424060 206310 424088 332590
rect 425072 329730 425100 463014
rect 425164 458182 425192 583034
rect 425152 458176 425204 458182
rect 425152 458118 425204 458124
rect 425060 329724 425112 329730
rect 425060 329666 425112 329672
rect 424048 206304 424100 206310
rect 424048 206246 424100 206252
rect 423956 205012 424008 205018
rect 423956 204954 424008 204960
rect 424048 204604 424100 204610
rect 424048 204546 424100 204552
rect 423864 201476 423916 201482
rect 423864 201418 423916 201424
rect 423680 201340 423732 201346
rect 423680 201282 423732 201288
rect 423692 200114 423720 201282
rect 423692 200086 423812 200114
rect 422668 75676 422720 75682
rect 422668 75618 422720 75624
rect 423784 74458 423812 200086
rect 423876 75886 423904 201418
rect 423864 75880 423916 75886
rect 423864 75822 423916 75828
rect 423772 74452 423824 74458
rect 423772 74394 423824 74400
rect 424060 74322 424088 204546
rect 425072 201278 425100 329666
rect 425152 284980 425204 284986
rect 425152 284922 425204 284928
rect 425164 204950 425192 284922
rect 425244 205012 425296 205018
rect 425244 204954 425296 204960
rect 425152 204944 425204 204950
rect 425152 204886 425204 204892
rect 425060 201272 425112 201278
rect 425060 201214 425112 201220
rect 425072 200114 425100 201214
rect 425072 200086 425192 200114
rect 425164 74390 425192 200086
rect 425152 74384 425204 74390
rect 425152 74326 425204 74332
rect 424048 74316 424100 74322
rect 424048 74258 424100 74264
rect 425256 74254 425284 204954
rect 425244 74248 425296 74254
rect 425244 74190 425296 74196
rect 422300 57248 422352 57254
rect 422300 57190 422352 57196
rect 396460 54726 396842 54754
rect 399484 53100 399536 53106
rect 399484 53042 399536 53048
rect 396842 24682 397224 24698
rect 399496 24682 399524 53042
rect 396842 24676 397236 24682
rect 396842 24670 397184 24676
rect 397184 24618 397236 24624
rect 399484 24676 399536 24682
rect 399484 24618 399536 24624
rect 356992 24274 357374 24290
rect 356980 24268 357374 24274
rect 357032 24262 357374 24268
rect 356980 24210 357032 24216
rect 360660 24200 360712 24206
rect 390006 24168 390062 24177
rect 360712 24148 360962 24154
rect 360660 24142 360962 24148
rect 360672 24126 360962 24142
rect 371344 24138 371726 24154
rect 371332 24132 371726 24138
rect 371384 24126 371726 24132
rect 389666 24126 390006 24154
rect 390006 24103 390062 24112
rect 371332 24074 371384 24080
rect 266360 23520 266412 23526
rect 266360 23462 266412 23468
rect 267372 23520 267424 23526
rect 267424 23468 267674 23474
rect 267372 23462 267674 23468
rect 202892 23310 203090 23338
rect 205652 23310 206678 23338
rect 200028 22092 200080 22098
rect 200028 22034 200080 22040
rect 199476 21820 199528 21826
rect 199476 21762 199528 21768
rect 184848 21480 184900 21486
rect 184848 21422 184900 21428
rect 151820 21412 151872 21418
rect 151820 21354 151872 21360
rect 132500 20120 132552 20126
rect 132500 20062 132552 20068
rect 131120 17332 131172 17338
rect 131120 17274 131172 17280
rect 131132 16574 131160 17274
rect 132512 16574 132540 20062
rect 142804 20052 142856 20058
rect 142804 19994 142856 20000
rect 135260 18692 135312 18698
rect 135260 18634 135312 18640
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 125600 11892 125652 11898
rect 125600 11834 125652 11840
rect 96620 4820 96672 4826
rect 96620 4762 96672 4768
rect 66260 3460 66312 3466
rect 66260 3402 66312 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 11834
rect 128176 7676 128228 7682
rect 128176 7618 128228 7624
rect 128188 480 128216 7618
rect 129372 4888 129424 4894
rect 129372 4830 129424 4836
rect 129384 480 129412 4830
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 135272 3602 135300 18634
rect 135352 15972 135404 15978
rect 135352 15914 135404 15920
rect 135260 3596 135312 3602
rect 135260 3538 135312 3544
rect 135364 3482 135392 15914
rect 139584 13252 139636 13258
rect 139584 13194 139636 13200
rect 138848 4004 138900 4010
rect 138848 3946 138900 3952
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3538
rect 138860 480 138888 3946
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 13194
rect 142816 4010 142844 19994
rect 150624 11960 150676 11966
rect 150624 11902 150676 11908
rect 145472 11756 145524 11762
rect 145472 11698 145524 11704
rect 143540 6384 143592 6390
rect 143540 6326 143592 6332
rect 142804 4004 142856 4010
rect 142804 3946 142856 3952
rect 142436 3596 142488 3602
rect 142436 3538 142488 3544
rect 142448 480 142476 3538
rect 143552 480 143580 6326
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 11698
rect 147128 10532 147180 10538
rect 147128 10474 147180 10480
rect 147140 480 147168 10474
rect 149520 10396 149572 10402
rect 149520 10338 149572 10344
rect 149532 480 149560 10338
rect 150636 480 150664 11902
rect 151832 3534 151860 21354
rect 167000 19984 167052 19990
rect 167000 19926 167052 19932
rect 160100 18624 160152 18630
rect 160100 18566 160152 18572
rect 157800 7744 157852 7750
rect 157800 7686 157852 7692
rect 154212 4956 154264 4962
rect 154212 4898 154264 4904
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 153028 480 153056 3470
rect 154224 480 154252 4898
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 156616 480 156644 3470
rect 157812 480 157840 7686
rect 160112 480 160140 18566
rect 167012 16574 167040 19926
rect 175280 18760 175332 18766
rect 175280 18702 175332 18708
rect 171140 17400 171192 17406
rect 171140 17342 171192 17348
rect 171152 16574 171180 17342
rect 175292 16574 175320 18702
rect 184860 18630 184888 21422
rect 184848 18624 184900 18630
rect 184848 18566 184900 18572
rect 184940 18624 184992 18630
rect 184940 18566 184992 18572
rect 167012 16546 167224 16574
rect 171152 16546 172008 16574
rect 175292 16546 175504 16574
rect 164424 14612 164476 14618
rect 164424 14554 164476 14560
rect 161296 13184 161348 13190
rect 161296 13126 161348 13132
rect 161308 480 161336 13126
rect 163688 9036 163740 9042
rect 163688 8978 163740 8984
rect 163700 480 163728 8978
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14554
rect 167196 480 167224 16546
rect 168380 16040 168432 16046
rect 168380 15982 168432 15988
rect 168392 480 168420 15982
rect 170772 9104 170824 9110
rect 170772 9046 170824 9052
rect 170784 480 170812 9046
rect 171980 480 172008 16546
rect 173900 14476 173952 14482
rect 173900 14418 173952 14424
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 14418
rect 175476 480 175504 16546
rect 178592 14544 178644 14550
rect 178592 14486 178644 14492
rect 176660 13116 176712 13122
rect 176660 13058 176712 13064
rect 176672 3398 176700 13058
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177868 480 177896 3334
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 14486
rect 181444 6316 181496 6322
rect 181444 6258 181496 6264
rect 181456 480 181484 6258
rect 182548 5024 182600 5030
rect 182548 4966 182600 4972
rect 182560 480 182588 4966
rect 184952 480 184980 18566
rect 202892 11898 202920 23310
rect 202880 11892 202932 11898
rect 202880 11834 202932 11840
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 186148 480 186176 11766
rect 188528 10464 188580 10470
rect 188528 10406 188580 10412
rect 188540 480 188568 10406
rect 205652 4894 205680 23310
rect 210252 20126 210280 23324
rect 210240 20120 210292 20126
rect 210240 20062 210292 20068
rect 213840 18698 213868 23324
rect 216692 23310 217442 23338
rect 220832 23310 221030 23338
rect 223592 23310 224618 23338
rect 227732 23310 228206 23338
rect 230492 23310 231794 23338
rect 234632 23310 235382 23338
rect 238772 23310 238970 23338
rect 241532 23310 242558 23338
rect 245672 23310 246146 23338
rect 213828 18692 213880 18698
rect 213828 18634 213880 18640
rect 216692 13258 216720 23310
rect 216680 13252 216732 13258
rect 216680 13194 216732 13200
rect 217324 13252 217376 13258
rect 217324 13194 217376 13200
rect 205640 4888 205692 4894
rect 205640 4830 205692 4836
rect 217336 3602 217364 13194
rect 220832 6390 220860 23310
rect 223592 10538 223620 23310
rect 227732 11966 227760 23310
rect 227720 11960 227772 11966
rect 227720 11902 227772 11908
rect 223580 10532 223632 10538
rect 223580 10474 223632 10480
rect 220820 6384 220872 6390
rect 220820 6326 220872 6332
rect 230492 4962 230520 23310
rect 234632 7750 234660 23310
rect 238772 13190 238800 23310
rect 241532 14618 241560 23310
rect 242900 17264 242952 17270
rect 242900 17206 242952 17212
rect 241520 14612 241572 14618
rect 241520 14554 241572 14560
rect 238760 13184 238812 13190
rect 238760 13126 238812 13132
rect 241704 8968 241756 8974
rect 241704 8910 241756 8916
rect 234620 7744 234672 7750
rect 234620 7686 234672 7692
rect 230480 4956 230532 4962
rect 230480 4898 230532 4904
rect 217324 3596 217376 3602
rect 217324 3538 217376 3544
rect 239312 3460 239364 3466
rect 239312 3402 239364 3408
rect 239324 480 239352 3402
rect 241716 480 241744 8910
rect 242912 480 242940 17206
rect 245672 16046 245700 23310
rect 249720 17406 249748 23324
rect 253308 18766 253336 23324
rect 256712 23310 256910 23338
rect 259472 23310 260498 23338
rect 263612 23310 264086 23338
rect 253296 18760 253348 18766
rect 253296 18702 253348 18708
rect 249708 17400 249760 17406
rect 249708 17342 249760 17348
rect 245660 16040 245712 16046
rect 245660 15982 245712 15988
rect 245936 15904 245988 15910
rect 245936 15846 245988 15852
rect 245200 7608 245252 7614
rect 245200 7550 245252 7556
rect 245212 480 245240 7550
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 15846
rect 256712 14550 256740 23310
rect 256700 14544 256752 14550
rect 256700 14486 256752 14492
rect 248788 6248 248840 6254
rect 248788 6190 248840 6196
rect 248800 480 248828 6190
rect 249984 6180 250036 6186
rect 249984 6122 250036 6128
rect 249996 480 250024 6122
rect 259472 5030 259500 23310
rect 263612 11830 263640 23310
rect 263600 11824 263652 11830
rect 263600 11766 263652 11772
rect 259460 5024 259512 5030
rect 259460 4966 259512 4972
rect 252376 4820 252428 4826
rect 252376 4762 252428 4768
rect 252388 480 252416 4762
rect 266372 3466 266400 23462
rect 267384 23446 267674 23462
rect 270512 23310 271262 23338
rect 270512 7682 270540 23310
rect 274836 17338 274864 23324
rect 277412 23310 278438 23338
rect 274824 17332 274876 17338
rect 274824 17274 274876 17280
rect 277412 15978 277440 23310
rect 282012 20058 282040 23324
rect 284312 23310 285614 23338
rect 288452 23310 289202 23338
rect 292592 23310 292790 23338
rect 282000 20052 282052 20058
rect 282000 19994 282052 20000
rect 277400 15972 277452 15978
rect 277400 15914 277452 15920
rect 284312 13258 284340 23310
rect 284300 13252 284352 13258
rect 284300 13194 284352 13200
rect 288452 11762 288480 23310
rect 288440 11756 288492 11762
rect 288440 11698 288492 11704
rect 292592 10402 292620 23310
rect 296364 21418 296392 23324
rect 299492 23310 299966 23338
rect 296352 21412 296404 21418
rect 296352 21354 296404 21360
rect 292580 10396 292632 10402
rect 292580 10338 292632 10344
rect 270500 7676 270552 7682
rect 270500 7618 270552 7624
rect 299492 3534 299520 23310
rect 303540 21486 303568 23324
rect 306392 23310 307142 23338
rect 303528 21480 303580 21486
rect 303528 21422 303580 21428
rect 306392 9042 306420 23310
rect 310716 19990 310744 23324
rect 313292 23310 314318 23338
rect 317432 23310 317906 23338
rect 320192 23310 321494 23338
rect 324332 23310 325082 23338
rect 310704 19984 310756 19990
rect 310704 19926 310756 19932
rect 313292 9110 313320 23310
rect 317432 14482 317460 23310
rect 317420 14476 317472 14482
rect 317420 14418 317472 14424
rect 320192 13122 320220 23310
rect 320180 13116 320232 13122
rect 320180 13058 320232 13064
rect 313280 9104 313332 9110
rect 313280 9046 313332 9052
rect 306380 9036 306432 9042
rect 306380 8978 306432 8984
rect 324332 6322 324360 23310
rect 328656 18630 328684 23324
rect 331232 23310 332258 23338
rect 328644 18624 328696 18630
rect 328644 18566 328696 18572
rect 331232 10470 331260 23310
rect 335832 22234 335860 23324
rect 338132 23310 339434 23338
rect 335820 22228 335872 22234
rect 335820 22170 335872 22176
rect 331220 10464 331272 10470
rect 331220 10406 331272 10412
rect 338132 10334 338160 23310
rect 343008 21962 343036 23324
rect 346596 22166 346624 23324
rect 346584 22160 346636 22166
rect 346584 22102 346636 22108
rect 342996 21956 343048 21962
rect 342996 21898 343048 21904
rect 350184 21826 350212 23324
rect 353772 22302 353800 23324
rect 353760 22296 353812 22302
rect 353760 22238 353812 22244
rect 364536 22030 364564 23324
rect 364524 22024 364576 22030
rect 368124 22001 368152 23324
rect 364524 21966 364576 21972
rect 368110 21992 368166 22001
rect 368110 21927 368166 21936
rect 375300 21894 375328 23324
rect 378888 22098 378916 23324
rect 378876 22092 378928 22098
rect 378876 22034 378928 22040
rect 382476 22001 382504 23324
rect 386064 22098 386092 23324
rect 393240 22137 393268 23324
rect 393226 22128 393282 22137
rect 386052 22092 386104 22098
rect 527836 22098 527864 697546
rect 542372 459377 542400 702406
rect 580172 697604 580224 697610
rect 580172 697546 580224 697552
rect 580184 697241 580212 697546
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580276 459513 580304 683839
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580354 524512 580410 524521
rect 580354 524447 580410 524456
rect 580262 459504 580318 459513
rect 580262 459439 580318 459448
rect 542358 459368 542414 459377
rect 542358 459303 542414 459312
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 580276 53106 580304 378383
rect 580368 204241 580396 524447
rect 580460 332489 580488 630799
rect 580920 591025 580948 643991
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580538 365120 580594 365129
rect 580538 365055 580594 365064
rect 580446 332480 580502 332489
rect 580446 332415 580502 332424
rect 580354 204232 580410 204241
rect 580354 204167 580410 204176
rect 580552 75954 580580 365055
rect 580644 332353 580672 577623
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 485081 580948 537775
rect 580906 485072 580962 485081
rect 580906 485007 580962 485016
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 378457 580948 431559
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580630 332344 580686 332353
rect 580630 332279 580686 332288
rect 580540 75948 580592 75954
rect 580540 75890 580592 75896
rect 580264 53100 580316 53106
rect 580264 53042 580316 53048
rect 393226 22063 393282 22072
rect 527824 22092 527876 22098
rect 386052 22034 386104 22040
rect 527824 22034 527876 22040
rect 382462 21992 382518 22001
rect 382462 21927 382518 21936
rect 375288 21888 375340 21894
rect 375288 21830 375340 21836
rect 350172 21820 350224 21826
rect 350172 21762 350224 21768
rect 338120 10328 338172 10334
rect 338120 10270 338172 10276
rect 324320 6316 324372 6322
rect 324320 6258 324372 6264
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 266360 3460 266412 3466
rect 266360 3402 266412 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 658144 2834 658200
rect 3606 619112 3662 619168
rect 2778 607144 2834 607200
rect 3422 607144 3478 607200
rect 3422 606056 3478 606112
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 2778 410488 2834 410544
rect 3330 345344 3386 345400
rect 2778 293120 2834 293176
rect 2778 267144 2834 267200
rect 2778 241032 2834 241088
rect 2778 214920 2834 214976
rect 2778 149776 2834 149832
rect 3330 136720 3386 136776
rect 3054 71576 3110 71632
rect 3330 45464 3386 45520
rect 3514 566888 3570 566944
rect 3698 553832 3754 553888
rect 3698 502424 3754 502480
rect 3698 501744 3754 501800
rect 3698 449520 3754 449576
rect 3698 397432 3754 397488
rect 3606 319232 3662 319288
rect 3514 204040 3570 204096
rect 3514 188808 3570 188864
rect 3606 110608 3662 110664
rect 3514 32408 3570 32464
rect 3698 84632 3754 84688
rect 4802 75792 4858 75848
rect 4986 75656 5042 75712
rect 15014 460128 15070 460184
rect 16394 203496 16450 203552
rect 17406 458224 17462 458280
rect 18878 459448 18934 459504
rect 18878 458224 18934 458280
rect 20166 585792 20222 585848
rect 19154 457952 19210 458008
rect 17590 204176 17646 204232
rect 20350 459312 20406 459368
rect 20166 457408 20222 457464
rect 18970 204448 19026 204504
rect 18786 204312 18842 204368
rect 17866 204176 17922 204232
rect 17866 203904 17922 203960
rect 18878 202816 18934 202872
rect 19246 202816 19302 202872
rect 19154 74296 19210 74352
rect 24766 586336 24822 586392
rect 21454 585656 21510 585712
rect 52550 585792 52606 585848
rect 55218 585656 55274 585712
rect 47398 582936 47454 582992
rect 88338 541728 88394 541784
rect 117226 585792 117282 585848
rect 133050 585656 133106 585712
rect 136638 541592 136694 541648
rect 23202 458224 23258 458280
rect 21454 458088 21510 458144
rect 29366 459312 29422 459368
rect 21362 457408 21418 457464
rect 21362 332424 21418 332480
rect 21086 331336 21142 331392
rect 20626 331200 20682 331256
rect 20994 329740 20996 329760
rect 20996 329740 21048 329760
rect 21048 329740 21050 329760
rect 20994 329704 21050 329740
rect 21178 331200 21234 331256
rect 41418 460128 41474 460184
rect 39670 457952 39726 458008
rect 62854 459448 62910 459504
rect 55218 458088 55274 458144
rect 52550 457408 52606 457464
rect 104714 458088 104770 458144
rect 109866 457952 109922 458008
rect 122746 460808 122802 460864
rect 127898 460672 127954 460728
rect 135718 458924 135774 458960
rect 135718 458904 135720 458924
rect 135720 458904 135772 458924
rect 135772 458904 135774 458924
rect 136546 458904 136602 458960
rect 133050 458768 133106 458824
rect 119986 457816 120042 457872
rect 137926 458224 137982 458280
rect 138294 457952 138350 458008
rect 136546 413888 136602 413944
rect 24214 333920 24270 333976
rect 27526 332324 27528 332344
rect 27528 332324 27580 332344
rect 27580 332324 27582 332344
rect 27526 332288 27582 332324
rect 21454 332152 21510 332208
rect 31114 332424 31170 332480
rect 31114 332152 31170 332208
rect 55310 332424 55366 332480
rect 52550 332288 52606 332344
rect 21454 331336 21510 331392
rect 21362 331200 21418 331256
rect 96526 332580 96582 332616
rect 96526 332560 96528 332580
rect 96528 332560 96580 332580
rect 96580 332560 96582 332580
rect 99194 331744 99250 331800
rect 133050 331880 133106 331936
rect 21086 202816 21142 202872
rect 22006 204212 22008 204232
rect 22008 204212 22060 204232
rect 22060 204212 22062 204232
rect 22006 204176 22062 204212
rect 21362 202680 21418 202736
rect 24214 204040 24270 204096
rect 34518 204448 34574 204504
rect 37278 204312 37334 204368
rect 44822 203904 44878 203960
rect 62854 204176 62910 204232
rect 55310 202816 55366 202872
rect 52550 202680 52606 202736
rect 29366 202544 29422 202600
rect 23294 202272 23350 202328
rect 104714 202816 104770 202872
rect 119986 204312 120042 204368
rect 109866 202680 109922 202736
rect 135626 204176 135682 204232
rect 133786 204040 133842 204096
rect 130014 203496 130070 203552
rect 119986 202544 120042 202600
rect 138570 460808 138626 460864
rect 138478 458088 138534 458144
rect 138846 460672 138902 460728
rect 139674 585792 139730 585848
rect 139858 457816 139914 457872
rect 138662 329704 138718 329760
rect 138386 204176 138442 204232
rect 138570 204176 138626 204232
rect 138386 203496 138442 203552
rect 138294 202816 138350 202872
rect 24214 75792 24270 75848
rect 21638 75656 21694 75712
rect 21362 74432 21418 74488
rect 39946 74296 40002 74352
rect 42062 74160 42118 74216
rect 53010 74432 53066 74488
rect 53010 73888 53066 73944
rect 65522 75656 65578 75712
rect 86682 75112 86738 75168
rect 77298 65456 77354 65512
rect 99286 61648 99342 61704
rect 57058 61512 57114 61568
rect 99286 60560 99342 60616
rect 102874 60696 102930 60752
rect 102782 57976 102838 58032
rect 102598 56616 102654 56672
rect 57518 56344 57574 56400
rect 102138 55528 102194 55584
rect 102138 54304 102194 54360
rect 102230 53080 102286 53136
rect 102138 52556 102194 52592
rect 102138 52536 102140 52556
rect 102140 52536 102192 52556
rect 102192 52536 102194 52556
rect 57058 51720 57114 51776
rect 102138 50088 102194 50144
rect 103150 59608 103206 59664
rect 103058 58520 103114 58576
rect 131118 75112 131174 75168
rect 142066 460964 142122 461000
rect 142066 460944 142068 460964
rect 142068 460944 142120 460964
rect 142120 460944 142122 460964
rect 142250 457952 142306 458008
rect 141514 329704 141570 329760
rect 139858 204312 139914 204368
rect 139766 204040 139822 204096
rect 139398 202544 139454 202600
rect 139858 75112 139914 75168
rect 142342 332560 142398 332616
rect 142250 202680 142306 202736
rect 143538 60560 143594 60616
rect 144826 60560 144882 60616
rect 144826 59880 144882 59936
rect 103242 51040 103298 51096
rect 102874 48728 102930 48784
rect 102598 46960 102654 47016
rect 57518 46860 57520 46880
rect 57520 46860 57572 46880
rect 57572 46860 57574 46880
rect 57518 46824 57574 46860
rect 57150 42064 57206 42120
rect 57058 36896 57114 36952
rect 57610 31592 57666 31648
rect 57242 27104 57298 27160
rect 102322 43288 102378 43344
rect 102138 42880 102194 42936
rect 102230 41384 102286 41440
rect 102138 40024 102194 40080
rect 102966 47640 103022 47696
rect 195978 52264 196034 52320
rect 196070 51720 196126 51776
rect 195978 50904 196034 50960
rect 103426 45600 103482 45656
rect 103610 44376 103666 44432
rect 195978 49544 196034 49600
rect 196070 49136 196126 49192
rect 195978 47776 196034 47832
rect 195978 46860 195980 46880
rect 195980 46860 196032 46880
rect 196032 46860 196034 46880
rect 195978 46824 196034 46860
rect 196622 48184 196678 48240
rect 196162 46144 196218 46200
rect 195978 45192 196034 45248
rect 195978 44004 195980 44024
rect 195980 44004 196032 44024
rect 196032 44004 196034 44024
rect 195978 43968 196034 44004
rect 196070 43560 196126 43616
rect 195978 42472 196034 42528
rect 196070 42064 196126 42120
rect 195978 41112 196034 41168
rect 195978 39924 195980 39944
rect 195980 39924 196032 39944
rect 196032 39924 196034 39944
rect 195978 39888 196034 39924
rect 196070 39480 196126 39536
rect 102782 38936 102838 38992
rect 102598 37848 102654 37904
rect 102690 36080 102746 36136
rect 102138 34584 102194 34640
rect 196162 38528 196218 38584
rect 195978 37984 196034 38040
rect 102874 37304 102930 37360
rect 195978 37032 196034 37088
rect 195978 35844 195980 35864
rect 195980 35844 196032 35864
rect 196032 35844 196034 35864
rect 195978 35808 196034 35844
rect 196070 35400 196126 35456
rect 195978 34348 195980 34368
rect 195980 34348 196032 34368
rect 196032 34348 196034 34368
rect 195978 34312 196034 34348
rect 196070 33904 196126 33960
rect 102322 33496 102378 33552
rect 102138 32408 102194 32464
rect 102230 31728 102286 31784
rect 102138 30504 102194 30560
rect 195978 32952 196034 33008
rect 195978 31628 195980 31648
rect 195980 31628 196032 31648
rect 196032 31628 196034 31648
rect 195978 31592 196034 31628
rect 196070 31456 196126 31512
rect 195978 30096 196034 30152
rect 196070 29688 196126 29744
rect 102138 29280 102194 29336
rect 195978 28908 195980 28928
rect 195980 28908 196032 28928
rect 196032 28908 196034 28928
rect 195978 28872 196034 28908
rect 102138 28464 102194 28520
rect 195978 28056 196034 28112
rect 102138 27648 102194 27704
rect 195978 27240 196034 27296
rect 102782 26288 102838 26344
rect 195978 26188 195980 26208
rect 195980 26188 196032 26208
rect 196032 26188 196034 26208
rect 195978 26152 196034 26188
rect 3422 6432 3478 6488
rect 418158 699760 418214 699816
rect 218058 586336 218114 586392
rect 298006 585792 298062 585848
rect 229742 331880 229798 331936
rect 226246 57296 226302 57352
rect 241518 331744 241574 331800
rect 230846 59880 230902 59936
rect 295982 541592 296038 541648
rect 269762 458768 269818 458824
rect 297638 285504 297694 285560
rect 300306 459176 300362 459232
rect 298926 331744 298982 331800
rect 298926 331200 298982 331256
rect 300398 458224 300454 458280
rect 300490 456864 300546 456920
rect 299386 331200 299442 331256
rect 301318 585656 301374 585712
rect 301318 460944 301374 461000
rect 338026 585928 338082 585984
rect 335450 585656 335506 585712
rect 327722 582936 327778 582992
rect 358634 585792 358690 585848
rect 361210 580216 361266 580272
rect 384394 585656 384450 585712
rect 412730 585792 412786 585848
rect 418250 585656 418306 585712
rect 417882 585112 417938 585168
rect 300766 458088 300822 458144
rect 300766 456864 300822 456920
rect 299202 203496 299258 203552
rect 302698 459584 302754 459640
rect 304538 459448 304594 459504
rect 301962 459312 302018 459368
rect 307114 459176 307170 459232
rect 309690 458088 309746 458144
rect 338026 461080 338082 461136
rect 335450 460944 335506 461000
rect 301502 456748 301558 456784
rect 301502 456728 301504 456748
rect 301504 456728 301556 456748
rect 301556 456728 301558 456748
rect 389546 461080 389602 461136
rect 386970 460944 387026 461000
rect 407026 459584 407082 459640
rect 418158 459584 418214 459640
rect 412730 458224 412786 458280
rect 422298 585112 422354 585168
rect 418710 459584 418766 459640
rect 301962 332424 302018 332480
rect 303526 332288 303582 332344
rect 304538 332288 304594 332344
rect 306746 331744 306802 331800
rect 303526 331064 303582 331120
rect 379426 329704 379482 329760
rect 353298 285504 353354 285560
rect 417882 331200 417938 331256
rect 301134 204040 301190 204096
rect 304538 204312 304594 204368
rect 301962 204176 302018 204232
rect 335450 204040 335506 204096
rect 303526 203804 303528 203824
rect 303528 203804 303580 203824
rect 303580 203804 303582 203824
rect 303526 203768 303582 203804
rect 319350 203496 319406 203552
rect 303526 158652 303528 158672
rect 303528 158652 303580 158672
rect 303580 158652 303582 158672
rect 303526 158616 303582 158652
rect 411258 203496 411314 203552
rect 416778 204040 416834 204096
rect 302054 78512 302110 78568
rect 302330 60596 302332 60616
rect 302332 60596 302384 60616
rect 302384 60596 302386 60616
rect 302330 60560 302386 60596
rect 333978 76608 334034 76664
rect 346766 73752 346822 73808
rect 355046 73888 355102 73944
rect 371146 77832 371202 77888
rect 366362 74432 366418 74488
rect 373998 76744 374054 76800
rect 372618 76608 372674 76664
rect 374090 74296 374146 74352
rect 374642 74296 374698 74352
rect 386510 76472 386566 76528
rect 420826 331336 420882 331392
rect 421378 461080 421434 461136
rect 421286 460944 421342 461000
rect 419814 203496 419870 203552
rect 421102 204040 421158 204096
rect 418526 74432 418582 74488
rect 421378 74296 421434 74352
rect 422390 331200 422446 331256
rect 422666 460944 422722 461000
rect 422482 329704 422538 329760
rect 390006 24112 390062 24168
rect 368110 21936 368166 21992
rect 393226 22072 393282 22128
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 579986 471416 580042 471472
rect 580906 644000 580962 644056
rect 580446 630808 580502 630864
rect 580354 524456 580410 524512
rect 580262 459448 580318 459504
rect 542358 459312 542414 459368
rect 580262 378392 580318 378448
rect 580906 590960 580962 591016
rect 580630 577632 580686 577688
rect 580538 365064 580594 365120
rect 580446 332424 580502 332480
rect 580354 204176 580410 204232
rect 580906 537784 580962 537840
rect 580906 485016 580962 485072
rect 580906 431568 580962 431624
rect 580906 378392 580962 378448
rect 580630 332288 580686 332344
rect 382462 21936 382518 21992
<< metal3 >>
rect 418153 699820 418219 699821
rect 418102 699818 418108 699820
rect 418062 699758 418108 699818
rect 418172 699816 418219 699820
rect 418214 699760 418219 699816
rect 418102 699756 418108 699758
rect 418172 699756 418219 699760
rect 418153 699755 418219 699756
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect -960 671198 674 671258
rect -960 671122 480 671198
rect 614 671122 674 671198
rect -960 671108 674 671122
rect 246 671062 674 671108
rect 246 670714 306 671062
rect 17166 670714 17172 670716
rect 246 670654 17172 670714
rect 17166 670652 17172 670654
rect 17236 670652 17242 670716
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 583520 617388 584960 617628
rect 2773 607202 2839 607205
rect 3417 607202 3483 607205
rect 2773 607200 3483 607202
rect 2773 607144 2778 607200
rect 2834 607144 3422 607200
rect 3478 607144 3483 607200
rect 2773 607142 3483 607144
rect 2773 607139 2839 607142
rect 3417 607139 3483 607142
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 420126 591228 420132 591292
rect 420196 591290 420202 591292
rect 420196 591230 567210 591290
rect 420196 591228 420202 591230
rect 567150 591018 567210 591230
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 567150 591016 584960 591018
rect 567150 590960 580906 591016
rect 580962 590960 584960 591016
rect 567150 590958 584960 590960
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect 24761 586394 24827 586397
rect 218053 586394 218119 586397
rect 24761 586392 218119 586394
rect 24761 586336 24766 586392
rect 24822 586336 218058 586392
rect 218114 586336 218119 586392
rect 24761 586334 218119 586336
rect 24761 586331 24827 586334
rect 218053 586331 218119 586334
rect 303470 585924 303476 585988
rect 303540 585986 303546 585988
rect 338021 585986 338087 585989
rect 303540 585984 338087 585986
rect 303540 585928 338026 585984
rect 338082 585928 338087 585984
rect 303540 585926 338087 585928
rect 303540 585924 303546 585926
rect 338021 585923 338087 585926
rect 20161 585850 20227 585853
rect 52545 585850 52611 585853
rect 20161 585848 52611 585850
rect 20161 585792 20166 585848
rect 20222 585792 52550 585848
rect 52606 585792 52611 585848
rect 20161 585790 52611 585792
rect 20161 585787 20227 585790
rect 52545 585787 52611 585790
rect 117221 585850 117287 585853
rect 139669 585850 139735 585853
rect 117221 585848 139735 585850
rect 117221 585792 117226 585848
rect 117282 585792 139674 585848
rect 139730 585792 139735 585848
rect 117221 585790 139735 585792
rect 117221 585787 117287 585790
rect 139669 585787 139735 585790
rect 298001 585850 298067 585853
rect 358629 585850 358695 585853
rect 298001 585848 358695 585850
rect 298001 585792 298006 585848
rect 298062 585792 358634 585848
rect 358690 585792 358695 585848
rect 298001 585790 358695 585792
rect 298001 585787 298067 585790
rect 358629 585787 358695 585790
rect 412725 585850 412791 585853
rect 422334 585850 422340 585852
rect 412725 585848 422340 585850
rect 412725 585792 412730 585848
rect 412786 585792 422340 585848
rect 412725 585790 422340 585792
rect 412725 585787 412791 585790
rect 422334 585788 422340 585790
rect 422404 585788 422410 585852
rect 21449 585714 21515 585717
rect 55213 585714 55279 585717
rect 21449 585712 55279 585714
rect 21449 585656 21454 585712
rect 21510 585656 55218 585712
rect 55274 585656 55279 585712
rect 21449 585654 55279 585656
rect 21449 585651 21515 585654
rect 55213 585651 55279 585654
rect 133045 585714 133111 585717
rect 299974 585714 299980 585716
rect 133045 585712 299980 585714
rect 133045 585656 133050 585712
rect 133106 585656 299980 585712
rect 133045 585654 299980 585656
rect 133045 585651 133111 585654
rect 299974 585652 299980 585654
rect 300044 585652 300050 585716
rect 301313 585714 301379 585717
rect 335445 585714 335511 585717
rect 301313 585712 335511 585714
rect 301313 585656 301318 585712
rect 301374 585656 335450 585712
rect 335506 585656 335511 585712
rect 301313 585654 335511 585656
rect 301313 585651 301379 585654
rect 335445 585651 335511 585654
rect 384389 585714 384455 585717
rect 418245 585714 418311 585717
rect 384389 585712 418311 585714
rect 384389 585656 384394 585712
rect 384450 585656 418250 585712
rect 418306 585656 418311 585712
rect 384389 585654 418311 585656
rect 384389 585651 384455 585654
rect 418245 585651 418311 585654
rect 417877 585170 417943 585173
rect 422293 585170 422359 585173
rect 417877 585168 422359 585170
rect 417877 585112 417882 585168
rect 417938 585112 422298 585168
rect 422354 585112 422359 585168
rect 417877 585110 422359 585112
rect 417877 585107 417943 585110
rect 422293 585107 422359 585110
rect 23238 582932 23244 582996
rect 23308 582994 23314 582996
rect 47393 582994 47459 582997
rect 23308 582992 47459 582994
rect 23308 582936 47398 582992
rect 47454 582936 47459 582992
rect 23308 582934 47459 582936
rect 23308 582932 23314 582934
rect 47393 582931 47459 582934
rect 299238 582932 299244 582996
rect 299308 582994 299314 582996
rect 327717 582994 327783 582997
rect 299308 582992 327783 582994
rect 299308 582936 327722 582992
rect 327778 582936 327783 582992
rect 299308 582934 327783 582936
rect 299308 582932 299314 582934
rect 327717 582931 327783 582934
rect 301446 580212 301452 580276
rect 301516 580274 301522 580276
rect 361205 580274 361271 580277
rect 301516 580272 361271 580274
rect 301516 580216 361210 580272
rect 361266 580216 361271 580272
rect 301516 580214 361271 580216
rect 301516 580212 301522 580214
rect 361205 580211 361271 580214
rect -960 579852 480 580092
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect 88333 541786 88399 541789
rect 138054 541786 138060 541788
rect 88333 541784 138060 541786
rect 88333 541728 88338 541784
rect 88394 541728 138060 541784
rect 88333 541726 138060 541728
rect 88333 541723 88399 541726
rect 138054 541724 138060 541726
rect 138124 541724 138130 541788
rect 136633 541650 136699 541653
rect 295977 541650 296043 541653
rect 136633 541648 296043 541650
rect 136633 541592 136638 541648
rect 136694 541592 295982 541648
rect 296038 541592 296043 541648
rect 136633 541590 296043 541592
rect 136633 541587 136699 541590
rect 295977 541587 296043 541590
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 580349 524514 580415 524517
rect 583520 524514 584960 524604
rect 580349 524512 584960 524514
rect 580349 524456 580354 524512
rect 580410 524456 584960 524512
rect 580349 524454 584960 524456
rect 580349 524451 580415 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 583520 511172 584960 511412
rect 3693 502482 3759 502485
rect 19558 502482 19564 502484
rect 3693 502480 19564 502482
rect 3693 502424 3698 502480
rect 3754 502424 19564 502480
rect 3693 502422 19564 502424
rect 3693 502419 3759 502422
rect 19558 502420 19564 502422
rect 19628 502420 19634 502484
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 418654 485012 418660 485076
rect 418724 485074 418730 485076
rect 580901 485074 580967 485077
rect 418724 485072 583586 485074
rect 418724 485016 580906 485072
rect 580962 485016 583586 485072
rect 418724 485014 583586 485016
rect 418724 485012 418730 485014
rect 580901 485011 580967 485014
rect 583526 484802 583586 485014
rect 583342 484756 583586 484802
rect 583342 484742 584960 484756
rect 583342 484666 583402 484742
rect 583520 484666 584960 484742
rect 583342 484606 584960 484666
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 303470 461076 303476 461140
rect 303540 461138 303546 461140
rect 338021 461138 338087 461141
rect 303540 461136 338087 461138
rect 303540 461080 338026 461136
rect 338082 461080 338087 461136
rect 303540 461078 338087 461080
rect 303540 461076 303546 461078
rect 338021 461075 338087 461078
rect 389541 461138 389607 461141
rect 421373 461138 421439 461141
rect 389541 461136 422310 461138
rect 389541 461080 389546 461136
rect 389602 461080 421378 461136
rect 421434 461080 422310 461136
rect 389541 461078 422310 461080
rect 389541 461075 389607 461078
rect 421373 461075 421439 461078
rect 142061 461004 142127 461005
rect 142061 461002 142108 461004
rect 142016 461000 142108 461002
rect 142172 461002 142178 461004
rect 301313 461002 301379 461005
rect 335445 461002 335511 461005
rect 142016 460944 142066 461000
rect 142016 460942 142108 460944
rect 142061 460940 142108 460942
rect 142172 460942 142254 461002
rect 301313 461000 335511 461002
rect 301313 460944 301318 461000
rect 301374 460944 335450 461000
rect 335506 460944 335511 461000
rect 301313 460942 335511 460944
rect 142172 460940 142178 460942
rect 142061 460939 142127 460940
rect 301313 460939 301379 460942
rect 335445 460939 335511 460942
rect 386965 461002 387031 461005
rect 421281 461002 421347 461005
rect 386965 461000 421347 461002
rect 386965 460944 386970 461000
rect 387026 460944 421286 461000
rect 421342 460944 421347 461000
rect 386965 460942 421347 460944
rect 422250 461002 422310 461078
rect 422661 461002 422727 461005
rect 422250 461000 422727 461002
rect 422250 460944 422666 461000
rect 422722 460944 422727 461000
rect 422250 460942 422727 460944
rect 386965 460939 387031 460942
rect 421281 460939 421347 460942
rect 422661 460939 422727 460942
rect 122741 460866 122807 460869
rect 138565 460866 138631 460869
rect 122741 460864 138631 460866
rect 122741 460808 122746 460864
rect 122802 460808 138570 460864
rect 138626 460808 138631 460864
rect 122741 460806 138631 460808
rect 122741 460803 122807 460806
rect 138565 460803 138631 460806
rect 127893 460730 127959 460733
rect 138841 460730 138907 460733
rect 127893 460728 138907 460730
rect 127893 460672 127898 460728
rect 127954 460672 138846 460728
rect 138902 460672 138907 460728
rect 127893 460670 138907 460672
rect 127893 460667 127959 460670
rect 138841 460667 138907 460670
rect 15009 460186 15075 460189
rect 23238 460186 23244 460188
rect 15009 460184 23244 460186
rect 15009 460128 15014 460184
rect 15070 460128 23244 460184
rect 15009 460126 23244 460128
rect 15009 460123 15075 460126
rect 23238 460124 23244 460126
rect 23308 460186 23314 460188
rect 41413 460186 41479 460189
rect 23308 460184 41479 460186
rect 23308 460128 41418 460184
rect 41474 460128 41479 460184
rect 23308 460126 41479 460128
rect 23308 460124 23314 460126
rect 41413 460123 41479 460126
rect 302693 459644 302759 459645
rect 302693 459640 302740 459644
rect 302804 459642 302810 459644
rect 407021 459642 407087 459645
rect 418153 459642 418219 459645
rect 418705 459642 418771 459645
rect 302693 459584 302698 459640
rect 302693 459580 302740 459584
rect 302804 459582 302850 459642
rect 407021 459640 418771 459642
rect 407021 459584 407026 459640
rect 407082 459584 418158 459640
rect 418214 459584 418710 459640
rect 418766 459584 418771 459640
rect 407021 459582 418771 459584
rect 302804 459580 302810 459582
rect 302693 459579 302759 459580
rect 407021 459579 407087 459582
rect 418153 459579 418219 459582
rect 418705 459579 418771 459582
rect 18873 459506 18939 459509
rect 62849 459506 62915 459509
rect 18873 459504 62915 459506
rect 18873 459448 18878 459504
rect 18934 459448 62854 459504
rect 62910 459448 62915 459504
rect 18873 459446 62915 459448
rect 18873 459443 18939 459446
rect 62849 459443 62915 459446
rect 304533 459506 304599 459509
rect 580257 459506 580323 459509
rect 304533 459504 580323 459506
rect 304533 459448 304538 459504
rect 304594 459448 580262 459504
rect 580318 459448 580323 459504
rect 304533 459446 580323 459448
rect 304533 459443 304599 459446
rect 580257 459443 580323 459446
rect 20345 459370 20411 459373
rect 29361 459370 29427 459373
rect 20345 459368 29427 459370
rect 20345 459312 20350 459368
rect 20406 459312 29366 459368
rect 29422 459312 29427 459368
rect 20345 459310 29427 459312
rect 20345 459307 20411 459310
rect 29361 459307 29427 459310
rect 301957 459370 302023 459373
rect 542353 459370 542419 459373
rect 301957 459368 542419 459370
rect 301957 459312 301962 459368
rect 302018 459312 542358 459368
rect 542414 459312 542419 459368
rect 301957 459310 542419 459312
rect 301957 459307 302023 459310
rect 542353 459307 542419 459310
rect 300301 459234 300367 459237
rect 307109 459234 307175 459237
rect 300301 459232 307175 459234
rect 300301 459176 300306 459232
rect 300362 459176 307114 459232
rect 307170 459176 307175 459232
rect 300301 459174 307175 459176
rect 300301 459171 300367 459174
rect 307109 459171 307175 459174
rect 135713 458962 135779 458965
rect 136541 458962 136607 458965
rect 138054 458962 138060 458964
rect 135713 458960 138060 458962
rect 135713 458904 135718 458960
rect 135774 458904 136546 458960
rect 136602 458904 138060 458960
rect 135713 458902 138060 458904
rect 135713 458899 135779 458902
rect 136541 458899 136607 458902
rect 138054 458900 138060 458902
rect 138124 458900 138130 458964
rect 133045 458826 133111 458829
rect 269757 458826 269823 458829
rect 133045 458824 269823 458826
rect 133045 458768 133050 458824
rect 133106 458768 269762 458824
rect 269818 458768 269823 458824
rect 133045 458766 269823 458768
rect 133045 458763 133111 458766
rect 269757 458763 269823 458766
rect 17401 458282 17467 458285
rect 18873 458282 18939 458285
rect 17401 458280 18939 458282
rect 17401 458224 17406 458280
rect 17462 458224 18878 458280
rect 18934 458224 18939 458280
rect 17401 458222 18939 458224
rect 17401 458219 17467 458222
rect 18873 458219 18939 458222
rect 23197 458284 23263 458285
rect 23197 458280 23244 458284
rect 23308 458282 23314 458284
rect 137921 458282 137987 458285
rect 138606 458282 138612 458284
rect 23197 458224 23202 458280
rect 23197 458220 23244 458224
rect 23308 458222 23354 458282
rect 137921 458280 138612 458282
rect 137921 458224 137926 458280
rect 137982 458224 138612 458280
rect 137921 458222 138612 458224
rect 23308 458220 23314 458222
rect 23197 458219 23263 458220
rect 137921 458219 137987 458222
rect 138606 458220 138612 458222
rect 138676 458220 138682 458284
rect 299238 458220 299244 458284
rect 299308 458282 299314 458284
rect 300393 458282 300459 458285
rect 299308 458280 300459 458282
rect 299308 458224 300398 458280
rect 300454 458224 300459 458280
rect 299308 458222 300459 458224
rect 299308 458220 299314 458222
rect 300393 458219 300459 458222
rect 412725 458282 412791 458285
rect 421046 458282 421052 458284
rect 412725 458280 421052 458282
rect 412725 458224 412730 458280
rect 412786 458224 421052 458280
rect 412725 458222 421052 458224
rect 412725 458219 412791 458222
rect 421046 458220 421052 458222
rect 421116 458220 421122 458284
rect 21449 458146 21515 458149
rect 55213 458146 55279 458149
rect 21449 458144 55279 458146
rect 21449 458088 21454 458144
rect 21510 458088 55218 458144
rect 55274 458088 55279 458144
rect 21449 458086 55279 458088
rect 21449 458083 21515 458086
rect 55213 458083 55279 458086
rect 104709 458146 104775 458149
rect 138473 458146 138539 458149
rect 104709 458144 138539 458146
rect 104709 458088 104714 458144
rect 104770 458088 138478 458144
rect 138534 458088 138539 458144
rect 104709 458086 138539 458088
rect 104709 458083 104775 458086
rect 138473 458083 138539 458086
rect 300761 458146 300827 458149
rect 309685 458146 309751 458149
rect 300761 458144 309751 458146
rect 300761 458088 300766 458144
rect 300822 458088 309690 458144
rect 309746 458088 309751 458144
rect 300761 458086 309751 458088
rect 300761 458083 300827 458086
rect 309685 458083 309751 458086
rect 19149 458010 19215 458013
rect 39665 458010 39731 458013
rect 19149 458008 39731 458010
rect 19149 457952 19154 458008
rect 19210 457952 39670 458008
rect 39726 457952 39731 458008
rect 19149 457950 39731 457952
rect 19149 457947 19215 457950
rect 39665 457947 39731 457950
rect 109861 458010 109927 458013
rect 138289 458010 138355 458013
rect 142245 458010 142311 458013
rect 109861 458008 142311 458010
rect 109861 457952 109866 458008
rect 109922 457952 138294 458008
rect 138350 457952 142250 458008
rect 142306 457952 142311 458008
rect 583520 457996 584960 458236
rect 109861 457950 142311 457952
rect 109861 457947 109927 457950
rect 138289 457947 138355 457950
rect 142245 457947 142311 457950
rect 119981 457874 120047 457877
rect 139853 457874 139919 457877
rect 119981 457872 139919 457874
rect 119981 457816 119986 457872
rect 120042 457816 139858 457872
rect 139914 457816 139919 457872
rect 119981 457814 139919 457816
rect 119981 457811 120047 457814
rect 139853 457811 139919 457814
rect 20161 457466 20227 457469
rect 21357 457466 21423 457469
rect 52545 457466 52611 457469
rect 20161 457464 52611 457466
rect 20161 457408 20166 457464
rect 20222 457408 21362 457464
rect 21418 457408 52550 457464
rect 52606 457408 52611 457464
rect 20161 457406 52611 457408
rect 20161 457403 20227 457406
rect 21357 457403 21423 457406
rect 52545 457403 52611 457406
rect 300485 456922 300551 456925
rect 300761 456922 300827 456925
rect 300485 456920 300827 456922
rect 300485 456864 300490 456920
rect 300546 456864 300766 456920
rect 300822 456864 300827 456920
rect 300485 456862 300827 456864
rect 300485 456859 300551 456862
rect 300761 456859 300827 456862
rect 301497 456788 301563 456789
rect 301446 456786 301452 456788
rect 301406 456726 301452 456786
rect 301516 456784 301563 456788
rect 301558 456728 301563 456784
rect 301446 456724 301452 456726
rect 301516 456724 301563 456728
rect 301497 456723 301563 456724
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 301998 418236 302004 418300
rect 302068 418298 302074 418300
rect 583520 418298 584960 418388
rect 302068 418238 584960 418298
rect 302068 418236 302074 418238
rect 583520 418148 584960 418238
rect 136541 413946 136607 413949
rect 138054 413946 138060 413948
rect 136541 413944 138060 413946
rect 136541 413888 136546 413944
rect 136602 413888 138060 413944
rect 136541 413886 138060 413888
rect 136541 413883 136607 413886
rect 138054 413884 138060 413886
rect 138124 413884 138130 413948
rect -960 410546 480 410636
rect 2773 410546 2839 410549
rect -960 410544 2839 410546
rect -960 410488 2778 410544
rect 2834 410488 2839 410544
rect -960 410486 2839 410488
rect -960 410396 480 410486
rect 2773 410483 2839 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 3693 397490 3759 397493
rect -960 397488 3759 397490
rect -960 397432 3698 397488
rect 3754 397432 3759 397488
rect -960 397430 3759 397432
rect -960 397340 480 397430
rect 3693 397427 3759 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580257 378450 580323 378453
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 580906 378448
rect 580962 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 580533 365122 580599 365125
rect 583520 365122 584960 365212
rect 580533 365120 584960 365122
rect 580533 365064 580538 365120
rect 580594 365064 584960 365120
rect 580533 365062 584960 365064
rect 580533 365059 580599 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 674 358458
rect -960 358322 480 358398
rect 614 358322 674 358398
rect -960 358308 674 358322
rect 246 358262 674 358308
rect 246 357778 306 358262
rect 246 357718 6930 357778
rect 6870 357506 6930 357718
rect 19374 357506 19380 357508
rect 6870 357446 19380 357506
rect 19374 357444 19380 357446
rect 19444 357444 19450 357508
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect 17166 333916 17172 333980
rect 17236 333978 17242 333980
rect 24209 333978 24275 333981
rect 17236 333976 24275 333978
rect 17236 333920 24214 333976
rect 24270 333920 24275 333976
rect 17236 333918 24275 333920
rect 17236 333916 17242 333918
rect 24209 333915 24275 333918
rect 96521 332618 96587 332621
rect 142337 332618 142403 332621
rect 96521 332616 142403 332618
rect 96521 332560 96526 332616
rect 96582 332560 142342 332616
rect 142398 332560 142403 332616
rect 96521 332558 142403 332560
rect 96521 332555 96587 332558
rect 142337 332555 142403 332558
rect 21357 332482 21423 332485
rect 31109 332482 31175 332485
rect 55305 332482 55371 332485
rect 21357 332480 31034 332482
rect -960 332196 480 332436
rect 21357 332424 21362 332480
rect 21418 332424 31034 332480
rect 21357 332422 31034 332424
rect 21357 332419 21423 332422
rect 23238 332284 23244 332348
rect 23308 332346 23314 332348
rect 27521 332346 27587 332349
rect 23308 332344 27587 332346
rect 23308 332288 27526 332344
rect 27582 332288 27587 332344
rect 23308 332286 27587 332288
rect 30974 332346 31034 332422
rect 31109 332480 55371 332482
rect 31109 332424 31114 332480
rect 31170 332424 55310 332480
rect 55366 332424 55371 332480
rect 31109 332422 55371 332424
rect 31109 332419 31175 332422
rect 55305 332419 55371 332422
rect 301957 332482 302023 332485
rect 580441 332482 580507 332485
rect 301957 332480 580507 332482
rect 301957 332424 301962 332480
rect 302018 332424 580446 332480
rect 580502 332424 580507 332480
rect 301957 332422 580507 332424
rect 301957 332419 302023 332422
rect 580441 332419 580507 332422
rect 52545 332346 52611 332349
rect 30974 332344 52611 332346
rect 30974 332288 52550 332344
rect 52606 332288 52611 332344
rect 30974 332286 52611 332288
rect 23308 332284 23314 332286
rect 27521 332283 27587 332286
rect 52545 332283 52611 332286
rect 302918 332284 302924 332348
rect 302988 332346 302994 332348
rect 303521 332346 303587 332349
rect 302988 332344 303587 332346
rect 302988 332288 303526 332344
rect 303582 332288 303587 332344
rect 302988 332286 303587 332288
rect 302988 332284 302994 332286
rect 303521 332283 303587 332286
rect 304533 332346 304599 332349
rect 580625 332346 580691 332349
rect 304533 332344 580691 332346
rect 304533 332288 304538 332344
rect 304594 332288 580630 332344
rect 580686 332288 580691 332344
rect 304533 332286 580691 332288
rect 304533 332283 304599 332286
rect 580625 332283 580691 332286
rect 21449 332210 21515 332213
rect 31109 332210 31175 332213
rect 21449 332208 31175 332210
rect 21449 332152 21454 332208
rect 21510 332152 31114 332208
rect 31170 332152 31175 332208
rect 21449 332150 31175 332152
rect 21449 332147 21515 332150
rect 31109 332147 31175 332150
rect 133045 331938 133111 331941
rect 229737 331938 229803 331941
rect 133045 331936 229803 331938
rect 133045 331880 133050 331936
rect 133106 331880 229742 331936
rect 229798 331880 229803 331936
rect 133045 331878 229803 331880
rect 133045 331875 133111 331878
rect 229737 331875 229803 331878
rect 99189 331802 99255 331805
rect 241513 331802 241579 331805
rect 99189 331800 241579 331802
rect 99189 331744 99194 331800
rect 99250 331744 241518 331800
rect 241574 331744 241579 331800
rect 99189 331742 241579 331744
rect 99189 331739 99255 331742
rect 241513 331739 241579 331742
rect 298921 331802 298987 331805
rect 306741 331802 306807 331805
rect 298921 331800 306807 331802
rect 298921 331744 298926 331800
rect 298982 331744 306746 331800
rect 306802 331744 306807 331800
rect 298921 331742 306807 331744
rect 298921 331739 298987 331742
rect 306741 331739 306807 331742
rect 21081 331394 21147 331397
rect 21449 331394 21515 331397
rect 21081 331392 21515 331394
rect 21081 331336 21086 331392
rect 21142 331336 21454 331392
rect 21510 331336 21515 331392
rect 21081 331334 21515 331336
rect 21081 331331 21147 331334
rect 21449 331331 21515 331334
rect 419574 331332 419580 331396
rect 419644 331394 419650 331396
rect 420821 331394 420887 331397
rect 419644 331392 420887 331394
rect 419644 331336 420826 331392
rect 420882 331336 420887 331392
rect 419644 331334 420887 331336
rect 419644 331332 419650 331334
rect 420821 331331 420887 331334
rect 19374 331196 19380 331260
rect 19444 331258 19450 331260
rect 20621 331258 20687 331261
rect 19444 331256 20687 331258
rect 19444 331200 20626 331256
rect 20682 331200 20687 331256
rect 19444 331198 20687 331200
rect 19444 331196 19450 331198
rect 20621 331195 20687 331198
rect 21173 331258 21239 331261
rect 21357 331258 21423 331261
rect 21173 331256 21423 331258
rect 21173 331200 21178 331256
rect 21234 331200 21362 331256
rect 21418 331200 21423 331256
rect 21173 331198 21423 331200
rect 21173 331195 21239 331198
rect 21357 331195 21423 331198
rect 298921 331258 298987 331261
rect 299381 331258 299447 331261
rect 298921 331256 299447 331258
rect 298921 331200 298926 331256
rect 298982 331200 299386 331256
rect 299442 331200 299447 331256
rect 298921 331198 299447 331200
rect 298921 331195 298987 331198
rect 299381 331195 299447 331198
rect 417877 331258 417943 331261
rect 422385 331258 422451 331261
rect 417877 331256 422451 331258
rect 417877 331200 417882 331256
rect 417938 331200 422390 331256
rect 422446 331200 422451 331256
rect 417877 331198 422451 331200
rect 417877 331195 417943 331198
rect 422385 331195 422451 331198
rect 302734 331060 302740 331124
rect 302804 331122 302810 331124
rect 303521 331122 303587 331125
rect 302804 331120 303587 331122
rect 302804 331064 303526 331120
rect 303582 331064 303587 331120
rect 302804 331062 303587 331064
rect 302804 331060 302810 331062
rect 303521 331059 303587 331062
rect 20989 329762 21055 329765
rect 21214 329762 21220 329764
rect 20989 329760 21220 329762
rect 20989 329704 20994 329760
rect 21050 329704 21220 329760
rect 20989 329702 21220 329704
rect 20989 329699 21055 329702
rect 21214 329700 21220 329702
rect 21284 329700 21290 329764
rect 138054 329700 138060 329764
rect 138124 329762 138130 329764
rect 138657 329762 138723 329765
rect 138124 329760 138723 329762
rect 138124 329704 138662 329760
rect 138718 329704 138723 329760
rect 138124 329702 138723 329704
rect 138124 329700 138130 329702
rect 138657 329699 138723 329702
rect 141509 329762 141575 329765
rect 141918 329762 141924 329764
rect 141509 329760 141924 329762
rect 141509 329704 141514 329760
rect 141570 329704 141924 329760
rect 141509 329702 141924 329704
rect 141509 329699 141575 329702
rect 141918 329700 141924 329702
rect 141988 329700 141994 329764
rect 379421 329762 379487 329765
rect 422477 329762 422543 329765
rect 379421 329760 422543 329762
rect 379421 329704 379426 329760
rect 379482 329704 422482 329760
rect 422538 329704 422543 329760
rect 379421 329702 422543 329704
rect 379421 329699 379487 329702
rect 422477 329699 422543 329702
rect 583520 325124 584960 325364
rect -960 319290 480 319380
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 297633 285562 297699 285565
rect 353293 285562 353359 285565
rect 297633 285560 353359 285562
rect 297633 285504 297638 285560
rect 297694 285504 353298 285560
rect 353354 285504 353359 285560
rect 297633 285502 353359 285504
rect 297633 285499 297699 285502
rect 353293 285499 353359 285502
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 583520 205580 584960 205820
rect 18965 204506 19031 204509
rect 34513 204506 34579 204509
rect 18965 204504 34579 204506
rect 18965 204448 18970 204504
rect 19026 204448 34518 204504
rect 34574 204448 34579 204504
rect 18965 204446 34579 204448
rect 18965 204443 19031 204446
rect 34513 204443 34579 204446
rect 18781 204370 18847 204373
rect 37273 204370 37339 204373
rect 18781 204368 37339 204370
rect 18781 204312 18786 204368
rect 18842 204312 37278 204368
rect 37334 204312 37339 204368
rect 18781 204310 37339 204312
rect 18781 204307 18847 204310
rect 37273 204307 37339 204310
rect 119981 204370 120047 204373
rect 139853 204370 139919 204373
rect 119981 204368 139919 204370
rect 119981 204312 119986 204368
rect 120042 204312 139858 204368
rect 139914 204312 139919 204368
rect 119981 204310 139919 204312
rect 119981 204307 120047 204310
rect 139853 204307 139919 204310
rect 304533 204370 304599 204373
rect 419574 204370 419580 204372
rect 304533 204368 419580 204370
rect 304533 204312 304538 204368
rect 304594 204312 419580 204368
rect 304533 204310 419580 204312
rect 304533 204307 304599 204310
rect 419574 204308 419580 204310
rect 419644 204308 419650 204372
rect 17585 204234 17651 204237
rect 17861 204234 17927 204237
rect 17585 204232 17927 204234
rect 17585 204176 17590 204232
rect 17646 204176 17866 204232
rect 17922 204176 17927 204232
rect 17585 204174 17927 204176
rect 17585 204171 17651 204174
rect 17861 204171 17927 204174
rect 21214 204172 21220 204236
rect 21284 204234 21290 204236
rect 22001 204234 22067 204237
rect 62849 204234 62915 204237
rect 21284 204232 22067 204234
rect 21284 204176 22006 204232
rect 22062 204176 22067 204232
rect 21284 204174 22067 204176
rect 21284 204172 21290 204174
rect 22001 204171 22067 204174
rect 26190 204232 62915 204234
rect 26190 204176 62854 204232
rect 62910 204176 62915 204232
rect 26190 204174 62915 204176
rect 3509 204098 3575 204101
rect 24209 204098 24275 204101
rect 3509 204096 24275 204098
rect 3509 204040 3514 204096
rect 3570 204040 24214 204096
rect 24270 204040 24275 204096
rect 3509 204038 24275 204040
rect 3509 204035 3575 204038
rect 24209 204035 24275 204038
rect 17861 203962 17927 203965
rect 26190 203962 26250 204174
rect 62849 204171 62915 204174
rect 135621 204234 135687 204237
rect 138381 204234 138447 204237
rect 138565 204234 138631 204237
rect 135621 204232 138631 204234
rect 135621 204176 135626 204232
rect 135682 204176 138386 204232
rect 138442 204176 138570 204232
rect 138626 204176 138631 204232
rect 135621 204174 138631 204176
rect 135621 204171 135687 204174
rect 138381 204171 138447 204174
rect 138565 204171 138631 204174
rect 301957 204234 302023 204237
rect 580349 204234 580415 204237
rect 301957 204232 580415 204234
rect 301957 204176 301962 204232
rect 302018 204176 580354 204232
rect 580410 204176 580415 204232
rect 301957 204174 580415 204176
rect 301957 204171 302023 204174
rect 580349 204171 580415 204174
rect 133781 204098 133847 204101
rect 139761 204098 139827 204101
rect 133781 204096 139827 204098
rect 133781 204040 133786 204096
rect 133842 204040 139766 204096
rect 139822 204040 139827 204096
rect 133781 204038 139827 204040
rect 133781 204035 133847 204038
rect 139761 204035 139827 204038
rect 301129 204098 301195 204101
rect 335445 204098 335511 204101
rect 301129 204096 335511 204098
rect 301129 204040 301134 204096
rect 301190 204040 335450 204096
rect 335506 204040 335511 204096
rect 301129 204038 335511 204040
rect 301129 204035 301195 204038
rect 335445 204035 335511 204038
rect 416773 204098 416839 204101
rect 421097 204098 421163 204101
rect 416773 204096 421163 204098
rect 416773 204040 416778 204096
rect 416834 204040 421102 204096
rect 421158 204040 421163 204096
rect 416773 204038 421163 204040
rect 416773 204035 416839 204038
rect 421097 204035 421163 204038
rect 44817 203962 44883 203965
rect 17861 203960 26250 203962
rect 17861 203904 17866 203960
rect 17922 203904 26250 203960
rect 17861 203902 26250 203904
rect 35850 203960 44883 203962
rect 35850 203904 44822 203960
rect 44878 203904 44883 203960
rect 35850 203902 44883 203904
rect 17861 203899 17927 203902
rect 16389 203554 16455 203557
rect 23238 203554 23244 203556
rect 16389 203552 23244 203554
rect 16389 203496 16394 203552
rect 16450 203496 23244 203552
rect 16389 203494 23244 203496
rect 16389 203491 16455 203494
rect 23238 203492 23244 203494
rect 23308 203554 23314 203556
rect 35850 203554 35910 203902
rect 44817 203899 44883 203902
rect 302918 203764 302924 203828
rect 302988 203826 302994 203828
rect 303521 203826 303587 203829
rect 302988 203824 303587 203826
rect 302988 203768 303526 203824
rect 303582 203768 303587 203824
rect 302988 203766 303587 203768
rect 302988 203764 302994 203766
rect 303521 203763 303587 203766
rect 23308 203494 35910 203554
rect 130009 203554 130075 203557
rect 138381 203554 138447 203557
rect 130009 203552 138447 203554
rect 130009 203496 130014 203552
rect 130070 203496 138386 203552
rect 138442 203496 138447 203552
rect 130009 203494 138447 203496
rect 23308 203492 23314 203494
rect 130009 203491 130075 203494
rect 138381 203491 138447 203494
rect 299197 203554 299263 203557
rect 319345 203554 319411 203557
rect 299197 203552 319411 203554
rect 299197 203496 299202 203552
rect 299258 203496 319350 203552
rect 319406 203496 319411 203552
rect 299197 203494 319411 203496
rect 299197 203491 299263 203494
rect 319345 203491 319411 203494
rect 411253 203554 411319 203557
rect 419809 203554 419875 203557
rect 411253 203552 419875 203554
rect 411253 203496 411258 203552
rect 411314 203496 419814 203552
rect 419870 203496 419875 203552
rect 411253 203494 419875 203496
rect 411253 203491 411319 203494
rect 419809 203491 419875 203494
rect 18873 202874 18939 202877
rect 19241 202874 19307 202877
rect 21081 202874 21147 202877
rect 55305 202874 55371 202877
rect 18873 202872 20914 202874
rect 18873 202816 18878 202872
rect 18934 202816 19246 202872
rect 19302 202816 20914 202872
rect 18873 202814 20914 202816
rect 18873 202811 18939 202814
rect 19241 202811 19307 202814
rect 20854 202602 20914 202814
rect 21081 202872 55371 202874
rect 21081 202816 21086 202872
rect 21142 202816 55310 202872
rect 55366 202816 55371 202872
rect 21081 202814 55371 202816
rect 21081 202811 21147 202814
rect 55305 202811 55371 202814
rect 104709 202874 104775 202877
rect 138289 202874 138355 202877
rect 104709 202872 138355 202874
rect 104709 202816 104714 202872
rect 104770 202816 138294 202872
rect 138350 202816 138355 202872
rect 104709 202814 138355 202816
rect 104709 202811 104775 202814
rect 138289 202811 138355 202814
rect 21357 202738 21423 202741
rect 52545 202738 52611 202741
rect 21357 202736 52611 202738
rect 21357 202680 21362 202736
rect 21418 202680 52550 202736
rect 52606 202680 52611 202736
rect 21357 202678 52611 202680
rect 21357 202675 21423 202678
rect 52545 202675 52611 202678
rect 109861 202738 109927 202741
rect 142245 202738 142311 202741
rect 109861 202736 142311 202738
rect 109861 202680 109866 202736
rect 109922 202680 142250 202736
rect 142306 202680 142311 202736
rect 109861 202678 142311 202680
rect 109861 202675 109927 202678
rect 142245 202675 142311 202678
rect 29361 202602 29427 202605
rect 20854 202600 29427 202602
rect 20854 202544 29366 202600
rect 29422 202544 29427 202600
rect 20854 202542 29427 202544
rect 29361 202539 29427 202542
rect 119981 202602 120047 202605
rect 139393 202602 139459 202605
rect 119981 202600 139459 202602
rect 119981 202544 119986 202600
rect 120042 202544 139398 202600
rect 139454 202544 139459 202600
rect 119981 202542 139459 202544
rect 119981 202539 120047 202542
rect 139393 202539 139459 202542
rect 23289 202332 23355 202333
rect 23238 202330 23244 202332
rect 23198 202270 23244 202330
rect 23308 202328 23355 202332
rect 23350 202272 23355 202328
rect 23238 202268 23244 202270
rect 23308 202268 23355 202272
rect 23289 202267 23355 202268
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 302734 158612 302740 158676
rect 302804 158674 302810 158676
rect 303521 158674 303587 158677
rect 302804 158672 303587 158674
rect 302804 158616 303526 158672
rect 303582 158616 303587 158672
rect 302804 158614 303587 158616
rect 302804 158612 302810 158614
rect 303521 158611 303587 158614
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110666 480 110756
rect 3601 110666 3667 110669
rect -960 110664 3667 110666
rect -960 110608 3606 110664
rect 3662 110608 3667 110664
rect -960 110606 3667 110608
rect -960 110516 480 110606
rect 3601 110603 3667 110606
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 302049 78572 302115 78573
rect 301998 78508 302004 78572
rect 302068 78570 302115 78572
rect 302068 78568 302160 78570
rect 302110 78512 302160 78568
rect 302068 78510 302160 78512
rect 302068 78508 302115 78510
rect 302049 78507 302115 78508
rect 299974 77828 299980 77892
rect 300044 77890 300050 77892
rect 371141 77890 371207 77893
rect 300044 77888 371207 77890
rect 300044 77832 371146 77888
rect 371202 77832 371207 77888
rect 300044 77830 371207 77832
rect 300044 77828 300050 77830
rect 371141 77827 371207 77830
rect 373993 76802 374059 76805
rect 421046 76802 421052 76804
rect 373993 76800 421052 76802
rect 373993 76744 373998 76800
rect 374054 76744 421052 76800
rect 373993 76742 421052 76744
rect 373993 76739 374059 76742
rect 421046 76740 421052 76742
rect 421116 76740 421122 76804
rect 303102 76604 303108 76668
rect 303172 76666 303178 76668
rect 333973 76666 334039 76669
rect 303172 76664 334039 76666
rect 303172 76608 333978 76664
rect 334034 76608 334039 76664
rect 303172 76606 334039 76608
rect 303172 76604 303178 76606
rect 333973 76603 334039 76606
rect 372613 76666 372679 76669
rect 422334 76666 422340 76668
rect 372613 76664 422340 76666
rect 372613 76608 372618 76664
rect 372674 76608 422340 76664
rect 372613 76606 422340 76608
rect 372613 76603 372679 76606
rect 422334 76604 422340 76606
rect 422404 76604 422410 76668
rect 138606 76468 138612 76532
rect 138676 76530 138682 76532
rect 386505 76530 386571 76533
rect 138676 76528 386571 76530
rect 138676 76472 386510 76528
rect 386566 76472 386571 76528
rect 138676 76470 386571 76472
rect 138676 76468 138682 76470
rect 386505 76467 386571 76470
rect 4797 75850 4863 75853
rect 24209 75850 24275 75853
rect 4797 75848 24275 75850
rect 4797 75792 4802 75848
rect 4858 75792 24214 75848
rect 24270 75792 24275 75848
rect 4797 75790 24275 75792
rect 4797 75787 4863 75790
rect 24209 75787 24275 75790
rect 4981 75714 5047 75717
rect 21633 75714 21699 75717
rect 4981 75712 21699 75714
rect 4981 75656 4986 75712
rect 5042 75656 21638 75712
rect 21694 75656 21699 75712
rect 4981 75654 21699 75656
rect 4981 75651 5047 75654
rect 21633 75651 21699 75654
rect 21950 75652 21956 75716
rect 22020 75714 22026 75716
rect 65517 75714 65583 75717
rect 22020 75712 65583 75714
rect 22020 75656 65522 75712
rect 65578 75656 65583 75712
rect 22020 75654 65583 75656
rect 22020 75652 22026 75654
rect 65517 75651 65583 75654
rect 86677 75170 86743 75173
rect 98494 75170 98500 75172
rect 86677 75168 98500 75170
rect 86677 75112 86682 75168
rect 86738 75112 98500 75168
rect 86677 75110 98500 75112
rect 86677 75107 86743 75110
rect 98494 75108 98500 75110
rect 98564 75108 98570 75172
rect 131113 75170 131179 75173
rect 139853 75170 139919 75173
rect 131113 75168 139919 75170
rect 131113 75112 131118 75168
rect 131174 75112 139858 75168
rect 139914 75112 139919 75168
rect 131113 75110 139919 75112
rect 131113 75107 131179 75110
rect 139853 75107 139919 75110
rect 21357 74490 21423 74493
rect 53005 74490 53071 74493
rect 21357 74488 53071 74490
rect 21357 74432 21362 74488
rect 21418 74432 53010 74488
rect 53066 74432 53071 74488
rect 21357 74430 53071 74432
rect 21357 74427 21423 74430
rect 53005 74427 53071 74430
rect 366357 74490 366423 74493
rect 418521 74490 418587 74493
rect 366357 74488 418587 74490
rect 366357 74432 366362 74488
rect 366418 74432 418526 74488
rect 418582 74432 418587 74488
rect 366357 74430 418587 74432
rect 366357 74427 366423 74430
rect 418521 74427 418587 74430
rect 19149 74354 19215 74357
rect 39941 74354 40007 74357
rect 374085 74354 374151 74357
rect 374637 74354 374703 74357
rect 421373 74354 421439 74357
rect 19149 74352 45570 74354
rect 19149 74296 19154 74352
rect 19210 74296 39946 74352
rect 40002 74296 45570 74352
rect 19149 74294 45570 74296
rect 19149 74291 19215 74294
rect 39941 74291 40007 74294
rect 23238 74156 23244 74220
rect 23308 74218 23314 74220
rect 42057 74218 42123 74221
rect 23308 74216 42123 74218
rect 23308 74160 42062 74216
rect 42118 74160 42123 74216
rect 23308 74158 42123 74160
rect 23308 74156 23314 74158
rect 42057 74155 42123 74158
rect 45510 73810 45570 74294
rect 374085 74352 421439 74354
rect 374085 74296 374090 74352
rect 374146 74296 374642 74352
rect 374698 74296 421378 74352
rect 421434 74296 421439 74352
rect 374085 74294 421439 74296
rect 374085 74291 374151 74294
rect 374637 74291 374703 74294
rect 421373 74291 421439 74294
rect 53005 73946 53071 73949
rect 355041 73946 355107 73949
rect 53005 73944 355107 73946
rect 53005 73888 53010 73944
rect 53066 73888 355046 73944
rect 355102 73888 355107 73944
rect 53005 73886 355107 73888
rect 53005 73883 53071 73886
rect 355041 73883 355107 73886
rect 346761 73810 346827 73813
rect 45510 73808 346827 73810
rect 45510 73752 346766 73808
rect 346822 73752 346827 73808
rect 45510 73750 346827 73752
rect 346761 73747 346827 73750
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 3049 71634 3115 71637
rect -960 71632 3115 71634
rect -960 71576 3054 71632
rect 3110 71576 3115 71632
rect -960 71574 3115 71576
rect -960 71484 480 71574
rect 3049 71571 3115 71574
rect 77293 65514 77359 65517
rect 98678 65514 98684 65516
rect 77293 65512 98684 65514
rect 77293 65456 77298 65512
rect 77354 65456 98684 65512
rect 77293 65454 98684 65456
rect 77293 65451 77359 65454
rect 98678 65452 98684 65454
rect 98748 65452 98754 65516
rect 98494 61644 98500 61708
rect 98564 61706 98570 61708
rect 99281 61706 99347 61709
rect 98564 61704 99347 61706
rect 98564 61648 99286 61704
rect 99342 61648 99347 61704
rect 98564 61646 99347 61648
rect 98564 61644 98570 61646
rect 99281 61643 99347 61646
rect 57053 61570 57119 61573
rect 57053 61568 60106 61570
rect 57053 61512 57058 61568
rect 57114 61512 60106 61568
rect 57053 61510 60106 61512
rect 57053 61507 57119 61510
rect 60046 61064 60106 61510
rect 99790 60754 99850 61336
rect 102869 60754 102935 60757
rect 99790 60752 102935 60754
rect 99790 60696 102874 60752
rect 102930 60696 102935 60752
rect 99790 60694 102935 60696
rect 102869 60691 102935 60694
rect 99281 60618 99347 60621
rect 143533 60618 143599 60621
rect 144821 60618 144887 60621
rect 99281 60616 144887 60618
rect 99281 60560 99286 60616
rect 99342 60560 143538 60616
rect 143594 60560 144826 60616
rect 144882 60560 144887 60616
rect 99281 60558 144887 60560
rect 99281 60555 99347 60558
rect 143533 60555 143599 60558
rect 144821 60555 144887 60558
rect 302325 60618 302391 60621
rect 302734 60618 302740 60620
rect 302325 60616 302740 60618
rect 302325 60560 302330 60616
rect 302386 60560 302740 60616
rect 302325 60558 302740 60560
rect 302325 60555 302391 60558
rect 302734 60556 302740 60558
rect 302804 60556 302810 60620
rect 99790 59666 99850 60248
rect 144821 59938 144887 59941
rect 230841 59938 230907 59941
rect 144821 59936 230907 59938
rect 144821 59880 144826 59936
rect 144882 59880 230846 59936
rect 230902 59880 230907 59936
rect 144821 59878 230907 59880
rect 144821 59875 144887 59878
rect 230841 59875 230907 59878
rect 103145 59666 103211 59669
rect 99790 59664 103211 59666
rect 99790 59608 103150 59664
rect 103206 59608 103211 59664
rect 99790 59606 103211 59608
rect 103145 59603 103211 59606
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 99790 58578 99850 59160
rect 103053 58578 103119 58581
rect 99790 58576 103119 58578
rect 99790 58520 103058 58576
rect 103114 58520 103119 58576
rect 99790 58518 103119 58520
rect 103053 58515 103119 58518
rect 99790 58034 99850 58072
rect 102777 58034 102843 58037
rect 99790 58032 102843 58034
rect 99790 57976 102782 58032
rect 102838 57976 102843 58032
rect 99790 57974 102843 57976
rect 102777 57971 102843 57974
rect 99414 57292 99420 57356
rect 99484 57354 99490 57356
rect 226241 57354 226307 57357
rect 99484 57352 226307 57354
rect 99484 57296 226246 57352
rect 226302 57296 226307 57352
rect 99484 57294 226307 57296
rect 99484 57292 99490 57294
rect 226241 57291 226307 57294
rect 99790 56674 99850 56984
rect 102593 56674 102659 56677
rect 99790 56672 102659 56674
rect 99790 56616 102598 56672
rect 102654 56616 102659 56672
rect 99790 56614 102659 56616
rect 102593 56611 102659 56614
rect 57513 56402 57579 56405
rect 57513 56400 60106 56402
rect 57513 56344 57518 56400
rect 57574 56344 60106 56400
rect 57513 56342 60106 56344
rect 57513 56339 57579 56342
rect 60046 56168 60106 56342
rect 99790 55586 99850 55896
rect 102133 55586 102199 55589
rect 99790 55584 102199 55586
rect 99790 55528 102138 55584
rect 102194 55528 102199 55584
rect 99790 55526 102199 55528
rect 102133 55523 102199 55526
rect 99790 54362 99850 54808
rect 102133 54362 102199 54365
rect 99790 54360 102199 54362
rect 99790 54304 102138 54360
rect 102194 54304 102199 54360
rect 99790 54302 102199 54304
rect 102133 54299 102199 54302
rect 99790 53138 99850 53720
rect 102225 53138 102291 53141
rect 99790 53136 102291 53138
rect 99790 53080 102230 53136
rect 102286 53080 102291 53136
rect 99790 53078 102291 53080
rect 102225 53075 102291 53078
rect 99790 52594 99850 52632
rect 102133 52594 102199 52597
rect 99790 52592 102199 52594
rect 99790 52536 102138 52592
rect 102194 52536 102199 52592
rect 99790 52534 102199 52536
rect 102133 52531 102199 52534
rect 195973 52322 196039 52325
rect 195973 52320 199394 52322
rect 195973 52264 195978 52320
rect 196034 52264 199394 52320
rect 195973 52262 199394 52264
rect 195973 52259 196039 52262
rect 199334 52088 199394 52262
rect 57053 51778 57119 51781
rect 196065 51778 196131 51781
rect 57053 51776 60106 51778
rect 57053 51720 57058 51776
rect 57114 51720 60106 51776
rect 57053 51718 60106 51720
rect 57053 51715 57119 51718
rect 60046 51272 60106 51718
rect 196065 51776 199394 51778
rect 196065 51720 196070 51776
rect 196126 51720 199394 51776
rect 196065 51718 199394 51720
rect 196065 51715 196131 51718
rect 99790 51098 99850 51544
rect 199334 51272 199394 51718
rect 103237 51098 103303 51101
rect 99790 51096 103303 51098
rect 99790 51040 103242 51096
rect 103298 51040 103303 51096
rect 99790 51038 103303 51040
rect 103237 51035 103303 51038
rect 195973 50962 196039 50965
rect 195973 50960 199394 50962
rect 195973 50904 195978 50960
rect 196034 50904 199394 50960
rect 195973 50902 199394 50904
rect 195973 50899 196039 50902
rect 199334 50456 199394 50902
rect 99790 50146 99850 50456
rect 102133 50146 102199 50149
rect 99790 50144 102199 50146
rect 99790 50088 102138 50144
rect 102194 50088 102199 50144
rect 99790 50086 102199 50088
rect 102133 50083 102199 50086
rect 195973 49602 196039 49605
rect 199334 49602 199394 49640
rect 195973 49600 199394 49602
rect 195973 49544 195978 49600
rect 196034 49544 199394 49600
rect 195973 49542 199394 49544
rect 195973 49539 196039 49542
rect 99790 48786 99850 49368
rect 196065 49194 196131 49197
rect 196065 49192 199394 49194
rect 196065 49136 196070 49192
rect 196126 49136 199394 49192
rect 196065 49134 199394 49136
rect 196065 49131 196131 49134
rect 199334 48824 199394 49134
rect 102869 48786 102935 48789
rect 99790 48784 102935 48786
rect 99790 48728 102874 48784
rect 102930 48728 102935 48784
rect 99790 48726 102935 48728
rect 102869 48723 102935 48726
rect 99790 47698 99850 48280
rect 196617 48242 196683 48245
rect 196617 48240 199394 48242
rect 196617 48184 196622 48240
rect 196678 48184 199394 48240
rect 196617 48182 199394 48184
rect 196617 48179 196683 48182
rect 199334 48008 199394 48182
rect 195973 47834 196039 47837
rect 195973 47832 199394 47834
rect 195973 47776 195978 47832
rect 196034 47776 199394 47832
rect 195973 47774 199394 47776
rect 195973 47771 196039 47774
rect 102961 47698 103027 47701
rect 99790 47696 103027 47698
rect 99790 47640 102966 47696
rect 103022 47640 103027 47696
rect 99790 47638 103027 47640
rect 102961 47635 103027 47638
rect 199334 47192 199394 47774
rect 99790 47018 99850 47192
rect 102593 47018 102659 47021
rect 99790 47016 102659 47018
rect 99790 46960 102598 47016
rect 102654 46960 102659 47016
rect 99790 46958 102659 46960
rect 102593 46955 102659 46958
rect 57513 46882 57579 46885
rect 195973 46882 196039 46885
rect 57513 46880 60106 46882
rect 57513 46824 57518 46880
rect 57574 46824 60106 46880
rect 57513 46822 60106 46824
rect 57513 46819 57579 46822
rect 60046 46376 60106 46822
rect 195973 46880 199394 46882
rect 195973 46824 195978 46880
rect 196034 46824 199394 46880
rect 195973 46822 199394 46824
rect 195973 46819 196039 46822
rect 199334 46376 199394 46822
rect 196157 46202 196223 46205
rect 196157 46200 199394 46202
rect 196157 46144 196162 46200
rect 196218 46144 199394 46200
rect 583520 46188 584960 46428
rect 196157 46142 199394 46144
rect 196157 46139 196223 46142
rect 99790 45658 99850 46104
rect 103421 45658 103487 45661
rect 99790 45656 103487 45658
rect -960 45522 480 45612
rect 99790 45600 103426 45656
rect 103482 45600 103487 45656
rect 99790 45598 103487 45600
rect 103421 45595 103487 45598
rect 199334 45560 199394 46142
rect 3325 45522 3391 45525
rect -960 45520 3391 45522
rect -960 45464 3330 45520
rect 3386 45464 3391 45520
rect -960 45462 3391 45464
rect -960 45372 480 45462
rect 3325 45459 3391 45462
rect 195973 45250 196039 45253
rect 195973 45248 199394 45250
rect 195973 45192 195978 45248
rect 196034 45192 199394 45248
rect 195973 45190 199394 45192
rect 195973 45187 196039 45190
rect 99790 44434 99850 45016
rect 199334 44744 199394 45190
rect 103605 44434 103671 44437
rect 99790 44432 103671 44434
rect 99790 44376 103610 44432
rect 103666 44376 103671 44432
rect 99790 44374 103671 44376
rect 103605 44371 103671 44374
rect 195973 44026 196039 44029
rect 195973 44024 199394 44026
rect 195973 43968 195978 44024
rect 196034 43968 199394 44024
rect 195973 43966 199394 43968
rect 195973 43963 196039 43966
rect 199334 43928 199394 43966
rect 99790 43346 99850 43928
rect 196065 43618 196131 43621
rect 196065 43616 199394 43618
rect 196065 43560 196070 43616
rect 196126 43560 199394 43616
rect 196065 43558 199394 43560
rect 196065 43555 196131 43558
rect 102317 43346 102383 43349
rect 99790 43344 102383 43346
rect 99790 43288 102322 43344
rect 102378 43288 102383 43344
rect 99790 43286 102383 43288
rect 102317 43283 102383 43286
rect 199334 43112 199394 43558
rect 102133 42938 102199 42941
rect 99790 42936 102199 42938
rect 99790 42880 102138 42936
rect 102194 42880 102199 42936
rect 99790 42878 102199 42880
rect 99790 42840 99850 42878
rect 102133 42875 102199 42878
rect 195973 42530 196039 42533
rect 195973 42528 199394 42530
rect 195973 42472 195978 42528
rect 196034 42472 199394 42528
rect 195973 42470 199394 42472
rect 195973 42467 196039 42470
rect 199334 42296 199394 42470
rect 57145 42122 57211 42125
rect 196065 42122 196131 42125
rect 57145 42120 60106 42122
rect 57145 42064 57150 42120
rect 57206 42064 60106 42120
rect 57145 42062 60106 42064
rect 57145 42059 57211 42062
rect 60046 41480 60106 42062
rect 196065 42120 199394 42122
rect 196065 42064 196070 42120
rect 196126 42064 199394 42120
rect 196065 42062 199394 42064
rect 196065 42059 196131 42062
rect 99790 41442 99850 41752
rect 199334 41480 199394 42062
rect 102225 41442 102291 41445
rect 99790 41440 102291 41442
rect 99790 41384 102230 41440
rect 102286 41384 102291 41440
rect 99790 41382 102291 41384
rect 102225 41379 102291 41382
rect 195973 41170 196039 41173
rect 195973 41168 199394 41170
rect 195973 41112 195978 41168
rect 196034 41112 199394 41168
rect 195973 41110 199394 41112
rect 195973 41107 196039 41110
rect 199334 40664 199394 41110
rect 99790 40082 99850 40664
rect 102133 40082 102199 40085
rect 99790 40080 102199 40082
rect 99790 40024 102138 40080
rect 102194 40024 102199 40080
rect 99790 40022 102199 40024
rect 102133 40019 102199 40022
rect 195973 39946 196039 39949
rect 195973 39944 199394 39946
rect 195973 39888 195978 39944
rect 196034 39888 199394 39944
rect 195973 39886 199394 39888
rect 195973 39883 196039 39886
rect 199334 39848 199394 39886
rect 99790 38994 99850 39576
rect 196065 39538 196131 39541
rect 196065 39536 199394 39538
rect 196065 39480 196070 39536
rect 196126 39480 199394 39536
rect 196065 39478 199394 39480
rect 196065 39475 196131 39478
rect 199334 39032 199394 39478
rect 102777 38994 102843 38997
rect 99790 38992 102843 38994
rect 99790 38936 102782 38992
rect 102838 38936 102843 38992
rect 99790 38934 102843 38936
rect 102777 38931 102843 38934
rect 196157 38586 196223 38589
rect 196157 38584 199394 38586
rect 196157 38528 196162 38584
rect 196218 38528 199394 38584
rect 196157 38526 199394 38528
rect 196157 38523 196223 38526
rect 99790 37906 99850 38488
rect 199334 38216 199394 38526
rect 195973 38042 196039 38045
rect 195973 38040 199394 38042
rect 195973 37984 195978 38040
rect 196034 37984 199394 38040
rect 195973 37982 199394 37984
rect 195973 37979 196039 37982
rect 102593 37906 102659 37909
rect 99790 37904 102659 37906
rect 99790 37848 102598 37904
rect 102654 37848 102659 37904
rect 99790 37846 102659 37848
rect 102593 37843 102659 37846
rect 199334 37400 199394 37982
rect 99790 37362 99850 37400
rect 102869 37362 102935 37365
rect 99790 37360 102935 37362
rect 99790 37304 102874 37360
rect 102930 37304 102935 37360
rect 99790 37302 102935 37304
rect 102869 37299 102935 37302
rect 195973 37090 196039 37093
rect 195973 37088 199394 37090
rect 195973 37032 195978 37088
rect 196034 37032 199394 37088
rect 195973 37030 199394 37032
rect 195973 37027 196039 37030
rect 57053 36954 57119 36957
rect 57053 36952 60106 36954
rect 57053 36896 57058 36952
rect 57114 36896 60106 36952
rect 57053 36894 60106 36896
rect 57053 36891 57119 36894
rect 60046 36584 60106 36894
rect 199334 36584 199394 37030
rect 99790 36138 99850 36312
rect 102685 36138 102751 36141
rect 99790 36136 102751 36138
rect 99790 36080 102690 36136
rect 102746 36080 102751 36136
rect 99790 36078 102751 36080
rect 102685 36075 102751 36078
rect 195973 35866 196039 35869
rect 195973 35864 199394 35866
rect 195973 35808 195978 35864
rect 196034 35808 199394 35864
rect 195973 35806 199394 35808
rect 195973 35803 196039 35806
rect 199334 35768 199394 35806
rect 196065 35458 196131 35461
rect 196065 35456 199394 35458
rect 196065 35400 196070 35456
rect 196126 35400 199394 35456
rect 196065 35398 199394 35400
rect 196065 35395 196131 35398
rect 99790 34642 99850 35224
rect 199334 34952 199394 35398
rect 102133 34642 102199 34645
rect 99790 34640 102199 34642
rect 99790 34584 102138 34640
rect 102194 34584 102199 34640
rect 99790 34582 102199 34584
rect 102133 34579 102199 34582
rect 195973 34370 196039 34373
rect 195973 34368 199394 34370
rect 195973 34312 195978 34368
rect 196034 34312 199394 34368
rect 195973 34310 199394 34312
rect 195973 34307 196039 34310
rect 199334 34136 199394 34310
rect 99790 33554 99850 34136
rect 196065 33962 196131 33965
rect 196065 33960 199394 33962
rect 196065 33904 196070 33960
rect 196126 33904 199394 33960
rect 196065 33902 199394 33904
rect 196065 33899 196131 33902
rect 102317 33554 102383 33557
rect 99790 33552 102383 33554
rect 99790 33496 102322 33552
rect 102378 33496 102383 33552
rect 99790 33494 102383 33496
rect 102317 33491 102383 33494
rect 199334 33320 199394 33902
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect 99790 32466 99850 33048
rect 195973 33010 196039 33013
rect 195973 33008 199394 33010
rect 195973 32952 195978 33008
rect 196034 32952 199394 33008
rect 583520 32996 584960 33236
rect 195973 32950 199394 32952
rect 195973 32947 196039 32950
rect 199334 32504 199394 32950
rect 102133 32466 102199 32469
rect 99790 32464 102199 32466
rect 99790 32408 102138 32464
rect 102194 32408 102199 32464
rect 99790 32406 102199 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 102133 32403 102199 32406
rect 99790 31786 99850 31960
rect 102225 31786 102291 31789
rect 99790 31784 102291 31786
rect 99790 31728 102230 31784
rect 102286 31728 102291 31784
rect 99790 31726 102291 31728
rect 102225 31723 102291 31726
rect 57605 31650 57671 31653
rect 60046 31650 60106 31688
rect 57605 31648 60106 31650
rect 57605 31592 57610 31648
rect 57666 31592 60106 31648
rect 57605 31590 60106 31592
rect 195973 31650 196039 31653
rect 199334 31650 199394 31688
rect 195973 31648 199394 31650
rect 195973 31592 195978 31648
rect 196034 31592 199394 31648
rect 195973 31590 199394 31592
rect 57605 31587 57671 31590
rect 195973 31587 196039 31590
rect 196065 31514 196131 31517
rect 196065 31512 199394 31514
rect 196065 31456 196070 31512
rect 196126 31456 199394 31512
rect 196065 31454 199394 31456
rect 196065 31451 196131 31454
rect 199334 30872 199394 31454
rect 99790 30562 99850 30872
rect 102133 30562 102199 30565
rect 99790 30560 102199 30562
rect 99790 30504 102138 30560
rect 102194 30504 102199 30560
rect 99790 30502 102199 30504
rect 102133 30499 102199 30502
rect 195973 30154 196039 30157
rect 195973 30152 199394 30154
rect 195973 30096 195978 30152
rect 196034 30096 199394 30152
rect 195973 30094 199394 30096
rect 195973 30091 196039 30094
rect 199334 30056 199394 30094
rect 99790 29338 99850 29784
rect 196065 29746 196131 29749
rect 196065 29744 199394 29746
rect 196065 29688 196070 29744
rect 196126 29688 199394 29744
rect 196065 29686 199394 29688
rect 196065 29683 196131 29686
rect 102133 29338 102199 29341
rect 99790 29336 102199 29338
rect 99790 29280 102138 29336
rect 102194 29280 102199 29336
rect 99790 29278 102199 29280
rect 102133 29275 102199 29278
rect 199334 29240 199394 29686
rect 195973 28930 196039 28933
rect 195973 28928 199394 28930
rect 195973 28872 195978 28928
rect 196034 28872 199394 28928
rect 195973 28870 199394 28872
rect 195973 28867 196039 28870
rect 99790 28522 99850 28696
rect 102133 28522 102199 28525
rect 99790 28520 102199 28522
rect 99790 28464 102138 28520
rect 102194 28464 102199 28520
rect 99790 28462 102199 28464
rect 102133 28459 102199 28462
rect 199334 28424 199394 28870
rect 195973 28114 196039 28117
rect 195973 28112 199394 28114
rect 195973 28056 195978 28112
rect 196034 28056 199394 28112
rect 195973 28054 199394 28056
rect 195973 28051 196039 28054
rect 102133 27706 102199 27709
rect 99790 27704 102199 27706
rect 99790 27648 102138 27704
rect 102194 27648 102199 27704
rect 99790 27646 102199 27648
rect 99790 27608 99850 27646
rect 102133 27643 102199 27646
rect 199334 27608 199394 28054
rect 195973 27298 196039 27301
rect 195973 27296 199394 27298
rect 195973 27240 195978 27296
rect 196034 27240 199394 27296
rect 195973 27238 199394 27240
rect 195973 27235 196039 27238
rect 57237 27162 57303 27165
rect 57237 27160 60106 27162
rect 57237 27104 57242 27160
rect 57298 27104 60106 27160
rect 57237 27102 60106 27104
rect 57237 27099 57303 27102
rect 60046 26792 60106 27102
rect 199334 26792 199394 27238
rect 99790 26346 99850 26520
rect 102777 26346 102843 26349
rect 99790 26344 102843 26346
rect 99790 26288 102782 26344
rect 102838 26288 102843 26344
rect 99790 26286 102843 26288
rect 102777 26283 102843 26286
rect 195973 26210 196039 26213
rect 195973 26208 199394 26210
rect 195973 26152 195978 26208
rect 196034 26152 199394 26208
rect 195973 26150 199394 26152
rect 195973 26147 196039 26150
rect 199334 25976 199394 26150
rect 390001 24170 390067 24173
rect 420126 24170 420132 24172
rect 390001 24168 420132 24170
rect 390001 24112 390006 24168
rect 390062 24112 420132 24168
rect 390001 24110 420132 24112
rect 390001 24107 390067 24110
rect 420126 24108 420132 24110
rect 420196 24108 420202 24172
rect 393221 22130 393287 22133
rect 418654 22130 418660 22132
rect 393221 22128 418660 22130
rect 393221 22072 393226 22128
rect 393282 22072 418660 22128
rect 393221 22070 418660 22072
rect 393221 22067 393287 22070
rect 418654 22068 418660 22070
rect 418724 22068 418730 22132
rect 19558 21932 19564 21996
rect 19628 21994 19634 21996
rect 368105 21994 368171 21997
rect 19628 21992 368171 21994
rect 19628 21936 368110 21992
rect 368166 21936 368171 21992
rect 19628 21934 368171 21936
rect 19628 21932 19634 21934
rect 368105 21931 368171 21934
rect 382457 21994 382523 21997
rect 418102 21994 418108 21996
rect 382457 21992 418108 21994
rect 382457 21936 382462 21992
rect 382518 21936 418108 21992
rect 382457 21934 418108 21936
rect 382457 21931 382523 21934
rect 418102 21932 418108 21934
rect 418172 21932 418178 21996
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 418108 699816 418172 699820
rect 418108 699760 418158 699816
rect 418158 699760 418172 699816
rect 418108 699756 418172 699760
rect 17172 670652 17236 670716
rect 420132 591228 420196 591292
rect 303476 585924 303540 585988
rect 422340 585788 422404 585852
rect 299980 585652 300044 585716
rect 23244 582932 23308 582996
rect 299244 582932 299308 582996
rect 301452 580212 301516 580276
rect 138060 541724 138124 541788
rect 19564 502420 19628 502484
rect 418660 485012 418724 485076
rect 303476 461076 303540 461140
rect 142108 461000 142172 461004
rect 142108 460944 142122 461000
rect 142122 460944 142172 461000
rect 142108 460940 142172 460944
rect 23244 460124 23308 460188
rect 302740 459640 302804 459644
rect 302740 459584 302754 459640
rect 302754 459584 302804 459640
rect 302740 459580 302804 459584
rect 138060 458900 138124 458964
rect 23244 458280 23308 458284
rect 23244 458224 23258 458280
rect 23258 458224 23308 458280
rect 23244 458220 23308 458224
rect 138612 458220 138676 458284
rect 299244 458220 299308 458284
rect 421052 458220 421116 458284
rect 301452 456784 301516 456788
rect 301452 456728 301502 456784
rect 301502 456728 301516 456784
rect 301452 456724 301516 456728
rect 302004 418236 302068 418300
rect 138060 413884 138124 413948
rect 19380 357444 19444 357508
rect 17172 333916 17236 333980
rect 23244 332284 23308 332348
rect 302924 332284 302988 332348
rect 419580 331332 419644 331396
rect 19380 331196 19444 331260
rect 302740 331060 302804 331124
rect 21220 329700 21284 329764
rect 138060 329700 138124 329764
rect 141924 329700 141988 329764
rect 419580 204308 419644 204372
rect 21220 204172 21284 204236
rect 23244 203492 23308 203556
rect 302924 203764 302988 203828
rect 23244 202328 23308 202332
rect 23244 202272 23294 202328
rect 23294 202272 23308 202328
rect 23244 202268 23308 202272
rect 302740 158612 302804 158676
rect 302004 78568 302068 78572
rect 302004 78512 302054 78568
rect 302054 78512 302068 78568
rect 302004 78508 302068 78512
rect 299980 77828 300044 77892
rect 421052 76740 421116 76804
rect 303108 76604 303172 76668
rect 422340 76604 422404 76668
rect 138612 76468 138676 76532
rect 21956 75652 22020 75716
rect 98500 75108 98564 75172
rect 23244 74156 23308 74220
rect 98684 65452 98748 65516
rect 98500 61644 98564 61708
rect 302740 60556 302804 60620
rect 99420 57292 99484 57356
rect 420132 24108 420196 24172
rect 418660 22068 418724 22132
rect 19564 21932 19628 21996
rect 418108 21932 418172 21996
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 17171 670716 17237 670717
rect 17171 670652 17172 670716
rect 17236 670652 17237 670716
rect 17171 670651 17237 670652
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 17174 333981 17234 670651
rect 24294 670000 24914 673398
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 670000 29414 677898
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 670000 33914 682398
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 670000 38414 686898
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 670000 42914 691398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 670000 47414 695898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 670000 51914 700398
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 670000 60914 673398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 670000 65414 677898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 670000 69914 682398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 670000 74414 686898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 670000 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 670000 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 670000 87914 700398
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 670000 96914 673398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 670000 101414 677898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 670000 105914 682398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 670000 110414 686898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 670000 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 670000 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 670000 123914 700398
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 670000 132914 673398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 670000 137414 677898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 670000 141914 682398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 33868 655954 34868 655986
rect 33868 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 34868 655954
rect 33868 655634 34868 655718
rect 33868 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 34868 655634
rect 33868 655366 34868 655398
rect 53868 655954 54868 655986
rect 53868 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 54868 655954
rect 53868 655634 54868 655718
rect 53868 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 54868 655634
rect 53868 655366 54868 655398
rect 73868 655954 74868 655986
rect 73868 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 74868 655954
rect 73868 655634 74868 655718
rect 73868 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 74868 655634
rect 73868 655366 74868 655398
rect 93868 655954 94868 655986
rect 93868 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 94868 655954
rect 93868 655634 94868 655718
rect 93868 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 94868 655634
rect 93868 655366 94868 655398
rect 113868 655954 114868 655986
rect 113868 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 114868 655954
rect 113868 655634 114868 655718
rect 113868 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 114868 655634
rect 113868 655366 114868 655398
rect 133868 655954 134868 655986
rect 133868 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 134868 655954
rect 133868 655634 134868 655718
rect 133868 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 134868 655634
rect 133868 655366 134868 655398
rect 23868 651454 24868 651486
rect 23868 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 24868 651454
rect 23868 651134 24868 651218
rect 23868 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 24868 651134
rect 23868 650866 24868 650898
rect 43868 651454 44868 651486
rect 43868 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 44868 651454
rect 43868 651134 44868 651218
rect 43868 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 44868 651134
rect 43868 650866 44868 650898
rect 63868 651454 64868 651486
rect 63868 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 64868 651454
rect 63868 651134 64868 651218
rect 63868 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 64868 651134
rect 63868 650866 64868 650898
rect 83868 651454 84868 651486
rect 83868 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 84868 651454
rect 83868 651134 84868 651218
rect 83868 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 84868 651134
rect 83868 650866 84868 650898
rect 103868 651454 104868 651486
rect 103868 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 104868 651454
rect 103868 651134 104868 651218
rect 103868 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 104868 651134
rect 103868 650866 104868 650898
rect 123868 651454 124868 651486
rect 123868 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 124868 651454
rect 123868 651134 124868 651218
rect 123868 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 124868 651134
rect 123868 650866 124868 650898
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 33868 619954 34868 619986
rect 33868 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 34868 619954
rect 33868 619634 34868 619718
rect 33868 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 34868 619634
rect 33868 619366 34868 619398
rect 53868 619954 54868 619986
rect 53868 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 54868 619954
rect 53868 619634 54868 619718
rect 53868 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 54868 619634
rect 53868 619366 54868 619398
rect 73868 619954 74868 619986
rect 73868 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 74868 619954
rect 73868 619634 74868 619718
rect 73868 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 74868 619634
rect 73868 619366 74868 619398
rect 93868 619954 94868 619986
rect 93868 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 94868 619954
rect 93868 619634 94868 619718
rect 93868 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 94868 619634
rect 93868 619366 94868 619398
rect 113868 619954 114868 619986
rect 113868 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 114868 619954
rect 113868 619634 114868 619718
rect 113868 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 114868 619634
rect 113868 619366 114868 619398
rect 133868 619954 134868 619986
rect 133868 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 134868 619954
rect 133868 619634 134868 619718
rect 133868 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 134868 619634
rect 133868 619366 134868 619398
rect 23868 615454 24868 615486
rect 23868 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 24868 615454
rect 23868 615134 24868 615218
rect 23868 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 24868 615134
rect 23868 614866 24868 614898
rect 43868 615454 44868 615486
rect 43868 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 44868 615454
rect 43868 615134 44868 615218
rect 43868 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 44868 615134
rect 43868 614866 44868 614898
rect 63868 615454 64868 615486
rect 63868 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 64868 615454
rect 63868 615134 64868 615218
rect 63868 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 64868 615134
rect 63868 614866 64868 614898
rect 83868 615454 84868 615486
rect 83868 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 84868 615454
rect 83868 615134 84868 615218
rect 83868 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 84868 615134
rect 83868 614866 84868 614898
rect 103868 615454 104868 615486
rect 103868 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 104868 615454
rect 103868 615134 104868 615218
rect 103868 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 104868 615134
rect 103868 614866 104868 614898
rect 123868 615454 124868 615486
rect 123868 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 124868 615454
rect 123868 615134 124868 615218
rect 123868 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 124868 615134
rect 123868 614866 124868 614898
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 42294 583954 42914 586000
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 23243 582996 23309 582997
rect 23243 582932 23244 582996
rect 23308 582932 23309 582996
rect 23243 582931 23309 582932
rect 19563 502484 19629 502485
rect 19563 502420 19564 502484
rect 19628 502420 19629 502484
rect 19563 502419 19629 502420
rect 19379 357508 19445 357509
rect 19379 357444 19380 357508
rect 19444 357444 19445 357508
rect 19379 357443 19445 357444
rect 17171 333980 17237 333981
rect 17171 333916 17172 333980
rect 17236 333916 17237 333980
rect 17171 333915 17237 333916
rect 19382 331261 19442 357443
rect 19379 331260 19445 331261
rect 19379 331196 19380 331260
rect 19444 331196 19445 331260
rect 19379 331195 19445 331196
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 19566 21997 19626 502419
rect 23246 460189 23306 582931
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 544000 42914 547398
rect 78294 583954 78914 586000
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 544000 78914 547398
rect 114294 583954 114914 586000
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 544000 114914 547398
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 138059 541788 138125 541789
rect 138059 541724 138060 541788
rect 138124 541724 138125 541788
rect 138059 541723 138125 541724
rect 33868 511954 34868 511986
rect 33868 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 34868 511954
rect 33868 511634 34868 511718
rect 33868 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 34868 511634
rect 33868 511366 34868 511398
rect 53868 511954 54868 511986
rect 53868 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 54868 511954
rect 53868 511634 54868 511718
rect 53868 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 54868 511634
rect 53868 511366 54868 511398
rect 73868 511954 74868 511986
rect 73868 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 74868 511954
rect 73868 511634 74868 511718
rect 73868 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 74868 511634
rect 73868 511366 74868 511398
rect 93868 511954 94868 511986
rect 93868 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 94868 511954
rect 93868 511634 94868 511718
rect 93868 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 94868 511634
rect 93868 511366 94868 511398
rect 113868 511954 114868 511986
rect 113868 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 114868 511954
rect 113868 511634 114868 511718
rect 113868 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 114868 511634
rect 113868 511366 114868 511398
rect 133868 511954 134868 511986
rect 133868 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 134868 511954
rect 133868 511634 134868 511718
rect 133868 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 134868 511634
rect 133868 511366 134868 511398
rect 23868 507454 24868 507486
rect 23868 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 24868 507454
rect 23868 507134 24868 507218
rect 23868 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 24868 507134
rect 23868 506866 24868 506898
rect 43868 507454 44868 507486
rect 43868 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 44868 507454
rect 43868 507134 44868 507218
rect 43868 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 44868 507134
rect 43868 506866 44868 506898
rect 63868 507454 64868 507486
rect 63868 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 64868 507454
rect 63868 507134 64868 507218
rect 63868 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 64868 507134
rect 63868 506866 64868 506898
rect 83868 507454 84868 507486
rect 83868 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 84868 507454
rect 83868 507134 84868 507218
rect 83868 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 84868 507134
rect 83868 506866 84868 506898
rect 103868 507454 104868 507486
rect 103868 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 104868 507454
rect 103868 507134 104868 507218
rect 103868 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 104868 507134
rect 103868 506866 104868 506898
rect 123868 507454 124868 507486
rect 123868 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 124868 507454
rect 123868 507134 124868 507218
rect 123868 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 124868 507134
rect 123868 506866 124868 506898
rect 33868 475954 34868 475986
rect 33868 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 34868 475954
rect 33868 475634 34868 475718
rect 33868 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 34868 475634
rect 33868 475366 34868 475398
rect 53868 475954 54868 475986
rect 53868 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 54868 475954
rect 53868 475634 54868 475718
rect 53868 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 54868 475634
rect 53868 475366 54868 475398
rect 73868 475954 74868 475986
rect 73868 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 74868 475954
rect 73868 475634 74868 475718
rect 73868 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 74868 475634
rect 73868 475366 74868 475398
rect 93868 475954 94868 475986
rect 93868 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 94868 475954
rect 93868 475634 94868 475718
rect 93868 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 94868 475634
rect 93868 475366 94868 475398
rect 113868 475954 114868 475986
rect 113868 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 114868 475954
rect 113868 475634 114868 475718
rect 113868 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 114868 475634
rect 113868 475366 114868 475398
rect 133868 475954 134868 475986
rect 133868 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 134868 475954
rect 133868 475634 134868 475718
rect 133868 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 134868 475634
rect 133868 475366 134868 475398
rect 23868 471454 24868 471486
rect 23868 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 24868 471454
rect 23868 471134 24868 471218
rect 23868 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 24868 471134
rect 23868 470866 24868 470898
rect 43868 471454 44868 471486
rect 43868 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 44868 471454
rect 43868 471134 44868 471218
rect 43868 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 44868 471134
rect 43868 470866 44868 470898
rect 63868 471454 64868 471486
rect 63868 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 64868 471454
rect 63868 471134 64868 471218
rect 63868 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 64868 471134
rect 63868 470866 64868 470898
rect 83868 471454 84868 471486
rect 83868 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 84868 471454
rect 83868 471134 84868 471218
rect 83868 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 84868 471134
rect 83868 470866 84868 470898
rect 103868 471454 104868 471486
rect 103868 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 104868 471454
rect 103868 471134 104868 471218
rect 103868 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 104868 471134
rect 103868 470866 104868 470898
rect 123868 471454 124868 471486
rect 123868 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 124868 471454
rect 123868 471134 124868 471218
rect 123868 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 124868 471134
rect 123868 470866 124868 470898
rect 23243 460188 23309 460189
rect 23243 460124 23244 460188
rect 23308 460124 23309 460188
rect 23243 460123 23309 460124
rect 19794 453454 20414 460000
rect 23243 458284 23309 458285
rect 23243 458220 23244 458284
rect 23308 458220 23309 458284
rect 23243 458219 23309 458220
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 416000 20414 416898
rect 23246 332349 23306 458219
rect 24294 457954 24914 460000
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 416000 24914 421398
rect 55794 453454 56414 460000
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 416000 56414 416898
rect 60294 457954 60914 460000
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 416000 60914 421398
rect 91794 453454 92414 460000
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 416000 92414 416898
rect 96294 457954 96914 460000
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 416000 96914 421398
rect 127794 453454 128414 460000
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 416000 128414 416898
rect 132294 457954 132914 460000
rect 138062 458965 138122 541723
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 142107 461004 142173 461005
rect 142107 460950 142108 461004
rect 141926 460940 142108 460950
rect 142172 460940 142173 461004
rect 141926 460939 142173 460940
rect 141926 460890 142170 460939
rect 138059 458964 138125 458965
rect 138059 458900 138060 458964
rect 138124 458900 138125 458964
rect 138059 458899 138125 458900
rect 138611 458284 138677 458285
rect 138611 458220 138612 458284
rect 138676 458220 138677 458284
rect 138611 458219 138677 458220
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 416000 132914 421398
rect 138059 413948 138125 413949
rect 138059 413884 138060 413948
rect 138124 413884 138125 413948
rect 138059 413883 138125 413884
rect 33868 403954 34868 403986
rect 33868 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 34868 403954
rect 33868 403634 34868 403718
rect 33868 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 34868 403634
rect 33868 403366 34868 403398
rect 53868 403954 54868 403986
rect 53868 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 54868 403954
rect 53868 403634 54868 403718
rect 53868 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 54868 403634
rect 53868 403366 54868 403398
rect 73868 403954 74868 403986
rect 73868 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 74868 403954
rect 73868 403634 74868 403718
rect 73868 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 74868 403634
rect 73868 403366 74868 403398
rect 93868 403954 94868 403986
rect 93868 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 94868 403954
rect 93868 403634 94868 403718
rect 93868 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 94868 403634
rect 93868 403366 94868 403398
rect 113868 403954 114868 403986
rect 113868 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 114868 403954
rect 113868 403634 114868 403718
rect 113868 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 114868 403634
rect 113868 403366 114868 403398
rect 133868 403954 134868 403986
rect 133868 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 134868 403954
rect 133868 403634 134868 403718
rect 133868 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 134868 403634
rect 133868 403366 134868 403398
rect 23868 399454 24868 399486
rect 23868 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 24868 399454
rect 23868 399134 24868 399218
rect 23868 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 24868 399134
rect 23868 398866 24868 398898
rect 43868 399454 44868 399486
rect 43868 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 44868 399454
rect 43868 399134 44868 399218
rect 43868 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 44868 399134
rect 43868 398866 44868 398898
rect 63868 399454 64868 399486
rect 63868 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 64868 399454
rect 63868 399134 64868 399218
rect 63868 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 64868 399134
rect 63868 398866 64868 398898
rect 83868 399454 84868 399486
rect 83868 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 84868 399454
rect 83868 399134 84868 399218
rect 83868 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 84868 399134
rect 83868 398866 84868 398898
rect 103868 399454 104868 399486
rect 103868 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 104868 399454
rect 103868 399134 104868 399218
rect 103868 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 104868 399134
rect 103868 398866 104868 398898
rect 123868 399454 124868 399486
rect 123868 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 124868 399454
rect 123868 399134 124868 399218
rect 123868 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 124868 399134
rect 123868 398866 124868 398898
rect 33868 367954 34868 367986
rect 33868 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 34868 367954
rect 33868 367634 34868 367718
rect 33868 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 34868 367634
rect 33868 367366 34868 367398
rect 53868 367954 54868 367986
rect 53868 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 54868 367954
rect 53868 367634 54868 367718
rect 53868 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 54868 367634
rect 53868 367366 54868 367398
rect 73868 367954 74868 367986
rect 73868 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 74868 367954
rect 73868 367634 74868 367718
rect 73868 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 74868 367634
rect 73868 367366 74868 367398
rect 93868 367954 94868 367986
rect 93868 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 94868 367954
rect 93868 367634 94868 367718
rect 93868 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 94868 367634
rect 93868 367366 94868 367398
rect 113868 367954 114868 367986
rect 113868 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 114868 367954
rect 113868 367634 114868 367718
rect 113868 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 114868 367634
rect 113868 367366 114868 367398
rect 133868 367954 134868 367986
rect 133868 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 134868 367954
rect 133868 367634 134868 367718
rect 133868 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 134868 367634
rect 133868 367366 134868 367398
rect 23868 363454 24868 363486
rect 23868 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 24868 363454
rect 23868 363134 24868 363218
rect 23868 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 24868 363134
rect 23868 362866 24868 362898
rect 43868 363454 44868 363486
rect 43868 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 44868 363454
rect 43868 363134 44868 363218
rect 43868 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 44868 363134
rect 43868 362866 44868 362898
rect 63868 363454 64868 363486
rect 63868 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 64868 363454
rect 63868 363134 64868 363218
rect 63868 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 64868 363134
rect 63868 362866 64868 362898
rect 83868 363454 84868 363486
rect 83868 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 84868 363454
rect 83868 363134 84868 363218
rect 83868 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 84868 363134
rect 83868 362866 84868 362898
rect 103868 363454 104868 363486
rect 103868 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 104868 363454
rect 103868 363134 104868 363218
rect 103868 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 104868 363134
rect 103868 362866 104868 362898
rect 123868 363454 124868 363486
rect 123868 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 124868 363454
rect 123868 363134 124868 363218
rect 123868 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 124868 363134
rect 123868 362866 124868 362898
rect 23243 332348 23309 332349
rect 23243 332284 23244 332348
rect 23308 332284 23309 332348
rect 23243 332283 23309 332284
rect 21219 329764 21285 329765
rect 21219 329700 21220 329764
rect 21284 329700 21285 329764
rect 21219 329699 21285 329700
rect 21222 204237 21282 329699
rect 21219 204236 21285 204237
rect 21219 204172 21220 204236
rect 21284 204172 21285 204236
rect 21219 204171 21285 204172
rect 19794 201454 20414 204000
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 21222 200130 21282 204171
rect 23246 203557 23306 332283
rect 37794 327454 38414 332000
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 288000 38414 290898
rect 42294 331954 42914 332000
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 288000 42914 295398
rect 73794 327454 74414 332000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 288000 74414 290898
rect 78294 331954 78914 332000
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 288000 78914 295398
rect 109794 327454 110414 332000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 288000 110414 290898
rect 114294 331954 114914 332000
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 138062 329765 138122 413883
rect 138059 329764 138125 329765
rect 138059 329700 138060 329764
rect 138124 329700 138125 329764
rect 138059 329699 138125 329700
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 288000 114914 295398
rect 33868 259954 34868 259986
rect 33868 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 34868 259954
rect 33868 259634 34868 259718
rect 33868 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 34868 259634
rect 33868 259366 34868 259398
rect 53868 259954 54868 259986
rect 53868 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 54868 259954
rect 53868 259634 54868 259718
rect 53868 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 54868 259634
rect 53868 259366 54868 259398
rect 73868 259954 74868 259986
rect 73868 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 74868 259954
rect 73868 259634 74868 259718
rect 73868 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 74868 259634
rect 73868 259366 74868 259398
rect 93868 259954 94868 259986
rect 93868 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 94868 259954
rect 93868 259634 94868 259718
rect 93868 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 94868 259634
rect 93868 259366 94868 259398
rect 113868 259954 114868 259986
rect 113868 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 114868 259954
rect 113868 259634 114868 259718
rect 113868 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 114868 259634
rect 113868 259366 114868 259398
rect 133868 259954 134868 259986
rect 133868 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 134868 259954
rect 133868 259634 134868 259718
rect 133868 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 134868 259634
rect 133868 259366 134868 259398
rect 23868 255454 24868 255486
rect 23868 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 24868 255454
rect 23868 255134 24868 255218
rect 23868 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 24868 255134
rect 23868 254866 24868 254898
rect 43868 255454 44868 255486
rect 43868 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 44868 255454
rect 43868 255134 44868 255218
rect 43868 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 44868 255134
rect 43868 254866 44868 254898
rect 63868 255454 64868 255486
rect 63868 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 64868 255454
rect 63868 255134 64868 255218
rect 63868 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 64868 255134
rect 63868 254866 64868 254898
rect 83868 255454 84868 255486
rect 83868 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 84868 255454
rect 83868 255134 84868 255218
rect 83868 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 84868 255134
rect 83868 254866 84868 254898
rect 103868 255454 104868 255486
rect 103868 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 104868 255454
rect 103868 255134 104868 255218
rect 103868 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 104868 255134
rect 103868 254866 104868 254898
rect 123868 255454 124868 255486
rect 123868 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 124868 255454
rect 123868 255134 124868 255218
rect 123868 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 124868 255134
rect 123868 254866 124868 254898
rect 33868 223954 34868 223986
rect 33868 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 34868 223954
rect 33868 223634 34868 223718
rect 33868 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 34868 223634
rect 33868 223366 34868 223398
rect 53868 223954 54868 223986
rect 53868 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 54868 223954
rect 53868 223634 54868 223718
rect 53868 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 54868 223634
rect 53868 223366 54868 223398
rect 73868 223954 74868 223986
rect 73868 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 74868 223954
rect 73868 223634 74868 223718
rect 73868 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 74868 223634
rect 73868 223366 74868 223398
rect 93868 223954 94868 223986
rect 93868 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 94868 223954
rect 93868 223634 94868 223718
rect 93868 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 94868 223634
rect 93868 223366 94868 223398
rect 113868 223954 114868 223986
rect 113868 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 114868 223954
rect 113868 223634 114868 223718
rect 113868 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 114868 223634
rect 113868 223366 114868 223398
rect 133868 223954 134868 223986
rect 133868 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 134868 223954
rect 133868 223634 134868 223718
rect 133868 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 134868 223634
rect 133868 223366 134868 223398
rect 23868 219454 24868 219486
rect 23868 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 24868 219454
rect 23868 219134 24868 219218
rect 23868 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 24868 219134
rect 23868 218866 24868 218898
rect 43868 219454 44868 219486
rect 43868 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 44868 219454
rect 43868 219134 44868 219218
rect 43868 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 44868 219134
rect 43868 218866 44868 218898
rect 63868 219454 64868 219486
rect 63868 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 64868 219454
rect 63868 219134 64868 219218
rect 63868 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 64868 219134
rect 63868 218866 64868 218898
rect 83868 219454 84868 219486
rect 83868 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 84868 219454
rect 83868 219134 84868 219218
rect 83868 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 84868 219134
rect 83868 218866 84868 218898
rect 103868 219454 104868 219486
rect 103868 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 104868 219454
rect 103868 219134 104868 219218
rect 103868 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 104868 219134
rect 103868 218866 104868 218898
rect 123868 219454 124868 219486
rect 123868 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 124868 219454
rect 123868 219134 124868 219218
rect 123868 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 124868 219134
rect 123868 218866 124868 218898
rect 23243 203556 23309 203557
rect 23243 203492 23244 203556
rect 23308 203492 23309 203556
rect 23243 203491 23309 203492
rect 23243 202332 23309 202333
rect 23243 202268 23244 202332
rect 23308 202268 23309 202332
rect 23243 202267 23309 202268
rect 21222 200070 22018 200130
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 160000 20414 164898
rect 19794 57454 20414 76000
rect 21958 75717 22018 200070
rect 21955 75716 22021 75717
rect 21955 75652 21956 75716
rect 22020 75652 22021 75716
rect 21955 75651 22021 75652
rect 23246 74221 23306 202267
rect 51294 196954 51914 204000
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 160000 51914 160398
rect 55794 201454 56414 204000
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 160000 56414 164898
rect 87294 196954 87914 204000
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 160000 87914 160398
rect 91794 201454 92414 204000
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 160000 92414 164898
rect 123294 196954 123914 204000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 160000 123914 160398
rect 127794 201454 128414 204000
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 160000 128414 164898
rect 33868 151954 34868 151986
rect 33868 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 34868 151954
rect 33868 151634 34868 151718
rect 33868 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 34868 151634
rect 33868 151366 34868 151398
rect 53868 151954 54868 151986
rect 53868 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 54868 151954
rect 53868 151634 54868 151718
rect 53868 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 54868 151634
rect 53868 151366 54868 151398
rect 73868 151954 74868 151986
rect 73868 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 74868 151954
rect 73868 151634 74868 151718
rect 73868 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 74868 151634
rect 73868 151366 74868 151398
rect 93868 151954 94868 151986
rect 93868 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 94868 151954
rect 93868 151634 94868 151718
rect 93868 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 94868 151634
rect 93868 151366 94868 151398
rect 113868 151954 114868 151986
rect 113868 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 114868 151954
rect 113868 151634 114868 151718
rect 113868 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 114868 151634
rect 113868 151366 114868 151398
rect 133868 151954 134868 151986
rect 133868 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 134868 151954
rect 133868 151634 134868 151718
rect 133868 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 134868 151634
rect 133868 151366 134868 151398
rect 23868 147454 24868 147486
rect 23868 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 24868 147454
rect 23868 147134 24868 147218
rect 23868 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 24868 147134
rect 23868 146866 24868 146898
rect 43868 147454 44868 147486
rect 43868 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 44868 147454
rect 43868 147134 44868 147218
rect 43868 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 44868 147134
rect 43868 146866 44868 146898
rect 63868 147454 64868 147486
rect 63868 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 64868 147454
rect 63868 147134 64868 147218
rect 63868 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 64868 147134
rect 63868 146866 64868 146898
rect 83868 147454 84868 147486
rect 83868 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 84868 147454
rect 83868 147134 84868 147218
rect 83868 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 84868 147134
rect 83868 146866 84868 146898
rect 103868 147454 104868 147486
rect 103868 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 104868 147454
rect 103868 147134 104868 147218
rect 103868 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 104868 147134
rect 103868 146866 104868 146898
rect 123868 147454 124868 147486
rect 123868 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 124868 147454
rect 123868 147134 124868 147218
rect 123868 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 124868 147134
rect 123868 146866 124868 146898
rect 33868 115954 34868 115986
rect 33868 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 34868 115954
rect 33868 115634 34868 115718
rect 33868 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 34868 115634
rect 33868 115366 34868 115398
rect 53868 115954 54868 115986
rect 53868 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 54868 115954
rect 53868 115634 54868 115718
rect 53868 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 54868 115634
rect 53868 115366 54868 115398
rect 73868 115954 74868 115986
rect 73868 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 74868 115954
rect 73868 115634 74868 115718
rect 73868 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 74868 115634
rect 73868 115366 74868 115398
rect 93868 115954 94868 115986
rect 93868 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 94868 115954
rect 93868 115634 94868 115718
rect 93868 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 94868 115634
rect 93868 115366 94868 115398
rect 113868 115954 114868 115986
rect 113868 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 114868 115954
rect 113868 115634 114868 115718
rect 113868 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 114868 115634
rect 113868 115366 114868 115398
rect 133868 115954 134868 115986
rect 133868 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 134868 115954
rect 133868 115634 134868 115718
rect 133868 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 134868 115634
rect 133868 115366 134868 115398
rect 23868 111454 24868 111486
rect 23868 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 24868 111454
rect 23868 111134 24868 111218
rect 23868 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 24868 111134
rect 23868 110866 24868 110898
rect 43868 111454 44868 111486
rect 43868 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 44868 111454
rect 43868 111134 44868 111218
rect 43868 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 44868 111134
rect 43868 110866 44868 110898
rect 63868 111454 64868 111486
rect 63868 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 64868 111454
rect 63868 111134 64868 111218
rect 63868 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 64868 111134
rect 63868 110866 64868 110898
rect 83868 111454 84868 111486
rect 83868 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 84868 111454
rect 83868 111134 84868 111218
rect 83868 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 84868 111134
rect 83868 110866 84868 110898
rect 103868 111454 104868 111486
rect 103868 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 104868 111454
rect 103868 111134 104868 111218
rect 103868 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 104868 111134
rect 103868 110866 104868 110898
rect 123868 111454 124868 111486
rect 123868 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 124868 111454
rect 123868 111134 124868 111218
rect 123868 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 124868 111134
rect 123868 110866 124868 110898
rect 138614 76533 138674 458219
rect 141926 329765 141986 460890
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 141923 329764 141989 329765
rect 141923 329700 141924 329764
rect 141988 329700 141989 329764
rect 141923 329699 141989 329700
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 138611 76532 138677 76533
rect 138611 76468 138612 76532
rect 138676 76468 138677 76532
rect 138611 76467 138677 76468
rect 23243 74220 23309 74221
rect 23243 74156 23244 74220
rect 23308 74156 23309 74220
rect 23243 74155 23309 74156
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19563 21996 19629 21997
rect 19563 21932 19564 21996
rect 19628 21932 19629 21996
rect 19563 21931 19629 21932
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 61954 24914 76000
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 66454 29414 76000
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 70954 33914 76000
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 75454 38414 76000
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 43954 42914 76000
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 48454 47414 76000
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 52954 51914 76000
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 76000
rect 98499 75172 98565 75173
rect 98499 75108 98500 75172
rect 98564 75108 98565 75172
rect 98499 75107 98565 75108
rect 98502 61709 98562 75107
rect 105294 70954 105914 76000
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 98683 65516 98749 65517
rect 98683 65452 98684 65516
rect 98748 65452 98749 65516
rect 98683 65451 98749 65452
rect 98499 61708 98565 61709
rect 98499 61644 98500 61708
rect 98564 61644 98565 61708
rect 98499 61643 98565 61644
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 98686 57490 98746 65451
rect 98686 57430 99482 57490
rect 99422 57357 99482 57430
rect 99419 57356 99485 57357
rect 99419 57292 99420 57356
rect 99484 57292 99485 57356
rect 99419 57291 99485 57292
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 79568 43954 79888 43986
rect 79568 43718 79610 43954
rect 79846 43718 79888 43954
rect 79568 43634 79888 43718
rect 79568 43398 79610 43634
rect 79846 43398 79888 43634
rect 79568 43366 79888 43398
rect 64208 39454 64528 39486
rect 64208 39218 64250 39454
rect 64486 39218 64528 39454
rect 64208 39134 64528 39218
rect 64208 38898 64250 39134
rect 64486 38898 64528 39134
rect 64208 38866 64528 38898
rect 94928 39454 95248 39486
rect 94928 39218 94970 39454
rect 95206 39218 95248 39454
rect 94928 39134 95248 39218
rect 94928 38898 94970 39134
rect 95206 38898 95248 39134
rect 94928 38866 95248 38898
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 73794 3454 74414 22000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 22000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 22000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 22000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 21454 92414 22000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 76000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 76000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 76000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 76000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 76000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 76000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 76000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 76000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 56000 200414 56898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 56000 204914 61398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 56000 209414 65898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 56000 213914 70398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 56000 218414 74898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 56000 222914 79398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 56000 227414 83898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 56000 231914 88398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 56000 236414 56898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 56000 240914 61398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 56000 245414 65898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 56000 249914 70398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 56000 254414 74898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 56000 258914 79398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 56000 263414 83898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 56000 267914 88398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 56000 272414 56898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 56000 276914 61398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 56000 281414 65898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 56000 285914 70398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 56000 290414 74898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 670000 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 670000 303914 700398
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 670000 312914 673398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 670000 317414 677898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 670000 321914 682398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 670000 326414 686898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 670000 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 670000 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 670000 339914 700398
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 670000 348914 673398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 670000 353414 677898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 670000 357914 682398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 670000 362414 686898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 670000 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 670000 371414 695898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 670000 375914 700398
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 670000 384914 673398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 670000 389414 677898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 670000 393914 682398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 670000 398414 686898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 670000 402914 691398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 670000 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 670000 411914 700398
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 418107 699820 418173 699821
rect 418107 699756 418108 699820
rect 418172 699756 418173 699820
rect 418107 699755 418173 699756
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 313868 655954 314868 655986
rect 313868 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 314868 655954
rect 313868 655634 314868 655718
rect 313868 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 314868 655634
rect 313868 655366 314868 655398
rect 333868 655954 334868 655986
rect 333868 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 334868 655954
rect 333868 655634 334868 655718
rect 333868 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 334868 655634
rect 333868 655366 334868 655398
rect 353868 655954 354868 655986
rect 353868 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 354868 655954
rect 353868 655634 354868 655718
rect 353868 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 354868 655634
rect 353868 655366 354868 655398
rect 373868 655954 374868 655986
rect 373868 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 374868 655954
rect 373868 655634 374868 655718
rect 373868 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 374868 655634
rect 373868 655366 374868 655398
rect 393868 655954 394868 655986
rect 393868 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 394868 655954
rect 393868 655634 394868 655718
rect 393868 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 394868 655634
rect 393868 655366 394868 655398
rect 413868 655954 414868 655986
rect 413868 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 414868 655954
rect 413868 655634 414868 655718
rect 413868 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 414868 655634
rect 413868 655366 414868 655398
rect 303868 651454 304868 651486
rect 303868 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 304868 651454
rect 303868 651134 304868 651218
rect 303868 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 304868 651134
rect 303868 650866 304868 650898
rect 323868 651454 324868 651486
rect 323868 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 324868 651454
rect 323868 651134 324868 651218
rect 323868 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 324868 651134
rect 323868 650866 324868 650898
rect 343868 651454 344868 651486
rect 343868 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 344868 651454
rect 343868 651134 344868 651218
rect 343868 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 344868 651134
rect 343868 650866 344868 650898
rect 363868 651454 364868 651486
rect 363868 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 364868 651454
rect 363868 651134 364868 651218
rect 363868 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 364868 651134
rect 363868 650866 364868 650898
rect 383868 651454 384868 651486
rect 383868 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 384868 651454
rect 383868 651134 384868 651218
rect 383868 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 384868 651134
rect 383868 650866 384868 650898
rect 403868 651454 404868 651486
rect 403868 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 404868 651454
rect 403868 651134 404868 651218
rect 403868 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 404868 651134
rect 403868 650866 404868 650898
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 313868 619954 314868 619986
rect 313868 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 314868 619954
rect 313868 619634 314868 619718
rect 313868 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 314868 619634
rect 313868 619366 314868 619398
rect 333868 619954 334868 619986
rect 333868 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 334868 619954
rect 333868 619634 334868 619718
rect 333868 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 334868 619634
rect 333868 619366 334868 619398
rect 353868 619954 354868 619986
rect 353868 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 354868 619954
rect 353868 619634 354868 619718
rect 353868 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 354868 619634
rect 353868 619366 354868 619398
rect 373868 619954 374868 619986
rect 373868 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 374868 619954
rect 373868 619634 374868 619718
rect 373868 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 374868 619634
rect 373868 619366 374868 619398
rect 393868 619954 394868 619986
rect 393868 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 394868 619954
rect 393868 619634 394868 619718
rect 393868 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 394868 619634
rect 393868 619366 394868 619398
rect 413868 619954 414868 619986
rect 413868 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 414868 619954
rect 413868 619634 414868 619718
rect 413868 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 414868 619634
rect 413868 619366 414868 619398
rect 303868 615454 304868 615486
rect 303868 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 304868 615454
rect 303868 615134 304868 615218
rect 303868 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 304868 615134
rect 303868 614866 304868 614898
rect 323868 615454 324868 615486
rect 323868 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 324868 615454
rect 323868 615134 324868 615218
rect 323868 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 324868 615134
rect 323868 614866 324868 614898
rect 343868 615454 344868 615486
rect 343868 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 344868 615454
rect 343868 615134 344868 615218
rect 343868 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 344868 615134
rect 343868 614866 344868 614898
rect 363868 615454 364868 615486
rect 363868 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 364868 615454
rect 363868 615134 364868 615218
rect 363868 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 364868 615134
rect 363868 614866 364868 614898
rect 383868 615454 384868 615486
rect 383868 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 384868 615454
rect 383868 615134 384868 615218
rect 383868 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 384868 615134
rect 383868 614866 384868 614898
rect 403868 615454 404868 615486
rect 403868 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 404868 615454
rect 403868 615134 404868 615218
rect 403868 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 404868 615134
rect 403868 614866 404868 614898
rect 303475 585988 303541 585989
rect 303475 585924 303476 585988
rect 303540 585924 303541 585988
rect 303475 585923 303541 585924
rect 299979 585716 300045 585717
rect 299979 585652 299980 585716
rect 300044 585652 300045 585716
rect 299979 585651 300045 585652
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 299243 582996 299309 582997
rect 299243 582932 299244 582996
rect 299308 582932 299309 582996
rect 299243 582931 299309 582932
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 299246 458285 299306 582931
rect 299243 458284 299309 458285
rect 299243 458220 299244 458284
rect 299308 458220 299309 458284
rect 299243 458219 299309 458220
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 56000 294914 79398
rect 299982 77893 300042 585651
rect 301451 580276 301517 580277
rect 301451 580212 301452 580276
rect 301516 580212 301517 580276
rect 301451 580211 301517 580212
rect 301454 456789 301514 580211
rect 303478 461141 303538 585923
rect 330294 583954 330914 586000
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 544000 330914 547398
rect 366294 583954 366914 586000
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 544000 366914 547398
rect 402294 583954 402914 586000
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 544000 402914 547398
rect 313868 511954 314868 511986
rect 313868 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 314868 511954
rect 313868 511634 314868 511718
rect 313868 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 314868 511634
rect 313868 511366 314868 511398
rect 333868 511954 334868 511986
rect 333868 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 334868 511954
rect 333868 511634 334868 511718
rect 333868 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 334868 511634
rect 333868 511366 334868 511398
rect 353868 511954 354868 511986
rect 353868 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 354868 511954
rect 353868 511634 354868 511718
rect 353868 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 354868 511634
rect 353868 511366 354868 511398
rect 373868 511954 374868 511986
rect 373868 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 374868 511954
rect 373868 511634 374868 511718
rect 373868 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 374868 511634
rect 373868 511366 374868 511398
rect 393868 511954 394868 511986
rect 393868 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 394868 511954
rect 393868 511634 394868 511718
rect 393868 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 394868 511634
rect 393868 511366 394868 511398
rect 413868 511954 414868 511986
rect 413868 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 414868 511954
rect 413868 511634 414868 511718
rect 413868 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 414868 511634
rect 413868 511366 414868 511398
rect 303868 507454 304868 507486
rect 303868 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 304868 507454
rect 303868 507134 304868 507218
rect 303868 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 304868 507134
rect 303868 506866 304868 506898
rect 323868 507454 324868 507486
rect 323868 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 324868 507454
rect 323868 507134 324868 507218
rect 323868 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 324868 507134
rect 323868 506866 324868 506898
rect 343868 507454 344868 507486
rect 343868 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 344868 507454
rect 343868 507134 344868 507218
rect 343868 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 344868 507134
rect 343868 506866 344868 506898
rect 363868 507454 364868 507486
rect 363868 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 364868 507454
rect 363868 507134 364868 507218
rect 363868 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 364868 507134
rect 363868 506866 364868 506898
rect 383868 507454 384868 507486
rect 383868 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 384868 507454
rect 383868 507134 384868 507218
rect 383868 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 384868 507134
rect 383868 506866 384868 506898
rect 403868 507454 404868 507486
rect 403868 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 404868 507454
rect 403868 507134 404868 507218
rect 403868 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 404868 507134
rect 403868 506866 404868 506898
rect 313868 475954 314868 475986
rect 313868 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 314868 475954
rect 313868 475634 314868 475718
rect 313868 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 314868 475634
rect 313868 475366 314868 475398
rect 333868 475954 334868 475986
rect 333868 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 334868 475954
rect 333868 475634 334868 475718
rect 333868 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 334868 475634
rect 333868 475366 334868 475398
rect 353868 475954 354868 475986
rect 353868 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 354868 475954
rect 353868 475634 354868 475718
rect 353868 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 354868 475634
rect 353868 475366 354868 475398
rect 373868 475954 374868 475986
rect 373868 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 374868 475954
rect 373868 475634 374868 475718
rect 373868 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 374868 475634
rect 373868 475366 374868 475398
rect 393868 475954 394868 475986
rect 393868 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 394868 475954
rect 393868 475634 394868 475718
rect 393868 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 394868 475634
rect 393868 475366 394868 475398
rect 413868 475954 414868 475986
rect 413868 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 414868 475954
rect 413868 475634 414868 475718
rect 413868 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 414868 475634
rect 413868 475366 414868 475398
rect 303868 471454 304868 471486
rect 303868 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 304868 471454
rect 303868 471134 304868 471218
rect 303868 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 304868 471134
rect 303868 470866 304868 470898
rect 323868 471454 324868 471486
rect 323868 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 324868 471454
rect 323868 471134 324868 471218
rect 323868 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 324868 471134
rect 323868 470866 324868 470898
rect 343868 471454 344868 471486
rect 343868 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 344868 471454
rect 343868 471134 344868 471218
rect 343868 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 344868 471134
rect 343868 470866 344868 470898
rect 363868 471454 364868 471486
rect 363868 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 364868 471454
rect 363868 471134 364868 471218
rect 363868 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 364868 471134
rect 363868 470866 364868 470898
rect 383868 471454 384868 471486
rect 383868 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 384868 471454
rect 383868 471134 384868 471218
rect 383868 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 384868 471134
rect 383868 470866 384868 470898
rect 403868 471454 404868 471486
rect 403868 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 404868 471454
rect 403868 471134 404868 471218
rect 403868 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 404868 471134
rect 403868 470866 404868 470898
rect 303475 461140 303541 461141
rect 303475 461076 303476 461140
rect 303540 461076 303541 461140
rect 303475 461075 303541 461076
rect 302739 459644 302805 459645
rect 302739 459580 302740 459644
rect 302804 459580 302805 459644
rect 302739 459579 302805 459580
rect 301451 456788 301517 456789
rect 301451 456724 301452 456788
rect 301516 456724 301517 456788
rect 301451 456723 301517 456724
rect 302003 418300 302069 418301
rect 302003 418236 302004 418300
rect 302068 418236 302069 418300
rect 302003 418235 302069 418236
rect 302006 78573 302066 418235
rect 302742 331125 302802 459579
rect 303478 335370 303538 461075
rect 307794 453454 308414 460000
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 416000 308414 416898
rect 312294 457954 312914 460000
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 416000 312914 421398
rect 343794 453454 344414 460000
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 416000 344414 416898
rect 348294 457954 348914 460000
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 416000 348914 421398
rect 379794 453454 380414 460000
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 416000 380414 416898
rect 384294 457954 384914 460000
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 416000 384914 421398
rect 415794 453454 416414 460000
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 416000 416414 416898
rect 313868 403954 314868 403986
rect 313868 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 314868 403954
rect 313868 403634 314868 403718
rect 313868 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 314868 403634
rect 313868 403366 314868 403398
rect 333868 403954 334868 403986
rect 333868 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 334868 403954
rect 333868 403634 334868 403718
rect 333868 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 334868 403634
rect 333868 403366 334868 403398
rect 353868 403954 354868 403986
rect 353868 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 354868 403954
rect 353868 403634 354868 403718
rect 353868 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 354868 403634
rect 353868 403366 354868 403398
rect 373868 403954 374868 403986
rect 373868 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 374868 403954
rect 373868 403634 374868 403718
rect 373868 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 374868 403634
rect 373868 403366 374868 403398
rect 393868 403954 394868 403986
rect 393868 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 394868 403954
rect 393868 403634 394868 403718
rect 393868 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 394868 403634
rect 393868 403366 394868 403398
rect 413868 403954 414868 403986
rect 413868 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 414868 403954
rect 413868 403634 414868 403718
rect 413868 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 414868 403634
rect 413868 403366 414868 403398
rect 303868 399454 304868 399486
rect 303868 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 304868 399454
rect 303868 399134 304868 399218
rect 303868 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 304868 399134
rect 303868 398866 304868 398898
rect 323868 399454 324868 399486
rect 323868 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 324868 399454
rect 323868 399134 324868 399218
rect 323868 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 324868 399134
rect 323868 398866 324868 398898
rect 343868 399454 344868 399486
rect 343868 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 344868 399454
rect 343868 399134 344868 399218
rect 343868 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 344868 399134
rect 343868 398866 344868 398898
rect 363868 399454 364868 399486
rect 363868 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 364868 399454
rect 363868 399134 364868 399218
rect 363868 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 364868 399134
rect 363868 398866 364868 398898
rect 383868 399454 384868 399486
rect 383868 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 384868 399454
rect 383868 399134 384868 399218
rect 383868 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 384868 399134
rect 383868 398866 384868 398898
rect 403868 399454 404868 399486
rect 403868 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 404868 399454
rect 403868 399134 404868 399218
rect 403868 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 404868 399134
rect 403868 398866 404868 398898
rect 313868 367954 314868 367986
rect 313868 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 314868 367954
rect 313868 367634 314868 367718
rect 313868 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 314868 367634
rect 313868 367366 314868 367398
rect 333868 367954 334868 367986
rect 333868 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 334868 367954
rect 333868 367634 334868 367718
rect 333868 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 334868 367634
rect 333868 367366 334868 367398
rect 353868 367954 354868 367986
rect 353868 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 354868 367954
rect 353868 367634 354868 367718
rect 353868 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 354868 367634
rect 353868 367366 354868 367398
rect 373868 367954 374868 367986
rect 373868 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 374868 367954
rect 373868 367634 374868 367718
rect 373868 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 374868 367634
rect 373868 367366 374868 367398
rect 393868 367954 394868 367986
rect 393868 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 394868 367954
rect 393868 367634 394868 367718
rect 393868 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 394868 367634
rect 393868 367366 394868 367398
rect 413868 367954 414868 367986
rect 413868 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 414868 367954
rect 413868 367634 414868 367718
rect 413868 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 414868 367634
rect 413868 367366 414868 367398
rect 303868 363454 304868 363486
rect 303868 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 304868 363454
rect 303868 363134 304868 363218
rect 303868 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 304868 363134
rect 303868 362866 304868 362898
rect 323868 363454 324868 363486
rect 323868 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 324868 363454
rect 323868 363134 324868 363218
rect 323868 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 324868 363134
rect 323868 362866 324868 362898
rect 343868 363454 344868 363486
rect 343868 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 344868 363454
rect 343868 363134 344868 363218
rect 343868 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 344868 363134
rect 343868 362866 344868 362898
rect 363868 363454 364868 363486
rect 363868 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 364868 363454
rect 363868 363134 364868 363218
rect 363868 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 364868 363134
rect 363868 362866 364868 362898
rect 383868 363454 384868 363486
rect 383868 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 384868 363454
rect 383868 363134 384868 363218
rect 383868 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 384868 363134
rect 383868 362866 384868 362898
rect 403868 363454 404868 363486
rect 403868 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 404868 363454
rect 403868 363134 404868 363218
rect 403868 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 404868 363134
rect 403868 362866 404868 362898
rect 302926 335310 303538 335370
rect 302926 332349 302986 335310
rect 302923 332348 302989 332349
rect 302923 332284 302924 332348
rect 302988 332284 302989 332348
rect 302923 332283 302989 332284
rect 302739 331124 302805 331125
rect 302739 331060 302740 331124
rect 302804 331060 302805 331124
rect 302739 331059 302805 331060
rect 302742 158677 302802 331059
rect 302926 203829 302986 332283
rect 325794 327454 326414 332000
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 288000 326414 290898
rect 330294 331954 330914 332000
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 288000 330914 295398
rect 361794 327454 362414 332000
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 288000 362414 290898
rect 366294 331954 366914 332000
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 288000 366914 295398
rect 397794 327454 398414 332000
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 288000 398414 290898
rect 402294 331954 402914 332000
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 288000 402914 295398
rect 313868 259954 314868 259986
rect 313868 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 314868 259954
rect 313868 259634 314868 259718
rect 313868 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 314868 259634
rect 313868 259366 314868 259398
rect 333868 259954 334868 259986
rect 333868 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 334868 259954
rect 333868 259634 334868 259718
rect 333868 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 334868 259634
rect 333868 259366 334868 259398
rect 353868 259954 354868 259986
rect 353868 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 354868 259954
rect 353868 259634 354868 259718
rect 353868 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 354868 259634
rect 353868 259366 354868 259398
rect 373868 259954 374868 259986
rect 373868 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 374868 259954
rect 373868 259634 374868 259718
rect 373868 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 374868 259634
rect 373868 259366 374868 259398
rect 393868 259954 394868 259986
rect 393868 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 394868 259954
rect 393868 259634 394868 259718
rect 393868 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 394868 259634
rect 393868 259366 394868 259398
rect 413868 259954 414868 259986
rect 413868 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 414868 259954
rect 413868 259634 414868 259718
rect 413868 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 414868 259634
rect 413868 259366 414868 259398
rect 303868 255454 304868 255486
rect 303868 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 304868 255454
rect 303868 255134 304868 255218
rect 303868 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 304868 255134
rect 303868 254866 304868 254898
rect 323868 255454 324868 255486
rect 323868 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 324868 255454
rect 323868 255134 324868 255218
rect 323868 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 324868 255134
rect 323868 254866 324868 254898
rect 343868 255454 344868 255486
rect 343868 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 344868 255454
rect 343868 255134 344868 255218
rect 343868 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 344868 255134
rect 343868 254866 344868 254898
rect 363868 255454 364868 255486
rect 363868 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 364868 255454
rect 363868 255134 364868 255218
rect 363868 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 364868 255134
rect 363868 254866 364868 254898
rect 383868 255454 384868 255486
rect 383868 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 384868 255454
rect 383868 255134 384868 255218
rect 383868 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 384868 255134
rect 383868 254866 384868 254898
rect 403868 255454 404868 255486
rect 403868 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 404868 255454
rect 403868 255134 404868 255218
rect 403868 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 404868 255134
rect 403868 254866 404868 254898
rect 313868 223954 314868 223986
rect 313868 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 314868 223954
rect 313868 223634 314868 223718
rect 313868 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 314868 223634
rect 313868 223366 314868 223398
rect 333868 223954 334868 223986
rect 333868 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 334868 223954
rect 333868 223634 334868 223718
rect 333868 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 334868 223634
rect 333868 223366 334868 223398
rect 353868 223954 354868 223986
rect 353868 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 354868 223954
rect 353868 223634 354868 223718
rect 353868 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 354868 223634
rect 353868 223366 354868 223398
rect 373868 223954 374868 223986
rect 373868 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 374868 223954
rect 373868 223634 374868 223718
rect 373868 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 374868 223634
rect 373868 223366 374868 223398
rect 393868 223954 394868 223986
rect 393868 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 394868 223954
rect 393868 223634 394868 223718
rect 393868 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 394868 223634
rect 393868 223366 394868 223398
rect 413868 223954 414868 223986
rect 413868 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 414868 223954
rect 413868 223634 414868 223718
rect 413868 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 414868 223634
rect 413868 223366 414868 223398
rect 303868 219454 304868 219486
rect 303868 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 304868 219454
rect 303868 219134 304868 219218
rect 303868 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 304868 219134
rect 303868 218866 304868 218898
rect 323868 219454 324868 219486
rect 323868 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 324868 219454
rect 323868 219134 324868 219218
rect 323868 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 324868 219134
rect 323868 218866 324868 218898
rect 343868 219454 344868 219486
rect 343868 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 344868 219454
rect 343868 219134 344868 219218
rect 343868 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 344868 219134
rect 343868 218866 344868 218898
rect 363868 219454 364868 219486
rect 363868 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 364868 219454
rect 363868 219134 364868 219218
rect 363868 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 364868 219134
rect 363868 218866 364868 218898
rect 383868 219454 384868 219486
rect 383868 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 384868 219454
rect 383868 219134 384868 219218
rect 383868 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 384868 219134
rect 383868 218866 384868 218898
rect 403868 219454 404868 219486
rect 403868 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 404868 219454
rect 403868 219134 404868 219218
rect 403868 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 404868 219134
rect 403868 218866 404868 218898
rect 302923 203828 302989 203829
rect 302923 203764 302924 203828
rect 302988 203764 302989 203828
rect 302923 203763 302989 203764
rect 302926 200130 302986 203763
rect 302926 200070 303170 200130
rect 302739 158676 302805 158677
rect 302739 158612 302740 158676
rect 302804 158612 302805 158676
rect 302739 158611 302805 158612
rect 302003 78572 302069 78573
rect 302003 78508 302004 78572
rect 302068 78508 302069 78572
rect 302003 78507 302069 78508
rect 299979 77892 300045 77893
rect 299979 77828 299980 77892
rect 300044 77828 300045 77892
rect 299979 77827 300045 77828
rect 302742 60621 302802 158611
rect 303110 76669 303170 200070
rect 303294 196954 303914 204000
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 160000 303914 160398
rect 307794 201454 308414 204000
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 160000 308414 164898
rect 339294 196954 339914 204000
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 160000 339914 160398
rect 343794 201454 344414 204000
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 160000 344414 164898
rect 375294 196954 375914 204000
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 160000 375914 160398
rect 379794 201454 380414 204000
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 160000 380414 164898
rect 411294 196954 411914 204000
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 160000 411914 160398
rect 415794 201454 416414 204000
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 160000 416414 164898
rect 313868 151954 314868 151986
rect 313868 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 314868 151954
rect 313868 151634 314868 151718
rect 313868 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 314868 151634
rect 313868 151366 314868 151398
rect 333868 151954 334868 151986
rect 333868 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 334868 151954
rect 333868 151634 334868 151718
rect 333868 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 334868 151634
rect 333868 151366 334868 151398
rect 353868 151954 354868 151986
rect 353868 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 354868 151954
rect 353868 151634 354868 151718
rect 353868 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 354868 151634
rect 353868 151366 354868 151398
rect 373868 151954 374868 151986
rect 373868 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 374868 151954
rect 373868 151634 374868 151718
rect 373868 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 374868 151634
rect 373868 151366 374868 151398
rect 393868 151954 394868 151986
rect 393868 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 394868 151954
rect 393868 151634 394868 151718
rect 393868 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 394868 151634
rect 393868 151366 394868 151398
rect 413868 151954 414868 151986
rect 413868 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 414868 151954
rect 413868 151634 414868 151718
rect 413868 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 414868 151634
rect 413868 151366 414868 151398
rect 303868 147454 304868 147486
rect 303868 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 304868 147454
rect 303868 147134 304868 147218
rect 303868 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 304868 147134
rect 303868 146866 304868 146898
rect 323868 147454 324868 147486
rect 323868 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 324868 147454
rect 323868 147134 324868 147218
rect 323868 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 324868 147134
rect 323868 146866 324868 146898
rect 343868 147454 344868 147486
rect 343868 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 344868 147454
rect 343868 147134 344868 147218
rect 343868 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 344868 147134
rect 343868 146866 344868 146898
rect 363868 147454 364868 147486
rect 363868 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 364868 147454
rect 363868 147134 364868 147218
rect 363868 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 364868 147134
rect 363868 146866 364868 146898
rect 383868 147454 384868 147486
rect 383868 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 384868 147454
rect 383868 147134 384868 147218
rect 383868 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 384868 147134
rect 383868 146866 384868 146898
rect 403868 147454 404868 147486
rect 403868 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 404868 147454
rect 403868 147134 404868 147218
rect 403868 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 404868 147134
rect 403868 146866 404868 146898
rect 313868 115954 314868 115986
rect 313868 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 314868 115954
rect 313868 115634 314868 115718
rect 313868 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 314868 115634
rect 313868 115366 314868 115398
rect 333868 115954 334868 115986
rect 333868 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 334868 115954
rect 333868 115634 334868 115718
rect 333868 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 334868 115634
rect 333868 115366 334868 115398
rect 353868 115954 354868 115986
rect 353868 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 354868 115954
rect 353868 115634 354868 115718
rect 353868 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 354868 115634
rect 353868 115366 354868 115398
rect 373868 115954 374868 115986
rect 373868 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 374868 115954
rect 373868 115634 374868 115718
rect 373868 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 374868 115634
rect 373868 115366 374868 115398
rect 393868 115954 394868 115986
rect 393868 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 394868 115954
rect 393868 115634 394868 115718
rect 393868 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 394868 115634
rect 393868 115366 394868 115398
rect 413868 115954 414868 115986
rect 413868 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 414868 115954
rect 413868 115634 414868 115718
rect 413868 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 414868 115634
rect 413868 115366 414868 115398
rect 303868 111454 304868 111486
rect 303868 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 304868 111454
rect 303868 111134 304868 111218
rect 303868 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 304868 111134
rect 303868 110866 304868 110898
rect 323868 111454 324868 111486
rect 323868 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 324868 111454
rect 323868 111134 324868 111218
rect 323868 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 324868 111134
rect 323868 110866 324868 110898
rect 343868 111454 344868 111486
rect 343868 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 344868 111454
rect 343868 111134 344868 111218
rect 343868 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 344868 111134
rect 343868 110866 344868 110898
rect 363868 111454 364868 111486
rect 363868 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 364868 111454
rect 363868 111134 364868 111218
rect 363868 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 364868 111134
rect 363868 110866 364868 110898
rect 383868 111454 384868 111486
rect 383868 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 384868 111454
rect 383868 111134 384868 111218
rect 383868 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 384868 111134
rect 383868 110866 384868 110898
rect 403868 111454 404868 111486
rect 403868 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 404868 111454
rect 403868 111134 404868 111218
rect 403868 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 404868 111134
rect 403868 110866 404868 110898
rect 303107 76668 303173 76669
rect 303107 76604 303108 76668
rect 303172 76604 303173 76668
rect 303107 76603 303173 76604
rect 302739 60620 302805 60621
rect 302739 60556 302740 60620
rect 302804 60556 302805 60620
rect 302739 60555 302805 60556
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 213868 43954 214868 43986
rect 213868 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 214868 43954
rect 213868 43634 214868 43718
rect 213868 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 214868 43634
rect 213868 43366 214868 43398
rect 233868 43954 234868 43986
rect 233868 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 234868 43954
rect 233868 43634 234868 43718
rect 233868 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 234868 43634
rect 233868 43366 234868 43398
rect 253868 43954 254868 43986
rect 253868 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 254868 43954
rect 253868 43634 254868 43718
rect 253868 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 254868 43634
rect 253868 43366 254868 43398
rect 273868 43954 274868 43986
rect 273868 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 274868 43954
rect 273868 43634 274868 43718
rect 273868 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 274868 43634
rect 273868 43366 274868 43398
rect 293868 43954 294868 43986
rect 293868 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 294868 43954
rect 293868 43634 294868 43718
rect 293868 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 294868 43634
rect 293868 43366 294868 43398
rect 313868 43954 314868 43986
rect 313868 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 314868 43954
rect 313868 43634 314868 43718
rect 313868 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 314868 43634
rect 313868 43366 314868 43398
rect 333868 43954 334868 43986
rect 333868 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 334868 43954
rect 333868 43634 334868 43718
rect 333868 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 334868 43634
rect 333868 43366 334868 43398
rect 353868 43954 354868 43986
rect 353868 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 354868 43954
rect 353868 43634 354868 43718
rect 353868 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 354868 43634
rect 353868 43366 354868 43398
rect 373868 43954 374868 43986
rect 373868 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 374868 43954
rect 373868 43634 374868 43718
rect 373868 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 374868 43634
rect 373868 43366 374868 43398
rect 393868 43954 394868 43986
rect 393868 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 394868 43954
rect 393868 43634 394868 43718
rect 393868 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 394868 43634
rect 393868 43366 394868 43398
rect 402294 43954 402914 76000
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 203868 39454 204868 39486
rect 203868 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 204868 39454
rect 203868 39134 204868 39218
rect 203868 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 204868 39134
rect 203868 38866 204868 38898
rect 223868 39454 224868 39486
rect 223868 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 224868 39454
rect 223868 39134 224868 39218
rect 223868 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 224868 39134
rect 223868 38866 224868 38898
rect 243868 39454 244868 39486
rect 243868 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 244868 39454
rect 243868 39134 244868 39218
rect 243868 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 244868 39134
rect 243868 38866 244868 38898
rect 263868 39454 264868 39486
rect 263868 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 264868 39454
rect 263868 39134 264868 39218
rect 263868 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 264868 39134
rect 263868 38866 264868 38898
rect 283868 39454 284868 39486
rect 283868 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 284868 39454
rect 283868 39134 284868 39218
rect 283868 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 284868 39134
rect 283868 38866 284868 38898
rect 303868 39454 304868 39486
rect 303868 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 304868 39454
rect 303868 39134 304868 39218
rect 303868 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 304868 39134
rect 303868 38866 304868 38898
rect 323868 39454 324868 39486
rect 323868 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 324868 39454
rect 323868 39134 324868 39218
rect 323868 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 324868 39134
rect 323868 38866 324868 38898
rect 343868 39454 344868 39486
rect 343868 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 344868 39454
rect 343868 39134 344868 39218
rect 343868 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 344868 39134
rect 343868 38866 344868 38898
rect 363868 39454 364868 39486
rect 363868 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 364868 39454
rect 363868 39134 364868 39218
rect 363868 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 364868 39134
rect 363868 38866 364868 38898
rect 383868 39454 384868 39486
rect 383868 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 384868 39454
rect 383868 39134 384868 39218
rect 383868 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 384868 39134
rect 383868 38866 384868 38898
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 22000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 217794 3454 218414 22000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 22000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 22000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 22000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 22000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 253794 3454 254414 22000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 22000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 22000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 22000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 22000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 289794 3454 290414 22000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 22000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 22000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 22000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 22000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 325794 3454 326414 22000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 22000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 22000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 22000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 22000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 361794 3454 362414 22000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 22000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 22000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 22000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 22000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 397794 3454 398414 22000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 48454 407414 76000
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 52954 411914 76000
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 57454 416414 76000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 418110 21997 418170 699755
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 670000 420914 673398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 420131 591292 420197 591293
rect 420131 591228 420132 591292
rect 420196 591228 420197 591292
rect 420131 591227 420197 591228
rect 418659 485076 418725 485077
rect 418659 485012 418660 485076
rect 418724 485012 418725 485076
rect 418659 485011 418725 485012
rect 418662 22133 418722 485011
rect 419579 331396 419645 331397
rect 419579 331332 419580 331396
rect 419644 331332 419645 331396
rect 419579 331331 419645 331332
rect 419582 204373 419642 331331
rect 419579 204372 419645 204373
rect 419579 204308 419580 204372
rect 419644 204308 419645 204372
rect 419579 204307 419645 204308
rect 420134 24173 420194 591227
rect 422339 585852 422405 585853
rect 422339 585788 422340 585852
rect 422404 585788 422405 585852
rect 422339 585787 422405 585788
rect 420294 457954 420914 460000
rect 421051 458284 421117 458285
rect 421051 458220 421052 458284
rect 421116 458220 421117 458284
rect 421051 458219 421117 458220
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 416000 420914 421398
rect 421054 76805 421114 458219
rect 421051 76804 421117 76805
rect 421051 76740 421052 76804
rect 421116 76740 421117 76804
rect 421051 76739 421117 76740
rect 422342 76669 422402 585787
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 422339 76668 422405 76669
rect 422339 76604 422340 76668
rect 422404 76604 422405 76668
rect 422339 76603 422405 76604
rect 420294 61954 420914 76000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420131 24172 420197 24173
rect 420131 24108 420132 24172
rect 420196 24108 420197 24172
rect 420131 24107 420197 24108
rect 418659 22132 418725 22133
rect 418659 22068 418660 22132
rect 418724 22068 418725 22132
rect 418659 22067 418725 22068
rect 418107 21996 418173 21997
rect 418107 21932 418108 21996
rect 418172 21932 418173 21996
rect 418107 21931 418173 21932
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 33930 655718 34166 655954
rect 34250 655718 34486 655954
rect 34570 655718 34806 655954
rect 33930 655398 34166 655634
rect 34250 655398 34486 655634
rect 34570 655398 34806 655634
rect 53930 655718 54166 655954
rect 54250 655718 54486 655954
rect 54570 655718 54806 655954
rect 53930 655398 54166 655634
rect 54250 655398 54486 655634
rect 54570 655398 54806 655634
rect 73930 655718 74166 655954
rect 74250 655718 74486 655954
rect 74570 655718 74806 655954
rect 73930 655398 74166 655634
rect 74250 655398 74486 655634
rect 74570 655398 74806 655634
rect 93930 655718 94166 655954
rect 94250 655718 94486 655954
rect 94570 655718 94806 655954
rect 93930 655398 94166 655634
rect 94250 655398 94486 655634
rect 94570 655398 94806 655634
rect 113930 655718 114166 655954
rect 114250 655718 114486 655954
rect 114570 655718 114806 655954
rect 113930 655398 114166 655634
rect 114250 655398 114486 655634
rect 114570 655398 114806 655634
rect 133930 655718 134166 655954
rect 134250 655718 134486 655954
rect 134570 655718 134806 655954
rect 133930 655398 134166 655634
rect 134250 655398 134486 655634
rect 134570 655398 134806 655634
rect 23930 651218 24166 651454
rect 24250 651218 24486 651454
rect 24570 651218 24806 651454
rect 23930 650898 24166 651134
rect 24250 650898 24486 651134
rect 24570 650898 24806 651134
rect 43930 651218 44166 651454
rect 44250 651218 44486 651454
rect 44570 651218 44806 651454
rect 43930 650898 44166 651134
rect 44250 650898 44486 651134
rect 44570 650898 44806 651134
rect 63930 651218 64166 651454
rect 64250 651218 64486 651454
rect 64570 651218 64806 651454
rect 63930 650898 64166 651134
rect 64250 650898 64486 651134
rect 64570 650898 64806 651134
rect 83930 651218 84166 651454
rect 84250 651218 84486 651454
rect 84570 651218 84806 651454
rect 83930 650898 84166 651134
rect 84250 650898 84486 651134
rect 84570 650898 84806 651134
rect 103930 651218 104166 651454
rect 104250 651218 104486 651454
rect 104570 651218 104806 651454
rect 103930 650898 104166 651134
rect 104250 650898 104486 651134
rect 104570 650898 104806 651134
rect 123930 651218 124166 651454
rect 124250 651218 124486 651454
rect 124570 651218 124806 651454
rect 123930 650898 124166 651134
rect 124250 650898 124486 651134
rect 124570 650898 124806 651134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 33930 619718 34166 619954
rect 34250 619718 34486 619954
rect 34570 619718 34806 619954
rect 33930 619398 34166 619634
rect 34250 619398 34486 619634
rect 34570 619398 34806 619634
rect 53930 619718 54166 619954
rect 54250 619718 54486 619954
rect 54570 619718 54806 619954
rect 53930 619398 54166 619634
rect 54250 619398 54486 619634
rect 54570 619398 54806 619634
rect 73930 619718 74166 619954
rect 74250 619718 74486 619954
rect 74570 619718 74806 619954
rect 73930 619398 74166 619634
rect 74250 619398 74486 619634
rect 74570 619398 74806 619634
rect 93930 619718 94166 619954
rect 94250 619718 94486 619954
rect 94570 619718 94806 619954
rect 93930 619398 94166 619634
rect 94250 619398 94486 619634
rect 94570 619398 94806 619634
rect 113930 619718 114166 619954
rect 114250 619718 114486 619954
rect 114570 619718 114806 619954
rect 113930 619398 114166 619634
rect 114250 619398 114486 619634
rect 114570 619398 114806 619634
rect 133930 619718 134166 619954
rect 134250 619718 134486 619954
rect 134570 619718 134806 619954
rect 133930 619398 134166 619634
rect 134250 619398 134486 619634
rect 134570 619398 134806 619634
rect 23930 615218 24166 615454
rect 24250 615218 24486 615454
rect 24570 615218 24806 615454
rect 23930 614898 24166 615134
rect 24250 614898 24486 615134
rect 24570 614898 24806 615134
rect 43930 615218 44166 615454
rect 44250 615218 44486 615454
rect 44570 615218 44806 615454
rect 43930 614898 44166 615134
rect 44250 614898 44486 615134
rect 44570 614898 44806 615134
rect 63930 615218 64166 615454
rect 64250 615218 64486 615454
rect 64570 615218 64806 615454
rect 63930 614898 64166 615134
rect 64250 614898 64486 615134
rect 64570 614898 64806 615134
rect 83930 615218 84166 615454
rect 84250 615218 84486 615454
rect 84570 615218 84806 615454
rect 83930 614898 84166 615134
rect 84250 614898 84486 615134
rect 84570 614898 84806 615134
rect 103930 615218 104166 615454
rect 104250 615218 104486 615454
rect 104570 615218 104806 615454
rect 103930 614898 104166 615134
rect 104250 614898 104486 615134
rect 104570 614898 104806 615134
rect 123930 615218 124166 615454
rect 124250 615218 124486 615454
rect 124570 615218 124806 615454
rect 123930 614898 124166 615134
rect 124250 614898 124486 615134
rect 124570 614898 124806 615134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 33930 511718 34166 511954
rect 34250 511718 34486 511954
rect 34570 511718 34806 511954
rect 33930 511398 34166 511634
rect 34250 511398 34486 511634
rect 34570 511398 34806 511634
rect 53930 511718 54166 511954
rect 54250 511718 54486 511954
rect 54570 511718 54806 511954
rect 53930 511398 54166 511634
rect 54250 511398 54486 511634
rect 54570 511398 54806 511634
rect 73930 511718 74166 511954
rect 74250 511718 74486 511954
rect 74570 511718 74806 511954
rect 73930 511398 74166 511634
rect 74250 511398 74486 511634
rect 74570 511398 74806 511634
rect 93930 511718 94166 511954
rect 94250 511718 94486 511954
rect 94570 511718 94806 511954
rect 93930 511398 94166 511634
rect 94250 511398 94486 511634
rect 94570 511398 94806 511634
rect 113930 511718 114166 511954
rect 114250 511718 114486 511954
rect 114570 511718 114806 511954
rect 113930 511398 114166 511634
rect 114250 511398 114486 511634
rect 114570 511398 114806 511634
rect 133930 511718 134166 511954
rect 134250 511718 134486 511954
rect 134570 511718 134806 511954
rect 133930 511398 134166 511634
rect 134250 511398 134486 511634
rect 134570 511398 134806 511634
rect 23930 507218 24166 507454
rect 24250 507218 24486 507454
rect 24570 507218 24806 507454
rect 23930 506898 24166 507134
rect 24250 506898 24486 507134
rect 24570 506898 24806 507134
rect 43930 507218 44166 507454
rect 44250 507218 44486 507454
rect 44570 507218 44806 507454
rect 43930 506898 44166 507134
rect 44250 506898 44486 507134
rect 44570 506898 44806 507134
rect 63930 507218 64166 507454
rect 64250 507218 64486 507454
rect 64570 507218 64806 507454
rect 63930 506898 64166 507134
rect 64250 506898 64486 507134
rect 64570 506898 64806 507134
rect 83930 507218 84166 507454
rect 84250 507218 84486 507454
rect 84570 507218 84806 507454
rect 83930 506898 84166 507134
rect 84250 506898 84486 507134
rect 84570 506898 84806 507134
rect 103930 507218 104166 507454
rect 104250 507218 104486 507454
rect 104570 507218 104806 507454
rect 103930 506898 104166 507134
rect 104250 506898 104486 507134
rect 104570 506898 104806 507134
rect 123930 507218 124166 507454
rect 124250 507218 124486 507454
rect 124570 507218 124806 507454
rect 123930 506898 124166 507134
rect 124250 506898 124486 507134
rect 124570 506898 124806 507134
rect 33930 475718 34166 475954
rect 34250 475718 34486 475954
rect 34570 475718 34806 475954
rect 33930 475398 34166 475634
rect 34250 475398 34486 475634
rect 34570 475398 34806 475634
rect 53930 475718 54166 475954
rect 54250 475718 54486 475954
rect 54570 475718 54806 475954
rect 53930 475398 54166 475634
rect 54250 475398 54486 475634
rect 54570 475398 54806 475634
rect 73930 475718 74166 475954
rect 74250 475718 74486 475954
rect 74570 475718 74806 475954
rect 73930 475398 74166 475634
rect 74250 475398 74486 475634
rect 74570 475398 74806 475634
rect 93930 475718 94166 475954
rect 94250 475718 94486 475954
rect 94570 475718 94806 475954
rect 93930 475398 94166 475634
rect 94250 475398 94486 475634
rect 94570 475398 94806 475634
rect 113930 475718 114166 475954
rect 114250 475718 114486 475954
rect 114570 475718 114806 475954
rect 113930 475398 114166 475634
rect 114250 475398 114486 475634
rect 114570 475398 114806 475634
rect 133930 475718 134166 475954
rect 134250 475718 134486 475954
rect 134570 475718 134806 475954
rect 133930 475398 134166 475634
rect 134250 475398 134486 475634
rect 134570 475398 134806 475634
rect 23930 471218 24166 471454
rect 24250 471218 24486 471454
rect 24570 471218 24806 471454
rect 23930 470898 24166 471134
rect 24250 470898 24486 471134
rect 24570 470898 24806 471134
rect 43930 471218 44166 471454
rect 44250 471218 44486 471454
rect 44570 471218 44806 471454
rect 43930 470898 44166 471134
rect 44250 470898 44486 471134
rect 44570 470898 44806 471134
rect 63930 471218 64166 471454
rect 64250 471218 64486 471454
rect 64570 471218 64806 471454
rect 63930 470898 64166 471134
rect 64250 470898 64486 471134
rect 64570 470898 64806 471134
rect 83930 471218 84166 471454
rect 84250 471218 84486 471454
rect 84570 471218 84806 471454
rect 83930 470898 84166 471134
rect 84250 470898 84486 471134
rect 84570 470898 84806 471134
rect 103930 471218 104166 471454
rect 104250 471218 104486 471454
rect 104570 471218 104806 471454
rect 103930 470898 104166 471134
rect 104250 470898 104486 471134
rect 104570 470898 104806 471134
rect 123930 471218 124166 471454
rect 124250 471218 124486 471454
rect 124570 471218 124806 471454
rect 123930 470898 124166 471134
rect 124250 470898 124486 471134
rect 124570 470898 124806 471134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 33930 403718 34166 403954
rect 34250 403718 34486 403954
rect 34570 403718 34806 403954
rect 33930 403398 34166 403634
rect 34250 403398 34486 403634
rect 34570 403398 34806 403634
rect 53930 403718 54166 403954
rect 54250 403718 54486 403954
rect 54570 403718 54806 403954
rect 53930 403398 54166 403634
rect 54250 403398 54486 403634
rect 54570 403398 54806 403634
rect 73930 403718 74166 403954
rect 74250 403718 74486 403954
rect 74570 403718 74806 403954
rect 73930 403398 74166 403634
rect 74250 403398 74486 403634
rect 74570 403398 74806 403634
rect 93930 403718 94166 403954
rect 94250 403718 94486 403954
rect 94570 403718 94806 403954
rect 93930 403398 94166 403634
rect 94250 403398 94486 403634
rect 94570 403398 94806 403634
rect 113930 403718 114166 403954
rect 114250 403718 114486 403954
rect 114570 403718 114806 403954
rect 113930 403398 114166 403634
rect 114250 403398 114486 403634
rect 114570 403398 114806 403634
rect 133930 403718 134166 403954
rect 134250 403718 134486 403954
rect 134570 403718 134806 403954
rect 133930 403398 134166 403634
rect 134250 403398 134486 403634
rect 134570 403398 134806 403634
rect 23930 399218 24166 399454
rect 24250 399218 24486 399454
rect 24570 399218 24806 399454
rect 23930 398898 24166 399134
rect 24250 398898 24486 399134
rect 24570 398898 24806 399134
rect 43930 399218 44166 399454
rect 44250 399218 44486 399454
rect 44570 399218 44806 399454
rect 43930 398898 44166 399134
rect 44250 398898 44486 399134
rect 44570 398898 44806 399134
rect 63930 399218 64166 399454
rect 64250 399218 64486 399454
rect 64570 399218 64806 399454
rect 63930 398898 64166 399134
rect 64250 398898 64486 399134
rect 64570 398898 64806 399134
rect 83930 399218 84166 399454
rect 84250 399218 84486 399454
rect 84570 399218 84806 399454
rect 83930 398898 84166 399134
rect 84250 398898 84486 399134
rect 84570 398898 84806 399134
rect 103930 399218 104166 399454
rect 104250 399218 104486 399454
rect 104570 399218 104806 399454
rect 103930 398898 104166 399134
rect 104250 398898 104486 399134
rect 104570 398898 104806 399134
rect 123930 399218 124166 399454
rect 124250 399218 124486 399454
rect 124570 399218 124806 399454
rect 123930 398898 124166 399134
rect 124250 398898 124486 399134
rect 124570 398898 124806 399134
rect 33930 367718 34166 367954
rect 34250 367718 34486 367954
rect 34570 367718 34806 367954
rect 33930 367398 34166 367634
rect 34250 367398 34486 367634
rect 34570 367398 34806 367634
rect 53930 367718 54166 367954
rect 54250 367718 54486 367954
rect 54570 367718 54806 367954
rect 53930 367398 54166 367634
rect 54250 367398 54486 367634
rect 54570 367398 54806 367634
rect 73930 367718 74166 367954
rect 74250 367718 74486 367954
rect 74570 367718 74806 367954
rect 73930 367398 74166 367634
rect 74250 367398 74486 367634
rect 74570 367398 74806 367634
rect 93930 367718 94166 367954
rect 94250 367718 94486 367954
rect 94570 367718 94806 367954
rect 93930 367398 94166 367634
rect 94250 367398 94486 367634
rect 94570 367398 94806 367634
rect 113930 367718 114166 367954
rect 114250 367718 114486 367954
rect 114570 367718 114806 367954
rect 113930 367398 114166 367634
rect 114250 367398 114486 367634
rect 114570 367398 114806 367634
rect 133930 367718 134166 367954
rect 134250 367718 134486 367954
rect 134570 367718 134806 367954
rect 133930 367398 134166 367634
rect 134250 367398 134486 367634
rect 134570 367398 134806 367634
rect 23930 363218 24166 363454
rect 24250 363218 24486 363454
rect 24570 363218 24806 363454
rect 23930 362898 24166 363134
rect 24250 362898 24486 363134
rect 24570 362898 24806 363134
rect 43930 363218 44166 363454
rect 44250 363218 44486 363454
rect 44570 363218 44806 363454
rect 43930 362898 44166 363134
rect 44250 362898 44486 363134
rect 44570 362898 44806 363134
rect 63930 363218 64166 363454
rect 64250 363218 64486 363454
rect 64570 363218 64806 363454
rect 63930 362898 64166 363134
rect 64250 362898 64486 363134
rect 64570 362898 64806 363134
rect 83930 363218 84166 363454
rect 84250 363218 84486 363454
rect 84570 363218 84806 363454
rect 83930 362898 84166 363134
rect 84250 362898 84486 363134
rect 84570 362898 84806 363134
rect 103930 363218 104166 363454
rect 104250 363218 104486 363454
rect 104570 363218 104806 363454
rect 103930 362898 104166 363134
rect 104250 362898 104486 363134
rect 104570 362898 104806 363134
rect 123930 363218 124166 363454
rect 124250 363218 124486 363454
rect 124570 363218 124806 363454
rect 123930 362898 124166 363134
rect 124250 362898 124486 363134
rect 124570 362898 124806 363134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 33930 259718 34166 259954
rect 34250 259718 34486 259954
rect 34570 259718 34806 259954
rect 33930 259398 34166 259634
rect 34250 259398 34486 259634
rect 34570 259398 34806 259634
rect 53930 259718 54166 259954
rect 54250 259718 54486 259954
rect 54570 259718 54806 259954
rect 53930 259398 54166 259634
rect 54250 259398 54486 259634
rect 54570 259398 54806 259634
rect 73930 259718 74166 259954
rect 74250 259718 74486 259954
rect 74570 259718 74806 259954
rect 73930 259398 74166 259634
rect 74250 259398 74486 259634
rect 74570 259398 74806 259634
rect 93930 259718 94166 259954
rect 94250 259718 94486 259954
rect 94570 259718 94806 259954
rect 93930 259398 94166 259634
rect 94250 259398 94486 259634
rect 94570 259398 94806 259634
rect 113930 259718 114166 259954
rect 114250 259718 114486 259954
rect 114570 259718 114806 259954
rect 113930 259398 114166 259634
rect 114250 259398 114486 259634
rect 114570 259398 114806 259634
rect 133930 259718 134166 259954
rect 134250 259718 134486 259954
rect 134570 259718 134806 259954
rect 133930 259398 134166 259634
rect 134250 259398 134486 259634
rect 134570 259398 134806 259634
rect 23930 255218 24166 255454
rect 24250 255218 24486 255454
rect 24570 255218 24806 255454
rect 23930 254898 24166 255134
rect 24250 254898 24486 255134
rect 24570 254898 24806 255134
rect 43930 255218 44166 255454
rect 44250 255218 44486 255454
rect 44570 255218 44806 255454
rect 43930 254898 44166 255134
rect 44250 254898 44486 255134
rect 44570 254898 44806 255134
rect 63930 255218 64166 255454
rect 64250 255218 64486 255454
rect 64570 255218 64806 255454
rect 63930 254898 64166 255134
rect 64250 254898 64486 255134
rect 64570 254898 64806 255134
rect 83930 255218 84166 255454
rect 84250 255218 84486 255454
rect 84570 255218 84806 255454
rect 83930 254898 84166 255134
rect 84250 254898 84486 255134
rect 84570 254898 84806 255134
rect 103930 255218 104166 255454
rect 104250 255218 104486 255454
rect 104570 255218 104806 255454
rect 103930 254898 104166 255134
rect 104250 254898 104486 255134
rect 104570 254898 104806 255134
rect 123930 255218 124166 255454
rect 124250 255218 124486 255454
rect 124570 255218 124806 255454
rect 123930 254898 124166 255134
rect 124250 254898 124486 255134
rect 124570 254898 124806 255134
rect 33930 223718 34166 223954
rect 34250 223718 34486 223954
rect 34570 223718 34806 223954
rect 33930 223398 34166 223634
rect 34250 223398 34486 223634
rect 34570 223398 34806 223634
rect 53930 223718 54166 223954
rect 54250 223718 54486 223954
rect 54570 223718 54806 223954
rect 53930 223398 54166 223634
rect 54250 223398 54486 223634
rect 54570 223398 54806 223634
rect 73930 223718 74166 223954
rect 74250 223718 74486 223954
rect 74570 223718 74806 223954
rect 73930 223398 74166 223634
rect 74250 223398 74486 223634
rect 74570 223398 74806 223634
rect 93930 223718 94166 223954
rect 94250 223718 94486 223954
rect 94570 223718 94806 223954
rect 93930 223398 94166 223634
rect 94250 223398 94486 223634
rect 94570 223398 94806 223634
rect 113930 223718 114166 223954
rect 114250 223718 114486 223954
rect 114570 223718 114806 223954
rect 113930 223398 114166 223634
rect 114250 223398 114486 223634
rect 114570 223398 114806 223634
rect 133930 223718 134166 223954
rect 134250 223718 134486 223954
rect 134570 223718 134806 223954
rect 133930 223398 134166 223634
rect 134250 223398 134486 223634
rect 134570 223398 134806 223634
rect 23930 219218 24166 219454
rect 24250 219218 24486 219454
rect 24570 219218 24806 219454
rect 23930 218898 24166 219134
rect 24250 218898 24486 219134
rect 24570 218898 24806 219134
rect 43930 219218 44166 219454
rect 44250 219218 44486 219454
rect 44570 219218 44806 219454
rect 43930 218898 44166 219134
rect 44250 218898 44486 219134
rect 44570 218898 44806 219134
rect 63930 219218 64166 219454
rect 64250 219218 64486 219454
rect 64570 219218 64806 219454
rect 63930 218898 64166 219134
rect 64250 218898 64486 219134
rect 64570 218898 64806 219134
rect 83930 219218 84166 219454
rect 84250 219218 84486 219454
rect 84570 219218 84806 219454
rect 83930 218898 84166 219134
rect 84250 218898 84486 219134
rect 84570 218898 84806 219134
rect 103930 219218 104166 219454
rect 104250 219218 104486 219454
rect 104570 219218 104806 219454
rect 103930 218898 104166 219134
rect 104250 218898 104486 219134
rect 104570 218898 104806 219134
rect 123930 219218 124166 219454
rect 124250 219218 124486 219454
rect 124570 219218 124806 219454
rect 123930 218898 124166 219134
rect 124250 218898 124486 219134
rect 124570 218898 124806 219134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 33930 151718 34166 151954
rect 34250 151718 34486 151954
rect 34570 151718 34806 151954
rect 33930 151398 34166 151634
rect 34250 151398 34486 151634
rect 34570 151398 34806 151634
rect 53930 151718 54166 151954
rect 54250 151718 54486 151954
rect 54570 151718 54806 151954
rect 53930 151398 54166 151634
rect 54250 151398 54486 151634
rect 54570 151398 54806 151634
rect 73930 151718 74166 151954
rect 74250 151718 74486 151954
rect 74570 151718 74806 151954
rect 73930 151398 74166 151634
rect 74250 151398 74486 151634
rect 74570 151398 74806 151634
rect 93930 151718 94166 151954
rect 94250 151718 94486 151954
rect 94570 151718 94806 151954
rect 93930 151398 94166 151634
rect 94250 151398 94486 151634
rect 94570 151398 94806 151634
rect 113930 151718 114166 151954
rect 114250 151718 114486 151954
rect 114570 151718 114806 151954
rect 113930 151398 114166 151634
rect 114250 151398 114486 151634
rect 114570 151398 114806 151634
rect 133930 151718 134166 151954
rect 134250 151718 134486 151954
rect 134570 151718 134806 151954
rect 133930 151398 134166 151634
rect 134250 151398 134486 151634
rect 134570 151398 134806 151634
rect 23930 147218 24166 147454
rect 24250 147218 24486 147454
rect 24570 147218 24806 147454
rect 23930 146898 24166 147134
rect 24250 146898 24486 147134
rect 24570 146898 24806 147134
rect 43930 147218 44166 147454
rect 44250 147218 44486 147454
rect 44570 147218 44806 147454
rect 43930 146898 44166 147134
rect 44250 146898 44486 147134
rect 44570 146898 44806 147134
rect 63930 147218 64166 147454
rect 64250 147218 64486 147454
rect 64570 147218 64806 147454
rect 63930 146898 64166 147134
rect 64250 146898 64486 147134
rect 64570 146898 64806 147134
rect 83930 147218 84166 147454
rect 84250 147218 84486 147454
rect 84570 147218 84806 147454
rect 83930 146898 84166 147134
rect 84250 146898 84486 147134
rect 84570 146898 84806 147134
rect 103930 147218 104166 147454
rect 104250 147218 104486 147454
rect 104570 147218 104806 147454
rect 103930 146898 104166 147134
rect 104250 146898 104486 147134
rect 104570 146898 104806 147134
rect 123930 147218 124166 147454
rect 124250 147218 124486 147454
rect 124570 147218 124806 147454
rect 123930 146898 124166 147134
rect 124250 146898 124486 147134
rect 124570 146898 124806 147134
rect 33930 115718 34166 115954
rect 34250 115718 34486 115954
rect 34570 115718 34806 115954
rect 33930 115398 34166 115634
rect 34250 115398 34486 115634
rect 34570 115398 34806 115634
rect 53930 115718 54166 115954
rect 54250 115718 54486 115954
rect 54570 115718 54806 115954
rect 53930 115398 54166 115634
rect 54250 115398 54486 115634
rect 54570 115398 54806 115634
rect 73930 115718 74166 115954
rect 74250 115718 74486 115954
rect 74570 115718 74806 115954
rect 73930 115398 74166 115634
rect 74250 115398 74486 115634
rect 74570 115398 74806 115634
rect 93930 115718 94166 115954
rect 94250 115718 94486 115954
rect 94570 115718 94806 115954
rect 93930 115398 94166 115634
rect 94250 115398 94486 115634
rect 94570 115398 94806 115634
rect 113930 115718 114166 115954
rect 114250 115718 114486 115954
rect 114570 115718 114806 115954
rect 113930 115398 114166 115634
rect 114250 115398 114486 115634
rect 114570 115398 114806 115634
rect 133930 115718 134166 115954
rect 134250 115718 134486 115954
rect 134570 115718 134806 115954
rect 133930 115398 134166 115634
rect 134250 115398 134486 115634
rect 134570 115398 134806 115634
rect 23930 111218 24166 111454
rect 24250 111218 24486 111454
rect 24570 111218 24806 111454
rect 23930 110898 24166 111134
rect 24250 110898 24486 111134
rect 24570 110898 24806 111134
rect 43930 111218 44166 111454
rect 44250 111218 44486 111454
rect 44570 111218 44806 111454
rect 43930 110898 44166 111134
rect 44250 110898 44486 111134
rect 44570 110898 44806 111134
rect 63930 111218 64166 111454
rect 64250 111218 64486 111454
rect 64570 111218 64806 111454
rect 63930 110898 64166 111134
rect 64250 110898 64486 111134
rect 64570 110898 64806 111134
rect 83930 111218 84166 111454
rect 84250 111218 84486 111454
rect 84570 111218 84806 111454
rect 83930 110898 84166 111134
rect 84250 110898 84486 111134
rect 84570 110898 84806 111134
rect 103930 111218 104166 111454
rect 104250 111218 104486 111454
rect 104570 111218 104806 111454
rect 103930 110898 104166 111134
rect 104250 110898 104486 111134
rect 104570 110898 104806 111134
rect 123930 111218 124166 111454
rect 124250 111218 124486 111454
rect 124570 111218 124806 111454
rect 123930 110898 124166 111134
rect 124250 110898 124486 111134
rect 124570 110898 124806 111134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 79610 43718 79846 43954
rect 79610 43398 79846 43634
rect 64250 39218 64486 39454
rect 64250 38898 64486 39134
rect 94970 39218 95206 39454
rect 94970 38898 95206 39134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 313930 655718 314166 655954
rect 314250 655718 314486 655954
rect 314570 655718 314806 655954
rect 313930 655398 314166 655634
rect 314250 655398 314486 655634
rect 314570 655398 314806 655634
rect 333930 655718 334166 655954
rect 334250 655718 334486 655954
rect 334570 655718 334806 655954
rect 333930 655398 334166 655634
rect 334250 655398 334486 655634
rect 334570 655398 334806 655634
rect 353930 655718 354166 655954
rect 354250 655718 354486 655954
rect 354570 655718 354806 655954
rect 353930 655398 354166 655634
rect 354250 655398 354486 655634
rect 354570 655398 354806 655634
rect 373930 655718 374166 655954
rect 374250 655718 374486 655954
rect 374570 655718 374806 655954
rect 373930 655398 374166 655634
rect 374250 655398 374486 655634
rect 374570 655398 374806 655634
rect 393930 655718 394166 655954
rect 394250 655718 394486 655954
rect 394570 655718 394806 655954
rect 393930 655398 394166 655634
rect 394250 655398 394486 655634
rect 394570 655398 394806 655634
rect 413930 655718 414166 655954
rect 414250 655718 414486 655954
rect 414570 655718 414806 655954
rect 413930 655398 414166 655634
rect 414250 655398 414486 655634
rect 414570 655398 414806 655634
rect 303930 651218 304166 651454
rect 304250 651218 304486 651454
rect 304570 651218 304806 651454
rect 303930 650898 304166 651134
rect 304250 650898 304486 651134
rect 304570 650898 304806 651134
rect 323930 651218 324166 651454
rect 324250 651218 324486 651454
rect 324570 651218 324806 651454
rect 323930 650898 324166 651134
rect 324250 650898 324486 651134
rect 324570 650898 324806 651134
rect 343930 651218 344166 651454
rect 344250 651218 344486 651454
rect 344570 651218 344806 651454
rect 343930 650898 344166 651134
rect 344250 650898 344486 651134
rect 344570 650898 344806 651134
rect 363930 651218 364166 651454
rect 364250 651218 364486 651454
rect 364570 651218 364806 651454
rect 363930 650898 364166 651134
rect 364250 650898 364486 651134
rect 364570 650898 364806 651134
rect 383930 651218 384166 651454
rect 384250 651218 384486 651454
rect 384570 651218 384806 651454
rect 383930 650898 384166 651134
rect 384250 650898 384486 651134
rect 384570 650898 384806 651134
rect 403930 651218 404166 651454
rect 404250 651218 404486 651454
rect 404570 651218 404806 651454
rect 403930 650898 404166 651134
rect 404250 650898 404486 651134
rect 404570 650898 404806 651134
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 313930 619718 314166 619954
rect 314250 619718 314486 619954
rect 314570 619718 314806 619954
rect 313930 619398 314166 619634
rect 314250 619398 314486 619634
rect 314570 619398 314806 619634
rect 333930 619718 334166 619954
rect 334250 619718 334486 619954
rect 334570 619718 334806 619954
rect 333930 619398 334166 619634
rect 334250 619398 334486 619634
rect 334570 619398 334806 619634
rect 353930 619718 354166 619954
rect 354250 619718 354486 619954
rect 354570 619718 354806 619954
rect 353930 619398 354166 619634
rect 354250 619398 354486 619634
rect 354570 619398 354806 619634
rect 373930 619718 374166 619954
rect 374250 619718 374486 619954
rect 374570 619718 374806 619954
rect 373930 619398 374166 619634
rect 374250 619398 374486 619634
rect 374570 619398 374806 619634
rect 393930 619718 394166 619954
rect 394250 619718 394486 619954
rect 394570 619718 394806 619954
rect 393930 619398 394166 619634
rect 394250 619398 394486 619634
rect 394570 619398 394806 619634
rect 413930 619718 414166 619954
rect 414250 619718 414486 619954
rect 414570 619718 414806 619954
rect 413930 619398 414166 619634
rect 414250 619398 414486 619634
rect 414570 619398 414806 619634
rect 303930 615218 304166 615454
rect 304250 615218 304486 615454
rect 304570 615218 304806 615454
rect 303930 614898 304166 615134
rect 304250 614898 304486 615134
rect 304570 614898 304806 615134
rect 323930 615218 324166 615454
rect 324250 615218 324486 615454
rect 324570 615218 324806 615454
rect 323930 614898 324166 615134
rect 324250 614898 324486 615134
rect 324570 614898 324806 615134
rect 343930 615218 344166 615454
rect 344250 615218 344486 615454
rect 344570 615218 344806 615454
rect 343930 614898 344166 615134
rect 344250 614898 344486 615134
rect 344570 614898 344806 615134
rect 363930 615218 364166 615454
rect 364250 615218 364486 615454
rect 364570 615218 364806 615454
rect 363930 614898 364166 615134
rect 364250 614898 364486 615134
rect 364570 614898 364806 615134
rect 383930 615218 384166 615454
rect 384250 615218 384486 615454
rect 384570 615218 384806 615454
rect 383930 614898 384166 615134
rect 384250 614898 384486 615134
rect 384570 614898 384806 615134
rect 403930 615218 404166 615454
rect 404250 615218 404486 615454
rect 404570 615218 404806 615454
rect 403930 614898 404166 615134
rect 404250 614898 404486 615134
rect 404570 614898 404806 615134
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 313930 511718 314166 511954
rect 314250 511718 314486 511954
rect 314570 511718 314806 511954
rect 313930 511398 314166 511634
rect 314250 511398 314486 511634
rect 314570 511398 314806 511634
rect 333930 511718 334166 511954
rect 334250 511718 334486 511954
rect 334570 511718 334806 511954
rect 333930 511398 334166 511634
rect 334250 511398 334486 511634
rect 334570 511398 334806 511634
rect 353930 511718 354166 511954
rect 354250 511718 354486 511954
rect 354570 511718 354806 511954
rect 353930 511398 354166 511634
rect 354250 511398 354486 511634
rect 354570 511398 354806 511634
rect 373930 511718 374166 511954
rect 374250 511718 374486 511954
rect 374570 511718 374806 511954
rect 373930 511398 374166 511634
rect 374250 511398 374486 511634
rect 374570 511398 374806 511634
rect 393930 511718 394166 511954
rect 394250 511718 394486 511954
rect 394570 511718 394806 511954
rect 393930 511398 394166 511634
rect 394250 511398 394486 511634
rect 394570 511398 394806 511634
rect 413930 511718 414166 511954
rect 414250 511718 414486 511954
rect 414570 511718 414806 511954
rect 413930 511398 414166 511634
rect 414250 511398 414486 511634
rect 414570 511398 414806 511634
rect 303930 507218 304166 507454
rect 304250 507218 304486 507454
rect 304570 507218 304806 507454
rect 303930 506898 304166 507134
rect 304250 506898 304486 507134
rect 304570 506898 304806 507134
rect 323930 507218 324166 507454
rect 324250 507218 324486 507454
rect 324570 507218 324806 507454
rect 323930 506898 324166 507134
rect 324250 506898 324486 507134
rect 324570 506898 324806 507134
rect 343930 507218 344166 507454
rect 344250 507218 344486 507454
rect 344570 507218 344806 507454
rect 343930 506898 344166 507134
rect 344250 506898 344486 507134
rect 344570 506898 344806 507134
rect 363930 507218 364166 507454
rect 364250 507218 364486 507454
rect 364570 507218 364806 507454
rect 363930 506898 364166 507134
rect 364250 506898 364486 507134
rect 364570 506898 364806 507134
rect 383930 507218 384166 507454
rect 384250 507218 384486 507454
rect 384570 507218 384806 507454
rect 383930 506898 384166 507134
rect 384250 506898 384486 507134
rect 384570 506898 384806 507134
rect 403930 507218 404166 507454
rect 404250 507218 404486 507454
rect 404570 507218 404806 507454
rect 403930 506898 404166 507134
rect 404250 506898 404486 507134
rect 404570 506898 404806 507134
rect 313930 475718 314166 475954
rect 314250 475718 314486 475954
rect 314570 475718 314806 475954
rect 313930 475398 314166 475634
rect 314250 475398 314486 475634
rect 314570 475398 314806 475634
rect 333930 475718 334166 475954
rect 334250 475718 334486 475954
rect 334570 475718 334806 475954
rect 333930 475398 334166 475634
rect 334250 475398 334486 475634
rect 334570 475398 334806 475634
rect 353930 475718 354166 475954
rect 354250 475718 354486 475954
rect 354570 475718 354806 475954
rect 353930 475398 354166 475634
rect 354250 475398 354486 475634
rect 354570 475398 354806 475634
rect 373930 475718 374166 475954
rect 374250 475718 374486 475954
rect 374570 475718 374806 475954
rect 373930 475398 374166 475634
rect 374250 475398 374486 475634
rect 374570 475398 374806 475634
rect 393930 475718 394166 475954
rect 394250 475718 394486 475954
rect 394570 475718 394806 475954
rect 393930 475398 394166 475634
rect 394250 475398 394486 475634
rect 394570 475398 394806 475634
rect 413930 475718 414166 475954
rect 414250 475718 414486 475954
rect 414570 475718 414806 475954
rect 413930 475398 414166 475634
rect 414250 475398 414486 475634
rect 414570 475398 414806 475634
rect 303930 471218 304166 471454
rect 304250 471218 304486 471454
rect 304570 471218 304806 471454
rect 303930 470898 304166 471134
rect 304250 470898 304486 471134
rect 304570 470898 304806 471134
rect 323930 471218 324166 471454
rect 324250 471218 324486 471454
rect 324570 471218 324806 471454
rect 323930 470898 324166 471134
rect 324250 470898 324486 471134
rect 324570 470898 324806 471134
rect 343930 471218 344166 471454
rect 344250 471218 344486 471454
rect 344570 471218 344806 471454
rect 343930 470898 344166 471134
rect 344250 470898 344486 471134
rect 344570 470898 344806 471134
rect 363930 471218 364166 471454
rect 364250 471218 364486 471454
rect 364570 471218 364806 471454
rect 363930 470898 364166 471134
rect 364250 470898 364486 471134
rect 364570 470898 364806 471134
rect 383930 471218 384166 471454
rect 384250 471218 384486 471454
rect 384570 471218 384806 471454
rect 383930 470898 384166 471134
rect 384250 470898 384486 471134
rect 384570 470898 384806 471134
rect 403930 471218 404166 471454
rect 404250 471218 404486 471454
rect 404570 471218 404806 471454
rect 403930 470898 404166 471134
rect 404250 470898 404486 471134
rect 404570 470898 404806 471134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 313930 403718 314166 403954
rect 314250 403718 314486 403954
rect 314570 403718 314806 403954
rect 313930 403398 314166 403634
rect 314250 403398 314486 403634
rect 314570 403398 314806 403634
rect 333930 403718 334166 403954
rect 334250 403718 334486 403954
rect 334570 403718 334806 403954
rect 333930 403398 334166 403634
rect 334250 403398 334486 403634
rect 334570 403398 334806 403634
rect 353930 403718 354166 403954
rect 354250 403718 354486 403954
rect 354570 403718 354806 403954
rect 353930 403398 354166 403634
rect 354250 403398 354486 403634
rect 354570 403398 354806 403634
rect 373930 403718 374166 403954
rect 374250 403718 374486 403954
rect 374570 403718 374806 403954
rect 373930 403398 374166 403634
rect 374250 403398 374486 403634
rect 374570 403398 374806 403634
rect 393930 403718 394166 403954
rect 394250 403718 394486 403954
rect 394570 403718 394806 403954
rect 393930 403398 394166 403634
rect 394250 403398 394486 403634
rect 394570 403398 394806 403634
rect 413930 403718 414166 403954
rect 414250 403718 414486 403954
rect 414570 403718 414806 403954
rect 413930 403398 414166 403634
rect 414250 403398 414486 403634
rect 414570 403398 414806 403634
rect 303930 399218 304166 399454
rect 304250 399218 304486 399454
rect 304570 399218 304806 399454
rect 303930 398898 304166 399134
rect 304250 398898 304486 399134
rect 304570 398898 304806 399134
rect 323930 399218 324166 399454
rect 324250 399218 324486 399454
rect 324570 399218 324806 399454
rect 323930 398898 324166 399134
rect 324250 398898 324486 399134
rect 324570 398898 324806 399134
rect 343930 399218 344166 399454
rect 344250 399218 344486 399454
rect 344570 399218 344806 399454
rect 343930 398898 344166 399134
rect 344250 398898 344486 399134
rect 344570 398898 344806 399134
rect 363930 399218 364166 399454
rect 364250 399218 364486 399454
rect 364570 399218 364806 399454
rect 363930 398898 364166 399134
rect 364250 398898 364486 399134
rect 364570 398898 364806 399134
rect 383930 399218 384166 399454
rect 384250 399218 384486 399454
rect 384570 399218 384806 399454
rect 383930 398898 384166 399134
rect 384250 398898 384486 399134
rect 384570 398898 384806 399134
rect 403930 399218 404166 399454
rect 404250 399218 404486 399454
rect 404570 399218 404806 399454
rect 403930 398898 404166 399134
rect 404250 398898 404486 399134
rect 404570 398898 404806 399134
rect 313930 367718 314166 367954
rect 314250 367718 314486 367954
rect 314570 367718 314806 367954
rect 313930 367398 314166 367634
rect 314250 367398 314486 367634
rect 314570 367398 314806 367634
rect 333930 367718 334166 367954
rect 334250 367718 334486 367954
rect 334570 367718 334806 367954
rect 333930 367398 334166 367634
rect 334250 367398 334486 367634
rect 334570 367398 334806 367634
rect 353930 367718 354166 367954
rect 354250 367718 354486 367954
rect 354570 367718 354806 367954
rect 353930 367398 354166 367634
rect 354250 367398 354486 367634
rect 354570 367398 354806 367634
rect 373930 367718 374166 367954
rect 374250 367718 374486 367954
rect 374570 367718 374806 367954
rect 373930 367398 374166 367634
rect 374250 367398 374486 367634
rect 374570 367398 374806 367634
rect 393930 367718 394166 367954
rect 394250 367718 394486 367954
rect 394570 367718 394806 367954
rect 393930 367398 394166 367634
rect 394250 367398 394486 367634
rect 394570 367398 394806 367634
rect 413930 367718 414166 367954
rect 414250 367718 414486 367954
rect 414570 367718 414806 367954
rect 413930 367398 414166 367634
rect 414250 367398 414486 367634
rect 414570 367398 414806 367634
rect 303930 363218 304166 363454
rect 304250 363218 304486 363454
rect 304570 363218 304806 363454
rect 303930 362898 304166 363134
rect 304250 362898 304486 363134
rect 304570 362898 304806 363134
rect 323930 363218 324166 363454
rect 324250 363218 324486 363454
rect 324570 363218 324806 363454
rect 323930 362898 324166 363134
rect 324250 362898 324486 363134
rect 324570 362898 324806 363134
rect 343930 363218 344166 363454
rect 344250 363218 344486 363454
rect 344570 363218 344806 363454
rect 343930 362898 344166 363134
rect 344250 362898 344486 363134
rect 344570 362898 344806 363134
rect 363930 363218 364166 363454
rect 364250 363218 364486 363454
rect 364570 363218 364806 363454
rect 363930 362898 364166 363134
rect 364250 362898 364486 363134
rect 364570 362898 364806 363134
rect 383930 363218 384166 363454
rect 384250 363218 384486 363454
rect 384570 363218 384806 363454
rect 383930 362898 384166 363134
rect 384250 362898 384486 363134
rect 384570 362898 384806 363134
rect 403930 363218 404166 363454
rect 404250 363218 404486 363454
rect 404570 363218 404806 363454
rect 403930 362898 404166 363134
rect 404250 362898 404486 363134
rect 404570 362898 404806 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 313930 259718 314166 259954
rect 314250 259718 314486 259954
rect 314570 259718 314806 259954
rect 313930 259398 314166 259634
rect 314250 259398 314486 259634
rect 314570 259398 314806 259634
rect 333930 259718 334166 259954
rect 334250 259718 334486 259954
rect 334570 259718 334806 259954
rect 333930 259398 334166 259634
rect 334250 259398 334486 259634
rect 334570 259398 334806 259634
rect 353930 259718 354166 259954
rect 354250 259718 354486 259954
rect 354570 259718 354806 259954
rect 353930 259398 354166 259634
rect 354250 259398 354486 259634
rect 354570 259398 354806 259634
rect 373930 259718 374166 259954
rect 374250 259718 374486 259954
rect 374570 259718 374806 259954
rect 373930 259398 374166 259634
rect 374250 259398 374486 259634
rect 374570 259398 374806 259634
rect 393930 259718 394166 259954
rect 394250 259718 394486 259954
rect 394570 259718 394806 259954
rect 393930 259398 394166 259634
rect 394250 259398 394486 259634
rect 394570 259398 394806 259634
rect 413930 259718 414166 259954
rect 414250 259718 414486 259954
rect 414570 259718 414806 259954
rect 413930 259398 414166 259634
rect 414250 259398 414486 259634
rect 414570 259398 414806 259634
rect 303930 255218 304166 255454
rect 304250 255218 304486 255454
rect 304570 255218 304806 255454
rect 303930 254898 304166 255134
rect 304250 254898 304486 255134
rect 304570 254898 304806 255134
rect 323930 255218 324166 255454
rect 324250 255218 324486 255454
rect 324570 255218 324806 255454
rect 323930 254898 324166 255134
rect 324250 254898 324486 255134
rect 324570 254898 324806 255134
rect 343930 255218 344166 255454
rect 344250 255218 344486 255454
rect 344570 255218 344806 255454
rect 343930 254898 344166 255134
rect 344250 254898 344486 255134
rect 344570 254898 344806 255134
rect 363930 255218 364166 255454
rect 364250 255218 364486 255454
rect 364570 255218 364806 255454
rect 363930 254898 364166 255134
rect 364250 254898 364486 255134
rect 364570 254898 364806 255134
rect 383930 255218 384166 255454
rect 384250 255218 384486 255454
rect 384570 255218 384806 255454
rect 383930 254898 384166 255134
rect 384250 254898 384486 255134
rect 384570 254898 384806 255134
rect 403930 255218 404166 255454
rect 404250 255218 404486 255454
rect 404570 255218 404806 255454
rect 403930 254898 404166 255134
rect 404250 254898 404486 255134
rect 404570 254898 404806 255134
rect 313930 223718 314166 223954
rect 314250 223718 314486 223954
rect 314570 223718 314806 223954
rect 313930 223398 314166 223634
rect 314250 223398 314486 223634
rect 314570 223398 314806 223634
rect 333930 223718 334166 223954
rect 334250 223718 334486 223954
rect 334570 223718 334806 223954
rect 333930 223398 334166 223634
rect 334250 223398 334486 223634
rect 334570 223398 334806 223634
rect 353930 223718 354166 223954
rect 354250 223718 354486 223954
rect 354570 223718 354806 223954
rect 353930 223398 354166 223634
rect 354250 223398 354486 223634
rect 354570 223398 354806 223634
rect 373930 223718 374166 223954
rect 374250 223718 374486 223954
rect 374570 223718 374806 223954
rect 373930 223398 374166 223634
rect 374250 223398 374486 223634
rect 374570 223398 374806 223634
rect 393930 223718 394166 223954
rect 394250 223718 394486 223954
rect 394570 223718 394806 223954
rect 393930 223398 394166 223634
rect 394250 223398 394486 223634
rect 394570 223398 394806 223634
rect 413930 223718 414166 223954
rect 414250 223718 414486 223954
rect 414570 223718 414806 223954
rect 413930 223398 414166 223634
rect 414250 223398 414486 223634
rect 414570 223398 414806 223634
rect 303930 219218 304166 219454
rect 304250 219218 304486 219454
rect 304570 219218 304806 219454
rect 303930 218898 304166 219134
rect 304250 218898 304486 219134
rect 304570 218898 304806 219134
rect 323930 219218 324166 219454
rect 324250 219218 324486 219454
rect 324570 219218 324806 219454
rect 323930 218898 324166 219134
rect 324250 218898 324486 219134
rect 324570 218898 324806 219134
rect 343930 219218 344166 219454
rect 344250 219218 344486 219454
rect 344570 219218 344806 219454
rect 343930 218898 344166 219134
rect 344250 218898 344486 219134
rect 344570 218898 344806 219134
rect 363930 219218 364166 219454
rect 364250 219218 364486 219454
rect 364570 219218 364806 219454
rect 363930 218898 364166 219134
rect 364250 218898 364486 219134
rect 364570 218898 364806 219134
rect 383930 219218 384166 219454
rect 384250 219218 384486 219454
rect 384570 219218 384806 219454
rect 383930 218898 384166 219134
rect 384250 218898 384486 219134
rect 384570 218898 384806 219134
rect 403930 219218 404166 219454
rect 404250 219218 404486 219454
rect 404570 219218 404806 219454
rect 403930 218898 404166 219134
rect 404250 218898 404486 219134
rect 404570 218898 404806 219134
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 313930 151718 314166 151954
rect 314250 151718 314486 151954
rect 314570 151718 314806 151954
rect 313930 151398 314166 151634
rect 314250 151398 314486 151634
rect 314570 151398 314806 151634
rect 333930 151718 334166 151954
rect 334250 151718 334486 151954
rect 334570 151718 334806 151954
rect 333930 151398 334166 151634
rect 334250 151398 334486 151634
rect 334570 151398 334806 151634
rect 353930 151718 354166 151954
rect 354250 151718 354486 151954
rect 354570 151718 354806 151954
rect 353930 151398 354166 151634
rect 354250 151398 354486 151634
rect 354570 151398 354806 151634
rect 373930 151718 374166 151954
rect 374250 151718 374486 151954
rect 374570 151718 374806 151954
rect 373930 151398 374166 151634
rect 374250 151398 374486 151634
rect 374570 151398 374806 151634
rect 393930 151718 394166 151954
rect 394250 151718 394486 151954
rect 394570 151718 394806 151954
rect 393930 151398 394166 151634
rect 394250 151398 394486 151634
rect 394570 151398 394806 151634
rect 413930 151718 414166 151954
rect 414250 151718 414486 151954
rect 414570 151718 414806 151954
rect 413930 151398 414166 151634
rect 414250 151398 414486 151634
rect 414570 151398 414806 151634
rect 303930 147218 304166 147454
rect 304250 147218 304486 147454
rect 304570 147218 304806 147454
rect 303930 146898 304166 147134
rect 304250 146898 304486 147134
rect 304570 146898 304806 147134
rect 323930 147218 324166 147454
rect 324250 147218 324486 147454
rect 324570 147218 324806 147454
rect 323930 146898 324166 147134
rect 324250 146898 324486 147134
rect 324570 146898 324806 147134
rect 343930 147218 344166 147454
rect 344250 147218 344486 147454
rect 344570 147218 344806 147454
rect 343930 146898 344166 147134
rect 344250 146898 344486 147134
rect 344570 146898 344806 147134
rect 363930 147218 364166 147454
rect 364250 147218 364486 147454
rect 364570 147218 364806 147454
rect 363930 146898 364166 147134
rect 364250 146898 364486 147134
rect 364570 146898 364806 147134
rect 383930 147218 384166 147454
rect 384250 147218 384486 147454
rect 384570 147218 384806 147454
rect 383930 146898 384166 147134
rect 384250 146898 384486 147134
rect 384570 146898 384806 147134
rect 403930 147218 404166 147454
rect 404250 147218 404486 147454
rect 404570 147218 404806 147454
rect 403930 146898 404166 147134
rect 404250 146898 404486 147134
rect 404570 146898 404806 147134
rect 313930 115718 314166 115954
rect 314250 115718 314486 115954
rect 314570 115718 314806 115954
rect 313930 115398 314166 115634
rect 314250 115398 314486 115634
rect 314570 115398 314806 115634
rect 333930 115718 334166 115954
rect 334250 115718 334486 115954
rect 334570 115718 334806 115954
rect 333930 115398 334166 115634
rect 334250 115398 334486 115634
rect 334570 115398 334806 115634
rect 353930 115718 354166 115954
rect 354250 115718 354486 115954
rect 354570 115718 354806 115954
rect 353930 115398 354166 115634
rect 354250 115398 354486 115634
rect 354570 115398 354806 115634
rect 373930 115718 374166 115954
rect 374250 115718 374486 115954
rect 374570 115718 374806 115954
rect 373930 115398 374166 115634
rect 374250 115398 374486 115634
rect 374570 115398 374806 115634
rect 393930 115718 394166 115954
rect 394250 115718 394486 115954
rect 394570 115718 394806 115954
rect 393930 115398 394166 115634
rect 394250 115398 394486 115634
rect 394570 115398 394806 115634
rect 413930 115718 414166 115954
rect 414250 115718 414486 115954
rect 414570 115718 414806 115954
rect 413930 115398 414166 115634
rect 414250 115398 414486 115634
rect 414570 115398 414806 115634
rect 303930 111218 304166 111454
rect 304250 111218 304486 111454
rect 304570 111218 304806 111454
rect 303930 110898 304166 111134
rect 304250 110898 304486 111134
rect 304570 110898 304806 111134
rect 323930 111218 324166 111454
rect 324250 111218 324486 111454
rect 324570 111218 324806 111454
rect 323930 110898 324166 111134
rect 324250 110898 324486 111134
rect 324570 110898 324806 111134
rect 343930 111218 344166 111454
rect 344250 111218 344486 111454
rect 344570 111218 344806 111454
rect 343930 110898 344166 111134
rect 344250 110898 344486 111134
rect 344570 110898 344806 111134
rect 363930 111218 364166 111454
rect 364250 111218 364486 111454
rect 364570 111218 364806 111454
rect 363930 110898 364166 111134
rect 364250 110898 364486 111134
rect 364570 110898 364806 111134
rect 383930 111218 384166 111454
rect 384250 111218 384486 111454
rect 384570 111218 384806 111454
rect 383930 110898 384166 111134
rect 384250 110898 384486 111134
rect 384570 110898 384806 111134
rect 403930 111218 404166 111454
rect 404250 111218 404486 111454
rect 404570 111218 404806 111454
rect 403930 110898 404166 111134
rect 404250 110898 404486 111134
rect 404570 110898 404806 111134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 213930 43718 214166 43954
rect 214250 43718 214486 43954
rect 214570 43718 214806 43954
rect 213930 43398 214166 43634
rect 214250 43398 214486 43634
rect 214570 43398 214806 43634
rect 233930 43718 234166 43954
rect 234250 43718 234486 43954
rect 234570 43718 234806 43954
rect 233930 43398 234166 43634
rect 234250 43398 234486 43634
rect 234570 43398 234806 43634
rect 253930 43718 254166 43954
rect 254250 43718 254486 43954
rect 254570 43718 254806 43954
rect 253930 43398 254166 43634
rect 254250 43398 254486 43634
rect 254570 43398 254806 43634
rect 273930 43718 274166 43954
rect 274250 43718 274486 43954
rect 274570 43718 274806 43954
rect 273930 43398 274166 43634
rect 274250 43398 274486 43634
rect 274570 43398 274806 43634
rect 293930 43718 294166 43954
rect 294250 43718 294486 43954
rect 294570 43718 294806 43954
rect 293930 43398 294166 43634
rect 294250 43398 294486 43634
rect 294570 43398 294806 43634
rect 313930 43718 314166 43954
rect 314250 43718 314486 43954
rect 314570 43718 314806 43954
rect 313930 43398 314166 43634
rect 314250 43398 314486 43634
rect 314570 43398 314806 43634
rect 333930 43718 334166 43954
rect 334250 43718 334486 43954
rect 334570 43718 334806 43954
rect 333930 43398 334166 43634
rect 334250 43398 334486 43634
rect 334570 43398 334806 43634
rect 353930 43718 354166 43954
rect 354250 43718 354486 43954
rect 354570 43718 354806 43954
rect 353930 43398 354166 43634
rect 354250 43398 354486 43634
rect 354570 43398 354806 43634
rect 373930 43718 374166 43954
rect 374250 43718 374486 43954
rect 374570 43718 374806 43954
rect 373930 43398 374166 43634
rect 374250 43398 374486 43634
rect 374570 43398 374806 43634
rect 393930 43718 394166 43954
rect 394250 43718 394486 43954
rect 394570 43718 394806 43954
rect 393930 43398 394166 43634
rect 394250 43398 394486 43634
rect 394570 43398 394806 43634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 203930 39218 204166 39454
rect 204250 39218 204486 39454
rect 204570 39218 204806 39454
rect 203930 38898 204166 39134
rect 204250 38898 204486 39134
rect 204570 38898 204806 39134
rect 223930 39218 224166 39454
rect 224250 39218 224486 39454
rect 224570 39218 224806 39454
rect 223930 38898 224166 39134
rect 224250 38898 224486 39134
rect 224570 38898 224806 39134
rect 243930 39218 244166 39454
rect 244250 39218 244486 39454
rect 244570 39218 244806 39454
rect 243930 38898 244166 39134
rect 244250 38898 244486 39134
rect 244570 38898 244806 39134
rect 263930 39218 264166 39454
rect 264250 39218 264486 39454
rect 264570 39218 264806 39454
rect 263930 38898 264166 39134
rect 264250 38898 264486 39134
rect 264570 38898 264806 39134
rect 283930 39218 284166 39454
rect 284250 39218 284486 39454
rect 284570 39218 284806 39454
rect 283930 38898 284166 39134
rect 284250 38898 284486 39134
rect 284570 38898 284806 39134
rect 303930 39218 304166 39454
rect 304250 39218 304486 39454
rect 304570 39218 304806 39454
rect 303930 38898 304166 39134
rect 304250 38898 304486 39134
rect 304570 38898 304806 39134
rect 323930 39218 324166 39454
rect 324250 39218 324486 39454
rect 324570 39218 324806 39454
rect 323930 38898 324166 39134
rect 324250 38898 324486 39134
rect 324570 38898 324806 39134
rect 343930 39218 344166 39454
rect 344250 39218 344486 39454
rect 344570 39218 344806 39454
rect 343930 38898 344166 39134
rect 344250 38898 344486 39134
rect 344570 38898 344806 39134
rect 363930 39218 364166 39454
rect 364250 39218 364486 39454
rect 364570 39218 364806 39454
rect 363930 38898 364166 39134
rect 364250 38898 364486 39134
rect 364570 38898 364806 39134
rect 383930 39218 384166 39454
rect 384250 39218 384486 39454
rect 384570 39218 384806 39454
rect 383930 38898 384166 39134
rect 384250 38898 384486 39134
rect 384570 38898 384806 39134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 79610 43954
rect 79846 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 79610 43634
rect 79846 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 64250 39454
rect 64486 39218 94970 39454
rect 95206 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 64250 39134
rect 64486 38898 94970 39134
rect 95206 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use controller_core  controller_core_mod
timestamp 0
transform 1 0 200000 0 1 24000
box -800 -800 198812 30800
use driver_core  driver_core_0
timestamp 0
transform 1 0 20000 0 1 78000
box 1066 -800 118902 77840
use driver_core  driver_core_1
timestamp 0
transform 1 0 20000 0 1 206000
box 1066 -800 118902 77840
use driver_core  driver_core_2
timestamp 0
transform 1 0 20000 0 1 334000
box 1066 -800 118902 77840
use driver_core  driver_core_3
timestamp 0
transform 1 0 20000 0 1 462000
box 1066 -800 118902 77840
use driver_core  driver_core_4
timestamp 0
transform 1 0 20000 0 1 588000
box 1066 -800 118902 77840
use driver_core  driver_core_5
timestamp 0
transform 1 0 300000 0 1 588000
box 1066 -800 118902 77840
use driver_core  driver_core_6
timestamp 0
transform 1 0 300000 0 1 462000
box 1066 -800 118902 77840
use driver_core  driver_core_7
timestamp 0
transform 1 0 300000 0 1 334000
box 1066 -800 118902 77840
use driver_core  driver_core_8
timestamp 0
transform 1 0 300000 0 1 206000
box 1066 -800 118902 77840
use driver_core  driver_core_9
timestamp 0
transform 1 0 300000 0 1 78000
box 1066 -800 118902 77840
use spi_controller  spi_controller_mod
timestamp 0
transform 1 0 60000 0 1 24000
box 0 0 40000 37584
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 288000 38414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 670000 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 288000 74414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 670000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 288000 110414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 670000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 56000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 56000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 56000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 288000 326414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 670000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 288000 362414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 670000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 288000 398414 332000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 670000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 670000 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 670000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 670000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 56000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 56000 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 670000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 670000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 670000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 670000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 160000 20414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 416000 20414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 160000 56414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 416000 56414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 160000 92414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 416000 92414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 160000 128414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 416000 128414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 56000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 56000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 56000 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 160000 308414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 416000 308414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 160000 344414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 416000 344414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 160000 380414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 416000 380414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 160000 416414 204000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 416000 416414 460000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 670000 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 670000 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 670000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 670000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 56000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 56000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 56000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 670000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 670000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 670000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 416000 24914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 670000 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 416000 60914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 670000 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 416000 96914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 670000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 416000 132914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 670000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 56000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 56000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 56000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 416000 312914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 670000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 416000 348914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 670000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 416000 384914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 670000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 416000 420914 460000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 670000 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 670000 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 670000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 670000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 670000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 56000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 56000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 56000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 670000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 670000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 670000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 288000 42914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 544000 42914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 670000 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 288000 78914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 544000 78914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 670000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 288000 114914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 544000 114914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 670000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 56000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 56000 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 56000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 288000 330914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 544000 330914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 670000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 288000 366914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 544000 366914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 670000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 288000 402914 332000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 544000 402914 586000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 670000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 160000 51914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 670000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 160000 87914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 670000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 160000 123914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 670000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 56000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 56000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 160000 303914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 670000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 160000 339914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 670000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 160000 375914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 670000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 160000 411914 204000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 670000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
