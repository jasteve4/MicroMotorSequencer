VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO controller_core
  CLASS BLOCK ;
  FOREIGN controller_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 150.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 -4.000 338.470 4.000 ;
    END
  END clock
  PIN clock_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 146.000 280.510 154.000 ;
    END
  END clock_out[0]
  PIN clock_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 146.000 288.790 154.000 ;
    END
  END clock_out[1]
  PIN clock_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 146.000 297.070 154.000 ;
    END
  END clock_out[2]
  PIN clock_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 146.000 305.350 154.000 ;
    END
  END clock_out[3]
  PIN clock_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 146.000 313.630 154.000 ;
    END
  END clock_out[4]
  PIN clock_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 146.000 321.910 154.000 ;
    END
  END clock_out[5]
  PIN clock_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 146.000 330.190 154.000 ;
    END
  END clock_out[6]
  PIN clock_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 146.000 338.470 154.000 ;
    END
  END clock_out[7]
  PIN clock_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 146.000 346.750 154.000 ;
    END
  END clock_out[8]
  PIN clock_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 146.000 355.030 154.000 ;
    END
  END clock_out[9]
  PIN col_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 146.000 512.350 154.000 ;
    END
  END col_select_left[0]
  PIN col_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 146.000 520.630 154.000 ;
    END
  END col_select_left[1]
  PIN col_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 146.000 528.910 154.000 ;
    END
  END col_select_left[2]
  PIN col_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 146.000 537.190 154.000 ;
    END
  END col_select_left[3]
  PIN col_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 146.000 545.470 154.000 ;
    END
  END col_select_left[4]
  PIN col_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 146.000 553.750 154.000 ;
    END
  END col_select_left[5]
  PIN col_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 146.000 462.670 154.000 ;
    END
  END col_select_right[0]
  PIN col_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 146.000 470.950 154.000 ;
    END
  END col_select_right[1]
  PIN col_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 146.000 479.230 154.000 ;
    END
  END col_select_right[2]
  PIN col_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 146.000 487.510 154.000 ;
    END
  END col_select_right[3]
  PIN col_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 146.000 495.790 154.000 ;
    END
  END col_select_right[4]
  PIN col_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 146.000 504.070 154.000 ;
    END
  END col_select_right[5]
  PIN data_out_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 146.000 694.510 154.000 ;
    END
  END data_out_left[0]
  PIN data_out_left[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 146.000 777.310 154.000 ;
    END
  END data_out_left[10]
  PIN data_out_left[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 146.000 785.590 154.000 ;
    END
  END data_out_left[11]
  PIN data_out_left[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 146.000 793.870 154.000 ;
    END
  END data_out_left[12]
  PIN data_out_left[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 146.000 802.150 154.000 ;
    END
  END data_out_left[13]
  PIN data_out_left[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 146.000 810.430 154.000 ;
    END
  END data_out_left[14]
  PIN data_out_left[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 146.000 818.710 154.000 ;
    END
  END data_out_left[15]
  PIN data_out_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 146.000 702.790 154.000 ;
    END
  END data_out_left[1]
  PIN data_out_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 146.000 711.070 154.000 ;
    END
  END data_out_left[2]
  PIN data_out_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 146.000 719.350 154.000 ;
    END
  END data_out_left[3]
  PIN data_out_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 146.000 727.630 154.000 ;
    END
  END data_out_left[4]
  PIN data_out_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 146.000 735.910 154.000 ;
    END
  END data_out_left[5]
  PIN data_out_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 146.000 744.190 154.000 ;
    END
  END data_out_left[6]
  PIN data_out_left[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 146.000 752.470 154.000 ;
    END
  END data_out_left[7]
  PIN data_out_left[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 146.000 760.750 154.000 ;
    END
  END data_out_left[8]
  PIN data_out_left[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 146.000 769.030 154.000 ;
    END
  END data_out_left[9]
  PIN data_out_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 146.000 562.030 154.000 ;
    END
  END data_out_right[0]
  PIN data_out_right[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 146.000 644.830 154.000 ;
    END
  END data_out_right[10]
  PIN data_out_right[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 146.000 653.110 154.000 ;
    END
  END data_out_right[11]
  PIN data_out_right[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 146.000 661.390 154.000 ;
    END
  END data_out_right[12]
  PIN data_out_right[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 146.000 669.670 154.000 ;
    END
  END data_out_right[13]
  PIN data_out_right[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 146.000 677.950 154.000 ;
    END
  END data_out_right[14]
  PIN data_out_right[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 146.000 686.230 154.000 ;
    END
  END data_out_right[15]
  PIN data_out_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 146.000 570.310 154.000 ;
    END
  END data_out_right[1]
  PIN data_out_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 146.000 578.590 154.000 ;
    END
  END data_out_right[2]
  PIN data_out_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 146.000 586.870 154.000 ;
    END
  END data_out_right[3]
  PIN data_out_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 146.000 595.150 154.000 ;
    END
  END data_out_right[4]
  PIN data_out_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 146.000 603.430 154.000 ;
    END
  END data_out_right[5]
  PIN data_out_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 146.000 611.710 154.000 ;
    END
  END data_out_right[6]
  PIN data_out_right[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 146.000 619.990 154.000 ;
    END
  END data_out_right[7]
  PIN data_out_right[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 146.000 628.270 154.000 ;
    END
  END data_out_right[8]
  PIN data_out_right[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 146.000 636.550 154.000 ;
    END
  END data_out_right[9]
  PIN inverter_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 146.000 909.790 154.000 ;
    END
  END inverter_select[0]
  PIN inverter_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 146.000 918.070 154.000 ;
    END
  END inverter_select[1]
  PIN inverter_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 146.000 926.350 154.000 ;
    END
  END inverter_select[2]
  PIN inverter_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 146.000 934.630 154.000 ;
    END
  END inverter_select[3]
  PIN inverter_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 146.000 942.910 154.000 ;
    END
  END inverter_select[4]
  PIN inverter_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 146.000 951.190 154.000 ;
    END
  END inverter_select[5]
  PIN inverter_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 146.000 959.470 154.000 ;
    END
  END inverter_select[6]
  PIN inverter_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 146.000 967.750 154.000 ;
    END
  END inverter_select[7]
  PIN inverter_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 146.000 976.030 154.000 ;
    END
  END inverter_select[8]
  PIN inverter_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 146.000 984.310 154.000 ;
    END
  END inverter_select[9]
  PIN io_control_trigger_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 -4.000 751.090 4.000 ;
    END
  END io_control_trigger_in
  PIN io_control_trigger_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 -4.000 769.030 4.000 ;
    END
  END io_control_trigger_oeb
  PIN io_driver_io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 -4.000 822.850 4.000 ;
    END
  END io_driver_io_oeb[0]
  PIN io_driver_io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 -4.000 840.790 4.000 ;
    END
  END io_driver_io_oeb[1]
  PIN io_driver_io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 -4.000 858.730 4.000 ;
    END
  END io_driver_io_oeb[2]
  PIN io_driver_io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 -4.000 876.670 4.000 ;
    END
  END io_driver_io_oeb[3]
  PIN io_driver_io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 -4.000 894.610 4.000 ;
    END
  END io_driver_io_oeb[4]
  PIN io_driver_io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 -4.000 912.550 4.000 ;
    END
  END io_driver_io_oeb[5]
  PIN io_driver_io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 -4.000 930.490 4.000 ;
    END
  END io_driver_io_oeb[6]
  PIN io_driver_io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 -4.000 948.430 4.000 ;
    END
  END io_driver_io_oeb[7]
  PIN io_driver_io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 -4.000 966.370 4.000 ;
    END
  END io_driver_io_oeb[8]
  PIN io_driver_io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 -4.000 984.310 4.000 ;
    END
  END io_driver_io_oeb[9]
  PIN io_latch_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 -4.000 715.210 4.000 ;
    END
  END io_latch_data_in
  PIN io_latch_data_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 -4.000 733.150 4.000 ;
    END
  END io_latch_data_oeb
  PIN io_reset_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 -4.000 679.330 4.000 ;
    END
  END io_reset_n_in
  PIN io_reset_n_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 -4.000 697.270 4.000 ;
    END
  END io_reset_n_oeb
  PIN io_update_cycle_complete_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 -4.000 804.910 4.000 ;
    END
  END io_update_cycle_complete_oeb
  PIN io_update_cycle_complete_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 -4.000 786.970 4.000 ;
    END
  END io_update_cycle_complete_out
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 -4.000 194.950 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 -4.000 212.890 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 -4.000 230.830 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 -4.000 248.770 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 -4.000 266.710 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 -4.000 284.650 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 -4.000 302.590 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 -4.000 320.530 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 -4.000 33.490 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 -4.000 51.430 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 -4.000 69.370 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 -4.000 105.250 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 -4.000 123.190 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 -4.000 141.130 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 -4.000 159.070 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 -4.000 177.010 4.000 ;
    END
  END la_data_in[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 -4.000 356.410 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 -4.000 535.810 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 -4.000 553.750 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 -4.000 571.690 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 -4.000 589.630 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 -4.000 607.570 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 -4.000 625.510 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 -4.000 643.450 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 -4.000 661.390 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 -4.000 374.350 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 -4.000 392.290 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 -4.000 410.230 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 -4.000 428.170 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 -4.000 446.110 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 -4.000 464.050 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 -4.000 481.990 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -4.000 499.930 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 -4.000 517.870 4.000 ;
    END
  END la_oenb[9]
  PIN mem_address_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 146.000 114.910 154.000 ;
    END
  END mem_address_left[0]
  PIN mem_address_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 146.000 123.190 154.000 ;
    END
  END mem_address_left[1]
  PIN mem_address_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 146.000 131.470 154.000 ;
    END
  END mem_address_left[2]
  PIN mem_address_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 146.000 139.750 154.000 ;
    END
  END mem_address_left[3]
  PIN mem_address_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 146.000 148.030 154.000 ;
    END
  END mem_address_left[4]
  PIN mem_address_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 146.000 156.310 154.000 ;
    END
  END mem_address_left[5]
  PIN mem_address_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 146.000 164.590 154.000 ;
    END
  END mem_address_left[6]
  PIN mem_address_left[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 146.000 172.870 154.000 ;
    END
  END mem_address_left[7]
  PIN mem_address_left[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 146.000 181.150 154.000 ;
    END
  END mem_address_left[8]
  PIN mem_address_left[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 146.000 189.430 154.000 ;
    END
  END mem_address_left[9]
  PIN mem_address_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 146.000 32.110 154.000 ;
    END
  END mem_address_right[0]
  PIN mem_address_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 146.000 40.390 154.000 ;
    END
  END mem_address_right[1]
  PIN mem_address_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 154.000 ;
    END
  END mem_address_right[2]
  PIN mem_address_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 146.000 56.950 154.000 ;
    END
  END mem_address_right[3]
  PIN mem_address_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 146.000 65.230 154.000 ;
    END
  END mem_address_right[4]
  PIN mem_address_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 146.000 73.510 154.000 ;
    END
  END mem_address_right[5]
  PIN mem_address_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 146.000 81.790 154.000 ;
    END
  END mem_address_right[6]
  PIN mem_address_right[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 146.000 90.070 154.000 ;
    END
  END mem_address_right[7]
  PIN mem_address_right[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 146.000 98.350 154.000 ;
    END
  END mem_address_right[8]
  PIN mem_address_right[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 146.000 106.630 154.000 ;
    END
  END mem_address_right[9]
  PIN mem_write_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 146.000 197.710 154.000 ;
    END
  END mem_write_n[0]
  PIN mem_write_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 146.000 205.990 154.000 ;
    END
  END mem_write_n[1]
  PIN mem_write_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 146.000 214.270 154.000 ;
    END
  END mem_write_n[2]
  PIN mem_write_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 146.000 222.550 154.000 ;
    END
  END mem_write_n[3]
  PIN mem_write_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 146.000 230.830 154.000 ;
    END
  END mem_write_n[4]
  PIN mem_write_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 146.000 239.110 154.000 ;
    END
  END mem_write_n[5]
  PIN mem_write_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 146.000 247.390 154.000 ;
    END
  END mem_write_n[6]
  PIN mem_write_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 146.000 255.670 154.000 ;
    END
  END mem_write_n[7]
  PIN mem_write_n[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 146.000 263.950 154.000 ;
    END
  END mem_write_n[8]
  PIN mem_write_n[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 146.000 272.230 154.000 ;
    END
  END mem_write_n[9]
  PIN output_active_left
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 146.000 23.830 154.000 ;
    END
  END output_active_left
  PIN output_active_right
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 146.000 15.550 154.000 ;
    END
  END output_active_right
  PIN row_col_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 146.000 826.990 154.000 ;
    END
  END row_col_select[0]
  PIN row_col_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 146.000 835.270 154.000 ;
    END
  END row_col_select[1]
  PIN row_col_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 146.000 843.550 154.000 ;
    END
  END row_col_select[2]
  PIN row_col_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 146.000 851.830 154.000 ;
    END
  END row_col_select[3]
  PIN row_col_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 146.000 860.110 154.000 ;
    END
  END row_col_select[4]
  PIN row_col_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 146.000 868.390 154.000 ;
    END
  END row_col_select[5]
  PIN row_col_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 146.000 876.670 154.000 ;
    END
  END row_col_select[6]
  PIN row_col_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 146.000 884.950 154.000 ;
    END
  END row_col_select[7]
  PIN row_col_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 146.000 893.230 154.000 ;
    END
  END row_col_select[8]
  PIN row_col_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 146.000 901.510 154.000 ;
    END
  END row_col_select[9]
  PIN row_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 146.000 412.990 154.000 ;
    END
  END row_select_left[0]
  PIN row_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 146.000 421.270 154.000 ;
    END
  END row_select_left[1]
  PIN row_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 146.000 429.550 154.000 ;
    END
  END row_select_left[2]
  PIN row_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 146.000 437.830 154.000 ;
    END
  END row_select_left[3]
  PIN row_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 146.000 446.110 154.000 ;
    END
  END row_select_left[4]
  PIN row_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 146.000 454.390 154.000 ;
    END
  END row_select_left[5]
  PIN row_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 146.000 363.310 154.000 ;
    END
  END row_select_right[0]
  PIN row_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 146.000 371.590 154.000 ;
    END
  END row_select_right[1]
  PIN row_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 146.000 379.870 154.000 ;
    END
  END row_select_right[2]
  PIN row_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 146.000 388.150 154.000 ;
    END
  END row_select_right[3]
  PIN row_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 146.000 396.430 154.000 ;
    END
  END row_select_right[4]
  PIN row_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 146.000 404.710 154.000 ;
    END
  END row_select_right[5]
  PIN spi_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 13.640 4.000 14.240 ;
    END
  END spi_data[0]
  PIN spi_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 54.440 4.000 55.040 ;
    END
  END spi_data[10]
  PIN spi_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 58.520 4.000 59.120 ;
    END
  END spi_data[11]
  PIN spi_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 62.600 4.000 63.200 ;
    END
  END spi_data[12]
  PIN spi_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 66.680 4.000 67.280 ;
    END
  END spi_data[13]
  PIN spi_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 70.760 4.000 71.360 ;
    END
  END spi_data[14]
  PIN spi_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 74.840 4.000 75.440 ;
    END
  END spi_data[15]
  PIN spi_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 78.920 4.000 79.520 ;
    END
  END spi_data[16]
  PIN spi_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 83.000 4.000 83.600 ;
    END
  END spi_data[17]
  PIN spi_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 87.080 4.000 87.680 ;
    END
  END spi_data[18]
  PIN spi_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 91.160 4.000 91.760 ;
    END
  END spi_data[19]
  PIN spi_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.720 4.000 18.320 ;
    END
  END spi_data[1]
  PIN spi_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 95.240 4.000 95.840 ;
    END
  END spi_data[20]
  PIN spi_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 99.320 4.000 99.920 ;
    END
  END spi_data[21]
  PIN spi_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 103.400 4.000 104.000 ;
    END
  END spi_data[22]
  PIN spi_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 107.480 4.000 108.080 ;
    END
  END spi_data[23]
  PIN spi_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 111.560 4.000 112.160 ;
    END
  END spi_data[24]
  PIN spi_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 115.640 4.000 116.240 ;
    END
  END spi_data[25]
  PIN spi_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 119.720 4.000 120.320 ;
    END
  END spi_data[26]
  PIN spi_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 123.800 4.000 124.400 ;
    END
  END spi_data[27]
  PIN spi_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 127.880 4.000 128.480 ;
    END
  END spi_data[28]
  PIN spi_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 131.960 4.000 132.560 ;
    END
  END spi_data[29]
  PIN spi_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 21.800 4.000 22.400 ;
    END
  END spi_data[2]
  PIN spi_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 136.040 4.000 136.640 ;
    END
  END spi_data[30]
  PIN spi_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 140.120 4.000 140.720 ;
    END
  END spi_data[31]
  PIN spi_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 25.880 4.000 26.480 ;
    END
  END spi_data[3]
  PIN spi_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.960 4.000 30.560 ;
    END
  END spi_data[4]
  PIN spi_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 34.040 4.000 34.640 ;
    END
  END spi_data[5]
  PIN spi_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 38.120 4.000 38.720 ;
    END
  END spi_data[6]
  PIN spi_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 42.200 4.000 42.800 ;
    END
  END spi_data[7]
  PIN spi_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 46.280 4.000 46.880 ;
    END
  END spi_data[8]
  PIN spi_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 50.360 4.000 50.960 ;
    END
  END spi_data[9]
  PIN spi_data_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 9.560 4.000 10.160 ;
    END
  END spi_data_clock
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.340 10.640 624.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.340 10.640 724.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.340 10.640 824.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 919.340 10.640 924.340 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 669.340 10.640 674.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.340 10.640 774.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 869.340 10.640 874.340 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 969.340 10.640 974.340 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 138.805 ;
      LAYER met1 ;
        RECT 5.520 5.480 994.060 142.420 ;
      LAYER met2 ;
        RECT 6.990 145.720 14.990 146.610 ;
        RECT 15.830 145.720 23.270 146.610 ;
        RECT 24.110 145.720 31.550 146.610 ;
        RECT 32.390 145.720 39.830 146.610 ;
        RECT 40.670 145.720 48.110 146.610 ;
        RECT 48.950 145.720 56.390 146.610 ;
        RECT 57.230 145.720 64.670 146.610 ;
        RECT 65.510 145.720 72.950 146.610 ;
        RECT 73.790 145.720 81.230 146.610 ;
        RECT 82.070 145.720 89.510 146.610 ;
        RECT 90.350 145.720 97.790 146.610 ;
        RECT 98.630 145.720 106.070 146.610 ;
        RECT 106.910 145.720 114.350 146.610 ;
        RECT 115.190 145.720 122.630 146.610 ;
        RECT 123.470 145.720 130.910 146.610 ;
        RECT 131.750 145.720 139.190 146.610 ;
        RECT 140.030 145.720 147.470 146.610 ;
        RECT 148.310 145.720 155.750 146.610 ;
        RECT 156.590 145.720 164.030 146.610 ;
        RECT 164.870 145.720 172.310 146.610 ;
        RECT 173.150 145.720 180.590 146.610 ;
        RECT 181.430 145.720 188.870 146.610 ;
        RECT 189.710 145.720 197.150 146.610 ;
        RECT 197.990 145.720 205.430 146.610 ;
        RECT 206.270 145.720 213.710 146.610 ;
        RECT 214.550 145.720 221.990 146.610 ;
        RECT 222.830 145.720 230.270 146.610 ;
        RECT 231.110 145.720 238.550 146.610 ;
        RECT 239.390 145.720 246.830 146.610 ;
        RECT 247.670 145.720 255.110 146.610 ;
        RECT 255.950 145.720 263.390 146.610 ;
        RECT 264.230 145.720 271.670 146.610 ;
        RECT 272.510 145.720 279.950 146.610 ;
        RECT 280.790 145.720 288.230 146.610 ;
        RECT 289.070 145.720 296.510 146.610 ;
        RECT 297.350 145.720 304.790 146.610 ;
        RECT 305.630 145.720 313.070 146.610 ;
        RECT 313.910 145.720 321.350 146.610 ;
        RECT 322.190 145.720 329.630 146.610 ;
        RECT 330.470 145.720 337.910 146.610 ;
        RECT 338.750 145.720 346.190 146.610 ;
        RECT 347.030 145.720 354.470 146.610 ;
        RECT 355.310 145.720 362.750 146.610 ;
        RECT 363.590 145.720 371.030 146.610 ;
        RECT 371.870 145.720 379.310 146.610 ;
        RECT 380.150 145.720 387.590 146.610 ;
        RECT 388.430 145.720 395.870 146.610 ;
        RECT 396.710 145.720 404.150 146.610 ;
        RECT 404.990 145.720 412.430 146.610 ;
        RECT 413.270 145.720 420.710 146.610 ;
        RECT 421.550 145.720 428.990 146.610 ;
        RECT 429.830 145.720 437.270 146.610 ;
        RECT 438.110 145.720 445.550 146.610 ;
        RECT 446.390 145.720 453.830 146.610 ;
        RECT 454.670 145.720 462.110 146.610 ;
        RECT 462.950 145.720 470.390 146.610 ;
        RECT 471.230 145.720 478.670 146.610 ;
        RECT 479.510 145.720 486.950 146.610 ;
        RECT 487.790 145.720 495.230 146.610 ;
        RECT 496.070 145.720 503.510 146.610 ;
        RECT 504.350 145.720 511.790 146.610 ;
        RECT 512.630 145.720 520.070 146.610 ;
        RECT 520.910 145.720 528.350 146.610 ;
        RECT 529.190 145.720 536.630 146.610 ;
        RECT 537.470 145.720 544.910 146.610 ;
        RECT 545.750 145.720 553.190 146.610 ;
        RECT 554.030 145.720 561.470 146.610 ;
        RECT 562.310 145.720 569.750 146.610 ;
        RECT 570.590 145.720 578.030 146.610 ;
        RECT 578.870 145.720 586.310 146.610 ;
        RECT 587.150 145.720 594.590 146.610 ;
        RECT 595.430 145.720 602.870 146.610 ;
        RECT 603.710 145.720 611.150 146.610 ;
        RECT 611.990 145.720 619.430 146.610 ;
        RECT 620.270 145.720 627.710 146.610 ;
        RECT 628.550 145.720 635.990 146.610 ;
        RECT 636.830 145.720 644.270 146.610 ;
        RECT 645.110 145.720 652.550 146.610 ;
        RECT 653.390 145.720 660.830 146.610 ;
        RECT 661.670 145.720 669.110 146.610 ;
        RECT 669.950 145.720 677.390 146.610 ;
        RECT 678.230 145.720 685.670 146.610 ;
        RECT 686.510 145.720 693.950 146.610 ;
        RECT 694.790 145.720 702.230 146.610 ;
        RECT 703.070 145.720 710.510 146.610 ;
        RECT 711.350 145.720 718.790 146.610 ;
        RECT 719.630 145.720 727.070 146.610 ;
        RECT 727.910 145.720 735.350 146.610 ;
        RECT 736.190 145.720 743.630 146.610 ;
        RECT 744.470 145.720 751.910 146.610 ;
        RECT 752.750 145.720 760.190 146.610 ;
        RECT 761.030 145.720 768.470 146.610 ;
        RECT 769.310 145.720 776.750 146.610 ;
        RECT 777.590 145.720 785.030 146.610 ;
        RECT 785.870 145.720 793.310 146.610 ;
        RECT 794.150 145.720 801.590 146.610 ;
        RECT 802.430 145.720 809.870 146.610 ;
        RECT 810.710 145.720 818.150 146.610 ;
        RECT 818.990 145.720 826.430 146.610 ;
        RECT 827.270 145.720 834.710 146.610 ;
        RECT 835.550 145.720 842.990 146.610 ;
        RECT 843.830 145.720 851.270 146.610 ;
        RECT 852.110 145.720 859.550 146.610 ;
        RECT 860.390 145.720 867.830 146.610 ;
        RECT 868.670 145.720 876.110 146.610 ;
        RECT 876.950 145.720 884.390 146.610 ;
        RECT 885.230 145.720 892.670 146.610 ;
        RECT 893.510 145.720 900.950 146.610 ;
        RECT 901.790 145.720 909.230 146.610 ;
        RECT 910.070 145.720 917.510 146.610 ;
        RECT 918.350 145.720 925.790 146.610 ;
        RECT 926.630 145.720 934.070 146.610 ;
        RECT 934.910 145.720 942.350 146.610 ;
        RECT 943.190 145.720 950.630 146.610 ;
        RECT 951.470 145.720 958.910 146.610 ;
        RECT 959.750 145.720 967.190 146.610 ;
        RECT 968.030 145.720 975.470 146.610 ;
        RECT 976.310 145.720 983.750 146.610 ;
        RECT 984.590 145.720 987.980 146.610 ;
        RECT 6.990 4.280 987.980 145.720 ;
        RECT 6.990 3.670 14.990 4.280 ;
        RECT 15.830 3.670 32.930 4.280 ;
        RECT 33.770 3.670 50.870 4.280 ;
        RECT 51.710 3.670 68.810 4.280 ;
        RECT 69.650 3.670 86.750 4.280 ;
        RECT 87.590 3.670 104.690 4.280 ;
        RECT 105.530 3.670 122.630 4.280 ;
        RECT 123.470 3.670 140.570 4.280 ;
        RECT 141.410 3.670 158.510 4.280 ;
        RECT 159.350 3.670 176.450 4.280 ;
        RECT 177.290 3.670 194.390 4.280 ;
        RECT 195.230 3.670 212.330 4.280 ;
        RECT 213.170 3.670 230.270 4.280 ;
        RECT 231.110 3.670 248.210 4.280 ;
        RECT 249.050 3.670 266.150 4.280 ;
        RECT 266.990 3.670 284.090 4.280 ;
        RECT 284.930 3.670 302.030 4.280 ;
        RECT 302.870 3.670 319.970 4.280 ;
        RECT 320.810 3.670 337.910 4.280 ;
        RECT 338.750 3.670 355.850 4.280 ;
        RECT 356.690 3.670 373.790 4.280 ;
        RECT 374.630 3.670 391.730 4.280 ;
        RECT 392.570 3.670 409.670 4.280 ;
        RECT 410.510 3.670 427.610 4.280 ;
        RECT 428.450 3.670 445.550 4.280 ;
        RECT 446.390 3.670 463.490 4.280 ;
        RECT 464.330 3.670 481.430 4.280 ;
        RECT 482.270 3.670 499.370 4.280 ;
        RECT 500.210 3.670 517.310 4.280 ;
        RECT 518.150 3.670 535.250 4.280 ;
        RECT 536.090 3.670 553.190 4.280 ;
        RECT 554.030 3.670 571.130 4.280 ;
        RECT 571.970 3.670 589.070 4.280 ;
        RECT 589.910 3.670 607.010 4.280 ;
        RECT 607.850 3.670 624.950 4.280 ;
        RECT 625.790 3.670 642.890 4.280 ;
        RECT 643.730 3.670 660.830 4.280 ;
        RECT 661.670 3.670 678.770 4.280 ;
        RECT 679.610 3.670 696.710 4.280 ;
        RECT 697.550 3.670 714.650 4.280 ;
        RECT 715.490 3.670 732.590 4.280 ;
        RECT 733.430 3.670 750.530 4.280 ;
        RECT 751.370 3.670 768.470 4.280 ;
        RECT 769.310 3.670 786.410 4.280 ;
        RECT 787.250 3.670 804.350 4.280 ;
        RECT 805.190 3.670 822.290 4.280 ;
        RECT 823.130 3.670 840.230 4.280 ;
        RECT 841.070 3.670 858.170 4.280 ;
        RECT 859.010 3.670 876.110 4.280 ;
        RECT 876.950 3.670 894.050 4.280 ;
        RECT 894.890 3.670 911.990 4.280 ;
        RECT 912.830 3.670 929.930 4.280 ;
        RECT 930.770 3.670 947.870 4.280 ;
        RECT 948.710 3.670 965.810 4.280 ;
        RECT 966.650 3.670 983.750 4.280 ;
        RECT 984.590 3.670 987.980 4.280 ;
      LAYER met3 ;
        RECT 4.400 139.720 982.035 140.585 ;
        RECT 4.000 137.040 982.035 139.720 ;
        RECT 4.400 135.640 982.035 137.040 ;
        RECT 4.000 132.960 982.035 135.640 ;
        RECT 4.400 131.560 982.035 132.960 ;
        RECT 4.000 128.880 982.035 131.560 ;
        RECT 4.400 127.480 982.035 128.880 ;
        RECT 4.000 124.800 982.035 127.480 ;
        RECT 4.400 123.400 982.035 124.800 ;
        RECT 4.000 120.720 982.035 123.400 ;
        RECT 4.400 119.320 982.035 120.720 ;
        RECT 4.000 116.640 982.035 119.320 ;
        RECT 4.400 115.240 982.035 116.640 ;
        RECT 4.000 112.560 982.035 115.240 ;
        RECT 4.400 111.160 982.035 112.560 ;
        RECT 4.000 108.480 982.035 111.160 ;
        RECT 4.400 107.080 982.035 108.480 ;
        RECT 4.000 104.400 982.035 107.080 ;
        RECT 4.400 103.000 982.035 104.400 ;
        RECT 4.000 100.320 982.035 103.000 ;
        RECT 4.400 98.920 982.035 100.320 ;
        RECT 4.000 96.240 982.035 98.920 ;
        RECT 4.400 94.840 982.035 96.240 ;
        RECT 4.000 92.160 982.035 94.840 ;
        RECT 4.400 90.760 982.035 92.160 ;
        RECT 4.000 88.080 982.035 90.760 ;
        RECT 4.400 86.680 982.035 88.080 ;
        RECT 4.000 84.000 982.035 86.680 ;
        RECT 4.400 82.600 982.035 84.000 ;
        RECT 4.000 79.920 982.035 82.600 ;
        RECT 4.400 78.520 982.035 79.920 ;
        RECT 4.000 75.840 982.035 78.520 ;
        RECT 4.400 74.440 982.035 75.840 ;
        RECT 4.000 71.760 982.035 74.440 ;
        RECT 4.400 70.360 982.035 71.760 ;
        RECT 4.000 67.680 982.035 70.360 ;
        RECT 4.400 66.280 982.035 67.680 ;
        RECT 4.000 63.600 982.035 66.280 ;
        RECT 4.400 62.200 982.035 63.600 ;
        RECT 4.000 59.520 982.035 62.200 ;
        RECT 4.400 58.120 982.035 59.520 ;
        RECT 4.000 55.440 982.035 58.120 ;
        RECT 4.400 54.040 982.035 55.440 ;
        RECT 4.000 51.360 982.035 54.040 ;
        RECT 4.400 49.960 982.035 51.360 ;
        RECT 4.000 47.280 982.035 49.960 ;
        RECT 4.400 45.880 982.035 47.280 ;
        RECT 4.000 43.200 982.035 45.880 ;
        RECT 4.400 41.800 982.035 43.200 ;
        RECT 4.000 39.120 982.035 41.800 ;
        RECT 4.400 37.720 982.035 39.120 ;
        RECT 4.000 35.040 982.035 37.720 ;
        RECT 4.400 33.640 982.035 35.040 ;
        RECT 4.000 30.960 982.035 33.640 ;
        RECT 4.400 29.560 982.035 30.960 ;
        RECT 4.000 26.880 982.035 29.560 ;
        RECT 4.400 25.480 982.035 26.880 ;
        RECT 4.000 22.800 982.035 25.480 ;
        RECT 4.400 21.400 982.035 22.800 ;
        RECT 4.000 18.720 982.035 21.400 ;
        RECT 4.400 17.320 982.035 18.720 ;
        RECT 4.000 14.640 982.035 17.320 ;
        RECT 4.400 13.240 982.035 14.640 ;
        RECT 4.000 10.560 982.035 13.240 ;
        RECT 4.400 9.695 982.035 10.560 ;
      LAYER met4 ;
        RECT 518.255 113.735 518.585 137.185 ;
  END
END controller_core
END LIBRARY

