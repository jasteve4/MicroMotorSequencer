VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO controller_unit
  CLASS BLOCK ;
  FOREIGN controller_unit ;
  ORIGIN 0.000 0.000 ;
  SIZE 1400.000 BY 140.000 ;
  PIN clock_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 136.000 594.230 144.000 ;
    END
  END clock_out[0]
  PIN clock_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 136.000 603.430 144.000 ;
    END
  END clock_out[1]
  PIN clock_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 136.000 612.630 144.000 ;
    END
  END clock_out[2]
  PIN clock_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 136.000 621.830 144.000 ;
    END
  END clock_out[3]
  PIN clock_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 136.000 631.030 144.000 ;
    END
  END clock_out[4]
  PIN clock_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 136.000 640.230 144.000 ;
    END
  END clock_out[5]
  PIN clock_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 136.000 649.430 144.000 ;
    END
  END clock_out[6]
  PIN clock_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 136.000 658.630 144.000 ;
    END
  END clock_out[7]
  PIN clock_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 136.000 667.830 144.000 ;
    END
  END clock_out[8]
  PIN clock_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 136.000 677.030 144.000 ;
    END
  END clock_out[9]
  PIN col_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 136.000 539.030 144.000 ;
    END
  END col_select_left[0]
  PIN col_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 136.000 548.230 144.000 ;
    END
  END col_select_left[1]
  PIN col_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 136.000 557.430 144.000 ;
    END
  END col_select_left[2]
  PIN col_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 136.000 566.630 144.000 ;
    END
  END col_select_left[3]
  PIN col_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 136.000 575.830 144.000 ;
    END
  END col_select_left[4]
  PIN col_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 136.000 585.030 144.000 ;
    END
  END col_select_left[5]
  PIN col_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 136.000 483.830 144.000 ;
    END
  END col_select_right[0]
  PIN col_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 136.000 493.030 144.000 ;
    END
  END col_select_right[1]
  PIN col_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 136.000 502.230 144.000 ;
    END
  END col_select_right[2]
  PIN col_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 136.000 511.430 144.000 ;
    END
  END col_select_right[3]
  PIN col_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 136.000 520.630 144.000 ;
    END
  END col_select_right[4]
  PIN col_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 136.000 529.830 144.000 ;
    END
  END col_select_right[5]
  PIN data_out_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 136.000 962.230 144.000 ;
    END
  END data_out_left[0]
  PIN data_out_left[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 136.000 1054.230 144.000 ;
    END
  END data_out_left[10]
  PIN data_out_left[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 136.000 1063.430 144.000 ;
    END
  END data_out_left[11]
  PIN data_out_left[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 136.000 1072.630 144.000 ;
    END
  END data_out_left[12]
  PIN data_out_left[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 136.000 1081.830 144.000 ;
    END
  END data_out_left[13]
  PIN data_out_left[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 136.000 1091.030 144.000 ;
    END
  END data_out_left[14]
  PIN data_out_left[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 136.000 1100.230 144.000 ;
    END
  END data_out_left[15]
  PIN data_out_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 136.000 971.430 144.000 ;
    END
  END data_out_left[1]
  PIN data_out_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 136.000 980.630 144.000 ;
    END
  END data_out_left[2]
  PIN data_out_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 136.000 989.830 144.000 ;
    END
  END data_out_left[3]
  PIN data_out_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 136.000 999.030 144.000 ;
    END
  END data_out_left[4]
  PIN data_out_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 136.000 1008.230 144.000 ;
    END
  END data_out_left[5]
  PIN data_out_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 136.000 1017.430 144.000 ;
    END
  END data_out_left[6]
  PIN data_out_left[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 136.000 1026.630 144.000 ;
    END
  END data_out_left[7]
  PIN data_out_left[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 136.000 1035.830 144.000 ;
    END
  END data_out_left[8]
  PIN data_out_left[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 136.000 1045.030 144.000 ;
    END
  END data_out_left[9]
  PIN data_out_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 136.000 815.030 144.000 ;
    END
  END data_out_right[0]
  PIN data_out_right[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 136.000 907.030 144.000 ;
    END
  END data_out_right[10]
  PIN data_out_right[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 136.000 916.230 144.000 ;
    END
  END data_out_right[11]
  PIN data_out_right[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.150 136.000 925.430 144.000 ;
    END
  END data_out_right[12]
  PIN data_out_right[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 136.000 934.630 144.000 ;
    END
  END data_out_right[13]
  PIN data_out_right[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 136.000 943.830 144.000 ;
    END
  END data_out_right[14]
  PIN data_out_right[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 136.000 953.030 144.000 ;
    END
  END data_out_right[15]
  PIN data_out_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 136.000 824.230 144.000 ;
    END
  END data_out_right[1]
  PIN data_out_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 136.000 833.430 144.000 ;
    END
  END data_out_right[2]
  PIN data_out_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 136.000 842.630 144.000 ;
    END
  END data_out_right[3]
  PIN data_out_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 136.000 851.830 144.000 ;
    END
  END data_out_right[4]
  PIN data_out_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 136.000 861.030 144.000 ;
    END
  END data_out_right[5]
  PIN data_out_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 136.000 870.230 144.000 ;
    END
  END data_out_right[6]
  PIN data_out_right[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 136.000 879.430 144.000 ;
    END
  END data_out_right[7]
  PIN data_out_right[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 136.000 888.630 144.000 ;
    END
  END data_out_right[8]
  PIN data_out_right[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 136.000 897.830 144.000 ;
    END
  END data_out_right[9]
  PIN inverter_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 136.000 1311.830 144.000 ;
    END
  END inverter_select[0]
  PIN inverter_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 136.000 1321.030 144.000 ;
    END
  END inverter_select[1]
  PIN inverter_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 136.000 1330.230 144.000 ;
    END
  END inverter_select[2]
  PIN inverter_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.150 136.000 1339.430 144.000 ;
    END
  END inverter_select[3]
  PIN inverter_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 136.000 1348.630 144.000 ;
    END
  END inverter_select[4]
  PIN inverter_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 136.000 1357.830 144.000 ;
    END
  END inverter_select[5]
  PIN inverter_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 136.000 1367.030 144.000 ;
    END
  END inverter_select[6]
  PIN inverter_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 136.000 1376.230 144.000 ;
    END
  END inverter_select[7]
  PIN inverter_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 136.000 1385.430 144.000 ;
    END
  END inverter_select[8]
  PIN inverter_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 136.000 1394.630 144.000 ;
    END
  END inverter_select[9]
  PIN io_control_trigger_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.280 4.000 29.880 ;
    END
  END io_control_trigger_in
  PIN io_control_trigger_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 34.040 4.000 34.640 ;
    END
  END io_control_trigger_oeb
  PIN io_driver_io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 38.800 4.000 39.400 ;
    END
  END io_driver_io_oeb[0]
  PIN io_driver_io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 43.560 4.000 44.160 ;
    END
  END io_driver_io_oeb[1]
  PIN io_driver_io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.320 4.000 48.920 ;
    END
  END io_driver_io_oeb[2]
  PIN io_driver_io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 53.080 4.000 53.680 ;
    END
  END io_driver_io_oeb[3]
  PIN io_driver_io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 57.840 4.000 58.440 ;
    END
  END io_driver_io_oeb[4]
  PIN io_driver_io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 62.600 4.000 63.200 ;
    END
  END io_driver_io_oeb[5]
  PIN io_driver_io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 67.360 4.000 67.960 ;
    END
  END io_driver_io_oeb[6]
  PIN io_driver_io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.120 4.000 72.720 ;
    END
  END io_driver_io_oeb[7]
  PIN io_driver_io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.880 4.000 77.480 ;
    END
  END io_driver_io_oeb[8]
  PIN io_driver_io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 81.640 4.000 82.240 ;
    END
  END io_driver_io_oeb[9]
  PIN io_latch_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 19.760 4.000 20.360 ;
    END
  END io_latch_data_in
  PIN io_latch_data_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 24.520 4.000 25.120 ;
    END
  END io_latch_data_oeb
  PIN io_miso_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 129.240 4.000 129.840 ;
    END
  END io_miso_oeb
  PIN io_miso_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 124.480 4.000 125.080 ;
    END
  END io_miso_out
  PIN io_mosi_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 105.440 4.000 106.040 ;
    END
  END io_mosi_in
  PIN io_mosi_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 110.200 4.000 110.800 ;
    END
  END io_mosi_oeb
  PIN io_reset_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.240 4.000 10.840 ;
    END
  END io_reset_n_in
  PIN io_reset_n_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 15.000 4.000 15.600 ;
    END
  END io_reset_n_oeb
  PIN io_sclk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 95.920 4.000 96.520 ;
    END
  END io_sclk_in
  PIN io_sclk_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.680 4.000 101.280 ;
    END
  END io_sclk_oeb
  PIN io_ss_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 114.960 4.000 115.560 ;
    END
  END io_ss_n_in
  PIN io_ss_n_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 119.720 4.000 120.320 ;
    END
  END io_ss_n_oeb
  PIN io_update_cycle_complete_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 91.160 4.000 91.760 ;
    END
  END io_update_cycle_complete_oeb
  PIN io_update_cycle_complete_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 86.400 4.000 87.000 ;
    END
  END io_update_cycle_complete_out
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 -4.000 54.650 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 -4.000 560.650 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 -4.000 565.710 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 -4.000 570.770 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 -4.000 575.830 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 -4.000 580.890 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 -4.000 585.950 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 -4.000 591.010 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 -4.000 596.070 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 -4.000 601.130 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 -4.000 606.190 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 -4.000 105.250 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 -4.000 611.250 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 -4.000 616.310 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 -4.000 621.370 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 -4.000 626.430 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 -4.000 631.490 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 -4.000 636.550 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 -4.000 641.610 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 -4.000 646.670 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 -4.000 651.730 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 -4.000 656.790 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 -4.000 110.310 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 -4.000 661.850 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 -4.000 666.910 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 -4.000 671.970 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 -4.000 677.030 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 -4.000 682.090 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 -4.000 687.150 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 -4.000 692.210 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 -4.000 697.270 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 -4.000 115.370 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 -4.000 120.430 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 -4.000 125.490 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 -4.000 130.550 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 -4.000 135.610 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 -4.000 140.670 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 -4.000 145.730 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 -4.000 150.790 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 -4.000 59.710 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 -4.000 155.850 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 -4.000 160.910 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 -4.000 165.970 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 -4.000 171.030 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 -4.000 176.090 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 -4.000 181.150 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -4.000 186.210 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 -4.000 191.270 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 -4.000 196.330 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 -4.000 201.390 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 -4.000 64.770 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 -4.000 206.450 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 -4.000 211.510 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 -4.000 216.570 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 -4.000 221.630 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 -4.000 226.690 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 -4.000 231.750 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 -4.000 236.810 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 -4.000 241.870 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 -4.000 246.930 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 -4.000 251.990 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 -4.000 69.830 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 -4.000 257.050 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 -4.000 262.110 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 -4.000 267.170 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 -4.000 272.230 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 -4.000 277.290 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 -4.000 282.350 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 -4.000 287.410 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 -4.000 292.470 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 -4.000 297.530 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 -4.000 302.590 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 -4.000 74.890 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 -4.000 307.650 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -4.000 312.710 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 -4.000 317.770 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 -4.000 322.830 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 -4.000 327.890 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 -4.000 332.950 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 -4.000 338.010 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 -4.000 343.070 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 -4.000 348.130 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 -4.000 353.190 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 -4.000 79.950 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 -4.000 358.250 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 -4.000 363.310 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 -4.000 368.370 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 -4.000 373.430 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 -4.000 378.490 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 -4.000 383.550 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 -4.000 388.610 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 -4.000 393.670 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 -4.000 398.730 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 -4.000 403.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 -4.000 85.010 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 -4.000 408.850 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 -4.000 413.910 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 -4.000 418.970 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 -4.000 424.030 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 -4.000 429.090 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 -4.000 434.150 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -4.000 439.210 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 -4.000 444.270 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 -4.000 449.330 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 -4.000 454.390 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 -4.000 90.070 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 -4.000 459.450 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 -4.000 464.510 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 -4.000 469.570 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 -4.000 474.630 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 -4.000 479.690 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 -4.000 484.750 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 -4.000 489.810 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 -4.000 494.870 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -4.000 499.930 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 -4.000 504.990 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 -4.000 95.130 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 -4.000 510.050 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 -4.000 515.110 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 -4.000 520.170 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 -4.000 525.230 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 -4.000 530.290 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 -4.000 535.350 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 -4.000 540.410 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 -4.000 545.470 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 -4.000 550.530 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 -4.000 555.590 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 -4.000 100.190 4.000 ;
    END
  END la_data_in[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 -4.000 702.330 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 -4.000 1208.330 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 -4.000 1213.390 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 -4.000 1218.450 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 -4.000 1223.510 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 -4.000 1228.570 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 -4.000 1233.630 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 -4.000 1238.690 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 -4.000 1243.750 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.530 -4.000 1248.810 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 -4.000 1253.870 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 -4.000 752.930 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 -4.000 1258.930 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 -4.000 1263.990 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 -4.000 1269.050 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 -4.000 1274.110 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 -4.000 1279.170 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 -4.000 1284.230 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 -4.000 1289.290 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 -4.000 1294.350 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 -4.000 1299.410 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 -4.000 1304.470 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 -4.000 757.990 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.250 -4.000 1309.530 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 -4.000 1314.590 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 -4.000 1319.650 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 -4.000 1324.710 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 -4.000 1329.770 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.550 -4.000 1334.830 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 -4.000 1339.890 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 -4.000 1344.950 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 -4.000 763.050 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 -4.000 768.110 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 -4.000 773.170 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 -4.000 778.230 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -4.000 783.290 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 -4.000 788.350 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 -4.000 793.410 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 -4.000 798.470 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 -4.000 707.390 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 -4.000 803.530 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 -4.000 808.590 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 -4.000 813.650 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 -4.000 818.710 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 -4.000 823.770 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 -4.000 828.830 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 -4.000 833.890 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 -4.000 838.950 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 -4.000 844.010 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 -4.000 849.070 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 -4.000 712.450 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 -4.000 854.130 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 -4.000 859.190 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 -4.000 864.250 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 -4.000 869.310 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 -4.000 874.370 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 -4.000 879.430 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 -4.000 884.490 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 -4.000 889.550 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 -4.000 894.610 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 -4.000 899.670 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 -4.000 717.510 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 -4.000 904.730 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 -4.000 909.790 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 -4.000 914.850 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 -4.000 919.910 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 -4.000 924.970 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 -4.000 930.030 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 -4.000 935.090 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 -4.000 940.150 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 -4.000 945.210 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 -4.000 950.270 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 -4.000 722.570 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 -4.000 955.330 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 -4.000 960.390 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 -4.000 965.450 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 -4.000 970.510 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 -4.000 975.570 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 -4.000 980.630 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 -4.000 985.690 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 -4.000 990.750 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 -4.000 995.810 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 -4.000 1000.870 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 -4.000 727.630 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 -4.000 1005.930 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 -4.000 1010.990 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 -4.000 1016.050 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 -4.000 1021.110 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 -4.000 1026.170 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 -4.000 1031.230 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 -4.000 1036.290 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 -4.000 1041.350 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 -4.000 1046.410 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 -4.000 1051.470 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 -4.000 732.690 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 -4.000 1056.530 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 -4.000 1061.590 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 -4.000 1066.650 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 -4.000 1071.710 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 -4.000 1076.770 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 -4.000 1081.830 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 -4.000 1086.890 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 -4.000 1091.950 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 -4.000 1097.010 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 -4.000 1102.070 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 -4.000 737.750 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 -4.000 1107.130 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 -4.000 1112.190 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 -4.000 1117.250 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 -4.000 1122.310 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 -4.000 1127.370 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 -4.000 1132.430 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 -4.000 1137.490 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 -4.000 1142.550 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 -4.000 1147.610 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 -4.000 1152.670 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 -4.000 742.810 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 -4.000 1157.730 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 -4.000 1162.790 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 -4.000 1167.850 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 -4.000 1172.910 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 -4.000 1177.970 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 -4.000 1183.030 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 -4.000 1188.090 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.870 -4.000 1193.150 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 -4.000 1198.210 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 -4.000 1203.270 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 -4.000 747.870 4.000 ;
    END
  END la_oenb[9]
  PIN mask_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 136.000 33.030 144.000 ;
    END
  END mask_select_left[0]
  PIN mask_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 136.000 42.230 144.000 ;
    END
  END mask_select_left[1]
  PIN mask_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 136.000 51.430 144.000 ;
    END
  END mask_select_left[2]
  PIN mask_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 136.000 5.430 144.000 ;
    END
  END mask_select_right[0]
  PIN mask_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 136.000 14.630 144.000 ;
    END
  END mask_select_right[1]
  PIN mask_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 136.000 23.830 144.000 ;
    END
  END mask_select_right[2]
  PIN mem_address_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 136.000 125.030 144.000 ;
    END
  END mem_address_left[0]
  PIN mem_address_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 136.000 134.230 144.000 ;
    END
  END mem_address_left[1]
  PIN mem_address_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 136.000 143.430 144.000 ;
    END
  END mem_address_left[2]
  PIN mem_address_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 136.000 152.630 144.000 ;
    END
  END mem_address_left[3]
  PIN mem_address_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 136.000 161.830 144.000 ;
    END
  END mem_address_left[4]
  PIN mem_address_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 136.000 171.030 144.000 ;
    END
  END mem_address_left[5]
  PIN mem_address_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 136.000 180.230 144.000 ;
    END
  END mem_address_left[6]
  PIN mem_address_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 136.000 60.630 144.000 ;
    END
  END mem_address_right[0]
  PIN mem_address_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 136.000 69.830 144.000 ;
    END
  END mem_address_right[1]
  PIN mem_address_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 136.000 79.030 144.000 ;
    END
  END mem_address_right[2]
  PIN mem_address_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 136.000 88.230 144.000 ;
    END
  END mem_address_right[3]
  PIN mem_address_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 136.000 97.430 144.000 ;
    END
  END mem_address_right[4]
  PIN mem_address_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 136.000 106.630 144.000 ;
    END
  END mem_address_right[5]
  PIN mem_address_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 136.000 115.830 144.000 ;
    END
  END mem_address_right[6]
  PIN mem_dot_write_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 136.000 281.430 144.000 ;
    END
  END mem_dot_write_n[0]
  PIN mem_dot_write_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 136.000 290.630 144.000 ;
    END
  END mem_dot_write_n[1]
  PIN mem_dot_write_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 136.000 299.830 144.000 ;
    END
  END mem_dot_write_n[2]
  PIN mem_dot_write_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 136.000 309.030 144.000 ;
    END
  END mem_dot_write_n[3]
  PIN mem_dot_write_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 136.000 318.230 144.000 ;
    END
  END mem_dot_write_n[4]
  PIN mem_dot_write_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 136.000 327.430 144.000 ;
    END
  END mem_dot_write_n[5]
  PIN mem_dot_write_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 136.000 336.630 144.000 ;
    END
  END mem_dot_write_n[6]
  PIN mem_dot_write_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 136.000 345.830 144.000 ;
    END
  END mem_dot_write_n[7]
  PIN mem_dot_write_n[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 136.000 355.030 144.000 ;
    END
  END mem_dot_write_n[8]
  PIN mem_dot_write_n[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 136.000 364.230 144.000 ;
    END
  END mem_dot_write_n[9]
  PIN mem_sel_col_address_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 136.000 750.630 144.000 ;
    END
  END mem_sel_col_address_left[0]
  PIN mem_sel_col_address_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 136.000 759.830 144.000 ;
    END
  END mem_sel_col_address_left[1]
  PIN mem_sel_col_address_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 136.000 769.030 144.000 ;
    END
  END mem_sel_col_address_left[2]
  PIN mem_sel_col_address_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 136.000 778.230 144.000 ;
    END
  END mem_sel_col_address_left[3]
  PIN mem_sel_col_address_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 136.000 787.430 144.000 ;
    END
  END mem_sel_col_address_left[4]
  PIN mem_sel_col_address_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 136.000 796.630 144.000 ;
    END
  END mem_sel_col_address_left[5]
  PIN mem_sel_col_address_left[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 136.000 805.830 144.000 ;
    END
  END mem_sel_col_address_left[6]
  PIN mem_sel_col_address_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 136.000 686.230 144.000 ;
    END
  END mem_sel_col_address_right[0]
  PIN mem_sel_col_address_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 136.000 695.430 144.000 ;
    END
  END mem_sel_col_address_right[1]
  PIN mem_sel_col_address_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 136.000 704.630 144.000 ;
    END
  END mem_sel_col_address_right[2]
  PIN mem_sel_col_address_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 136.000 713.830 144.000 ;
    END
  END mem_sel_col_address_right[3]
  PIN mem_sel_col_address_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 136.000 723.030 144.000 ;
    END
  END mem_sel_col_address_right[4]
  PIN mem_sel_col_address_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 136.000 732.230 144.000 ;
    END
  END mem_sel_col_address_right[5]
  PIN mem_sel_col_address_right[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 136.000 741.430 144.000 ;
    END
  END mem_sel_col_address_right[6]
  PIN mem_sel_write_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 136.000 1109.430 144.000 ;
    END
  END mem_sel_write_n[0]
  PIN mem_sel_write_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 136.000 1118.630 144.000 ;
    END
  END mem_sel_write_n[1]
  PIN mem_sel_write_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 136.000 1127.830 144.000 ;
    END
  END mem_sel_write_n[2]
  PIN mem_sel_write_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 136.000 1137.030 144.000 ;
    END
  END mem_sel_write_n[3]
  PIN mem_sel_write_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 136.000 1146.230 144.000 ;
    END
  END mem_sel_write_n[4]
  PIN mem_sel_write_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 136.000 1155.430 144.000 ;
    END
  END mem_sel_write_n[5]
  PIN mem_sel_write_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 136.000 1164.630 144.000 ;
    END
  END mem_sel_write_n[6]
  PIN mem_sel_write_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 136.000 1173.830 144.000 ;
    END
  END mem_sel_write_n[7]
  PIN mem_sel_write_n[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 136.000 1183.030 144.000 ;
    END
  END mem_sel_write_n[8]
  PIN mem_sel_write_n[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 136.000 1192.230 144.000 ;
    END
  END mem_sel_write_n[9]
  PIN mem_write_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 136.000 189.430 144.000 ;
    END
  END mem_write_n[0]
  PIN mem_write_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 136.000 198.630 144.000 ;
    END
  END mem_write_n[1]
  PIN mem_write_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 136.000 207.830 144.000 ;
    END
  END mem_write_n[2]
  PIN mem_write_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 136.000 217.030 144.000 ;
    END
  END mem_write_n[3]
  PIN mem_write_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 136.000 226.230 144.000 ;
    END
  END mem_write_n[4]
  PIN mem_write_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 136.000 235.430 144.000 ;
    END
  END mem_write_n[5]
  PIN mem_write_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 136.000 244.630 144.000 ;
    END
  END mem_write_n[6]
  PIN mem_write_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 136.000 253.830 144.000 ;
    END
  END mem_write_n[7]
  PIN mem_write_n[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 136.000 263.030 144.000 ;
    END
  END mem_write_n[8]
  PIN mem_write_n[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 136.000 272.230 144.000 ;
    END
  END mem_write_n[9]
  PIN output_active_left
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 136.000 1302.630 144.000 ;
    END
  END output_active_left
  PIN output_active_right
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 136.000 1293.430 144.000 ;
    END
  END output_active_right
  PIN row_col_select[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 136.000 1201.430 144.000 ;
    END
  END row_col_select[0]
  PIN row_col_select[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 136.000 1210.630 144.000 ;
    END
  END row_col_select[1]
  PIN row_col_select[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 136.000 1219.830 144.000 ;
    END
  END row_col_select[2]
  PIN row_col_select[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 136.000 1229.030 144.000 ;
    END
  END row_col_select[3]
  PIN row_col_select[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 136.000 1238.230 144.000 ;
    END
  END row_col_select[4]
  PIN row_col_select[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 136.000 1247.430 144.000 ;
    END
  END row_col_select[5]
  PIN row_col_select[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 136.000 1256.630 144.000 ;
    END
  END row_col_select[6]
  PIN row_col_select[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 136.000 1265.830 144.000 ;
    END
  END row_col_select[7]
  PIN row_col_select[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.750 136.000 1275.030 144.000 ;
    END
  END row_col_select[8]
  PIN row_col_select[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 136.000 1284.230 144.000 ;
    END
  END row_col_select[9]
  PIN row_select_left[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 136.000 428.630 144.000 ;
    END
  END row_select_left[0]
  PIN row_select_left[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 136.000 437.830 144.000 ;
    END
  END row_select_left[1]
  PIN row_select_left[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 136.000 447.030 144.000 ;
    END
  END row_select_left[2]
  PIN row_select_left[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 136.000 456.230 144.000 ;
    END
  END row_select_left[3]
  PIN row_select_left[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 136.000 465.430 144.000 ;
    END
  END row_select_left[4]
  PIN row_select_left[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 136.000 474.630 144.000 ;
    END
  END row_select_left[5]
  PIN row_select_right[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 136.000 373.430 144.000 ;
    END
  END row_select_right[0]
  PIN row_select_right[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 136.000 382.630 144.000 ;
    END
  END row_select_right[1]
  PIN row_select_right[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 136.000 391.830 144.000 ;
    END
  END row_select_right[2]
  PIN row_select_right[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 136.000 401.030 144.000 ;
    END
  END row_select_right[3]
  PIN row_select_right[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 136.000 410.230 144.000 ;
    END
  END row_select_right[4]
  PIN row_select_right[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 136.000 419.430 144.000 ;
    END
  END row_select_right[5]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 69.400 1404.000 70.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.340 10.640 624.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.340 10.640 724.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.340 10.640 824.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 919.340 10.640 924.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.340 10.640 1024.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1119.340 10.640 1124.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1219.340 10.640 1224.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1319.340 10.640 1324.340 128.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 669.340 10.640 674.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.340 10.640 774.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 869.340 10.640 874.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 969.340 10.640 974.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1069.340 10.640 1074.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1169.340 10.640 1174.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.340 10.640 1274.340 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1369.340 10.640 1374.340 128.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1394.260 127.925 ;
      LAYER met1 ;
        RECT 5.130 7.520 1394.650 130.180 ;
      LAYER met2 ;
        RECT 5.710 135.720 14.070 136.410 ;
        RECT 14.910 135.720 23.270 136.410 ;
        RECT 24.110 135.720 32.470 136.410 ;
        RECT 33.310 135.720 41.670 136.410 ;
        RECT 42.510 135.720 50.870 136.410 ;
        RECT 51.710 135.720 60.070 136.410 ;
        RECT 60.910 135.720 69.270 136.410 ;
        RECT 70.110 135.720 78.470 136.410 ;
        RECT 79.310 135.720 87.670 136.410 ;
        RECT 88.510 135.720 96.870 136.410 ;
        RECT 97.710 135.720 106.070 136.410 ;
        RECT 106.910 135.720 115.270 136.410 ;
        RECT 116.110 135.720 124.470 136.410 ;
        RECT 125.310 135.720 133.670 136.410 ;
        RECT 134.510 135.720 142.870 136.410 ;
        RECT 143.710 135.720 152.070 136.410 ;
        RECT 152.910 135.720 161.270 136.410 ;
        RECT 162.110 135.720 170.470 136.410 ;
        RECT 171.310 135.720 179.670 136.410 ;
        RECT 180.510 135.720 188.870 136.410 ;
        RECT 189.710 135.720 198.070 136.410 ;
        RECT 198.910 135.720 207.270 136.410 ;
        RECT 208.110 135.720 216.470 136.410 ;
        RECT 217.310 135.720 225.670 136.410 ;
        RECT 226.510 135.720 234.870 136.410 ;
        RECT 235.710 135.720 244.070 136.410 ;
        RECT 244.910 135.720 253.270 136.410 ;
        RECT 254.110 135.720 262.470 136.410 ;
        RECT 263.310 135.720 271.670 136.410 ;
        RECT 272.510 135.720 280.870 136.410 ;
        RECT 281.710 135.720 290.070 136.410 ;
        RECT 290.910 135.720 299.270 136.410 ;
        RECT 300.110 135.720 308.470 136.410 ;
        RECT 309.310 135.720 317.670 136.410 ;
        RECT 318.510 135.720 326.870 136.410 ;
        RECT 327.710 135.720 336.070 136.410 ;
        RECT 336.910 135.720 345.270 136.410 ;
        RECT 346.110 135.720 354.470 136.410 ;
        RECT 355.310 135.720 363.670 136.410 ;
        RECT 364.510 135.720 372.870 136.410 ;
        RECT 373.710 135.720 382.070 136.410 ;
        RECT 382.910 135.720 391.270 136.410 ;
        RECT 392.110 135.720 400.470 136.410 ;
        RECT 401.310 135.720 409.670 136.410 ;
        RECT 410.510 135.720 418.870 136.410 ;
        RECT 419.710 135.720 428.070 136.410 ;
        RECT 428.910 135.720 437.270 136.410 ;
        RECT 438.110 135.720 446.470 136.410 ;
        RECT 447.310 135.720 455.670 136.410 ;
        RECT 456.510 135.720 464.870 136.410 ;
        RECT 465.710 135.720 474.070 136.410 ;
        RECT 474.910 135.720 483.270 136.410 ;
        RECT 484.110 135.720 492.470 136.410 ;
        RECT 493.310 135.720 501.670 136.410 ;
        RECT 502.510 135.720 510.870 136.410 ;
        RECT 511.710 135.720 520.070 136.410 ;
        RECT 520.910 135.720 529.270 136.410 ;
        RECT 530.110 135.720 538.470 136.410 ;
        RECT 539.310 135.720 547.670 136.410 ;
        RECT 548.510 135.720 556.870 136.410 ;
        RECT 557.710 135.720 566.070 136.410 ;
        RECT 566.910 135.720 575.270 136.410 ;
        RECT 576.110 135.720 584.470 136.410 ;
        RECT 585.310 135.720 593.670 136.410 ;
        RECT 594.510 135.720 602.870 136.410 ;
        RECT 603.710 135.720 612.070 136.410 ;
        RECT 612.910 135.720 621.270 136.410 ;
        RECT 622.110 135.720 630.470 136.410 ;
        RECT 631.310 135.720 639.670 136.410 ;
        RECT 640.510 135.720 648.870 136.410 ;
        RECT 649.710 135.720 658.070 136.410 ;
        RECT 658.910 135.720 667.270 136.410 ;
        RECT 668.110 135.720 676.470 136.410 ;
        RECT 677.310 135.720 685.670 136.410 ;
        RECT 686.510 135.720 694.870 136.410 ;
        RECT 695.710 135.720 704.070 136.410 ;
        RECT 704.910 135.720 713.270 136.410 ;
        RECT 714.110 135.720 722.470 136.410 ;
        RECT 723.310 135.720 731.670 136.410 ;
        RECT 732.510 135.720 740.870 136.410 ;
        RECT 741.710 135.720 750.070 136.410 ;
        RECT 750.910 135.720 759.270 136.410 ;
        RECT 760.110 135.720 768.470 136.410 ;
        RECT 769.310 135.720 777.670 136.410 ;
        RECT 778.510 135.720 786.870 136.410 ;
        RECT 787.710 135.720 796.070 136.410 ;
        RECT 796.910 135.720 805.270 136.410 ;
        RECT 806.110 135.720 814.470 136.410 ;
        RECT 815.310 135.720 823.670 136.410 ;
        RECT 824.510 135.720 832.870 136.410 ;
        RECT 833.710 135.720 842.070 136.410 ;
        RECT 842.910 135.720 851.270 136.410 ;
        RECT 852.110 135.720 860.470 136.410 ;
        RECT 861.310 135.720 869.670 136.410 ;
        RECT 870.510 135.720 878.870 136.410 ;
        RECT 879.710 135.720 888.070 136.410 ;
        RECT 888.910 135.720 897.270 136.410 ;
        RECT 898.110 135.720 906.470 136.410 ;
        RECT 907.310 135.720 915.670 136.410 ;
        RECT 916.510 135.720 924.870 136.410 ;
        RECT 925.710 135.720 934.070 136.410 ;
        RECT 934.910 135.720 943.270 136.410 ;
        RECT 944.110 135.720 952.470 136.410 ;
        RECT 953.310 135.720 961.670 136.410 ;
        RECT 962.510 135.720 970.870 136.410 ;
        RECT 971.710 135.720 980.070 136.410 ;
        RECT 980.910 135.720 989.270 136.410 ;
        RECT 990.110 135.720 998.470 136.410 ;
        RECT 999.310 135.720 1007.670 136.410 ;
        RECT 1008.510 135.720 1016.870 136.410 ;
        RECT 1017.710 135.720 1026.070 136.410 ;
        RECT 1026.910 135.720 1035.270 136.410 ;
        RECT 1036.110 135.720 1044.470 136.410 ;
        RECT 1045.310 135.720 1053.670 136.410 ;
        RECT 1054.510 135.720 1062.870 136.410 ;
        RECT 1063.710 135.720 1072.070 136.410 ;
        RECT 1072.910 135.720 1081.270 136.410 ;
        RECT 1082.110 135.720 1090.470 136.410 ;
        RECT 1091.310 135.720 1099.670 136.410 ;
        RECT 1100.510 135.720 1108.870 136.410 ;
        RECT 1109.710 135.720 1118.070 136.410 ;
        RECT 1118.910 135.720 1127.270 136.410 ;
        RECT 1128.110 135.720 1136.470 136.410 ;
        RECT 1137.310 135.720 1145.670 136.410 ;
        RECT 1146.510 135.720 1154.870 136.410 ;
        RECT 1155.710 135.720 1164.070 136.410 ;
        RECT 1164.910 135.720 1173.270 136.410 ;
        RECT 1174.110 135.720 1182.470 136.410 ;
        RECT 1183.310 135.720 1191.670 136.410 ;
        RECT 1192.510 135.720 1200.870 136.410 ;
        RECT 1201.710 135.720 1210.070 136.410 ;
        RECT 1210.910 135.720 1219.270 136.410 ;
        RECT 1220.110 135.720 1228.470 136.410 ;
        RECT 1229.310 135.720 1237.670 136.410 ;
        RECT 1238.510 135.720 1246.870 136.410 ;
        RECT 1247.710 135.720 1256.070 136.410 ;
        RECT 1256.910 135.720 1265.270 136.410 ;
        RECT 1266.110 135.720 1274.470 136.410 ;
        RECT 1275.310 135.720 1283.670 136.410 ;
        RECT 1284.510 135.720 1292.870 136.410 ;
        RECT 1293.710 135.720 1302.070 136.410 ;
        RECT 1302.910 135.720 1311.270 136.410 ;
        RECT 1312.110 135.720 1320.470 136.410 ;
        RECT 1321.310 135.720 1329.670 136.410 ;
        RECT 1330.510 135.720 1338.870 136.410 ;
        RECT 1339.710 135.720 1348.070 136.410 ;
        RECT 1348.910 135.720 1357.270 136.410 ;
        RECT 1358.110 135.720 1366.470 136.410 ;
        RECT 1367.310 135.720 1375.670 136.410 ;
        RECT 1376.510 135.720 1384.870 136.410 ;
        RECT 1385.710 135.720 1394.070 136.410 ;
        RECT 5.160 4.280 1394.620 135.720 ;
        RECT 5.160 3.670 54.090 4.280 ;
        RECT 54.930 3.670 59.150 4.280 ;
        RECT 59.990 3.670 64.210 4.280 ;
        RECT 65.050 3.670 69.270 4.280 ;
        RECT 70.110 3.670 74.330 4.280 ;
        RECT 75.170 3.670 79.390 4.280 ;
        RECT 80.230 3.670 84.450 4.280 ;
        RECT 85.290 3.670 89.510 4.280 ;
        RECT 90.350 3.670 94.570 4.280 ;
        RECT 95.410 3.670 99.630 4.280 ;
        RECT 100.470 3.670 104.690 4.280 ;
        RECT 105.530 3.670 109.750 4.280 ;
        RECT 110.590 3.670 114.810 4.280 ;
        RECT 115.650 3.670 119.870 4.280 ;
        RECT 120.710 3.670 124.930 4.280 ;
        RECT 125.770 3.670 129.990 4.280 ;
        RECT 130.830 3.670 135.050 4.280 ;
        RECT 135.890 3.670 140.110 4.280 ;
        RECT 140.950 3.670 145.170 4.280 ;
        RECT 146.010 3.670 150.230 4.280 ;
        RECT 151.070 3.670 155.290 4.280 ;
        RECT 156.130 3.670 160.350 4.280 ;
        RECT 161.190 3.670 165.410 4.280 ;
        RECT 166.250 3.670 170.470 4.280 ;
        RECT 171.310 3.670 175.530 4.280 ;
        RECT 176.370 3.670 180.590 4.280 ;
        RECT 181.430 3.670 185.650 4.280 ;
        RECT 186.490 3.670 190.710 4.280 ;
        RECT 191.550 3.670 195.770 4.280 ;
        RECT 196.610 3.670 200.830 4.280 ;
        RECT 201.670 3.670 205.890 4.280 ;
        RECT 206.730 3.670 210.950 4.280 ;
        RECT 211.790 3.670 216.010 4.280 ;
        RECT 216.850 3.670 221.070 4.280 ;
        RECT 221.910 3.670 226.130 4.280 ;
        RECT 226.970 3.670 231.190 4.280 ;
        RECT 232.030 3.670 236.250 4.280 ;
        RECT 237.090 3.670 241.310 4.280 ;
        RECT 242.150 3.670 246.370 4.280 ;
        RECT 247.210 3.670 251.430 4.280 ;
        RECT 252.270 3.670 256.490 4.280 ;
        RECT 257.330 3.670 261.550 4.280 ;
        RECT 262.390 3.670 266.610 4.280 ;
        RECT 267.450 3.670 271.670 4.280 ;
        RECT 272.510 3.670 276.730 4.280 ;
        RECT 277.570 3.670 281.790 4.280 ;
        RECT 282.630 3.670 286.850 4.280 ;
        RECT 287.690 3.670 291.910 4.280 ;
        RECT 292.750 3.670 296.970 4.280 ;
        RECT 297.810 3.670 302.030 4.280 ;
        RECT 302.870 3.670 307.090 4.280 ;
        RECT 307.930 3.670 312.150 4.280 ;
        RECT 312.990 3.670 317.210 4.280 ;
        RECT 318.050 3.670 322.270 4.280 ;
        RECT 323.110 3.670 327.330 4.280 ;
        RECT 328.170 3.670 332.390 4.280 ;
        RECT 333.230 3.670 337.450 4.280 ;
        RECT 338.290 3.670 342.510 4.280 ;
        RECT 343.350 3.670 347.570 4.280 ;
        RECT 348.410 3.670 352.630 4.280 ;
        RECT 353.470 3.670 357.690 4.280 ;
        RECT 358.530 3.670 362.750 4.280 ;
        RECT 363.590 3.670 367.810 4.280 ;
        RECT 368.650 3.670 372.870 4.280 ;
        RECT 373.710 3.670 377.930 4.280 ;
        RECT 378.770 3.670 382.990 4.280 ;
        RECT 383.830 3.670 388.050 4.280 ;
        RECT 388.890 3.670 393.110 4.280 ;
        RECT 393.950 3.670 398.170 4.280 ;
        RECT 399.010 3.670 403.230 4.280 ;
        RECT 404.070 3.670 408.290 4.280 ;
        RECT 409.130 3.670 413.350 4.280 ;
        RECT 414.190 3.670 418.410 4.280 ;
        RECT 419.250 3.670 423.470 4.280 ;
        RECT 424.310 3.670 428.530 4.280 ;
        RECT 429.370 3.670 433.590 4.280 ;
        RECT 434.430 3.670 438.650 4.280 ;
        RECT 439.490 3.670 443.710 4.280 ;
        RECT 444.550 3.670 448.770 4.280 ;
        RECT 449.610 3.670 453.830 4.280 ;
        RECT 454.670 3.670 458.890 4.280 ;
        RECT 459.730 3.670 463.950 4.280 ;
        RECT 464.790 3.670 469.010 4.280 ;
        RECT 469.850 3.670 474.070 4.280 ;
        RECT 474.910 3.670 479.130 4.280 ;
        RECT 479.970 3.670 484.190 4.280 ;
        RECT 485.030 3.670 489.250 4.280 ;
        RECT 490.090 3.670 494.310 4.280 ;
        RECT 495.150 3.670 499.370 4.280 ;
        RECT 500.210 3.670 504.430 4.280 ;
        RECT 505.270 3.670 509.490 4.280 ;
        RECT 510.330 3.670 514.550 4.280 ;
        RECT 515.390 3.670 519.610 4.280 ;
        RECT 520.450 3.670 524.670 4.280 ;
        RECT 525.510 3.670 529.730 4.280 ;
        RECT 530.570 3.670 534.790 4.280 ;
        RECT 535.630 3.670 539.850 4.280 ;
        RECT 540.690 3.670 544.910 4.280 ;
        RECT 545.750 3.670 549.970 4.280 ;
        RECT 550.810 3.670 555.030 4.280 ;
        RECT 555.870 3.670 560.090 4.280 ;
        RECT 560.930 3.670 565.150 4.280 ;
        RECT 565.990 3.670 570.210 4.280 ;
        RECT 571.050 3.670 575.270 4.280 ;
        RECT 576.110 3.670 580.330 4.280 ;
        RECT 581.170 3.670 585.390 4.280 ;
        RECT 586.230 3.670 590.450 4.280 ;
        RECT 591.290 3.670 595.510 4.280 ;
        RECT 596.350 3.670 600.570 4.280 ;
        RECT 601.410 3.670 605.630 4.280 ;
        RECT 606.470 3.670 610.690 4.280 ;
        RECT 611.530 3.670 615.750 4.280 ;
        RECT 616.590 3.670 620.810 4.280 ;
        RECT 621.650 3.670 625.870 4.280 ;
        RECT 626.710 3.670 630.930 4.280 ;
        RECT 631.770 3.670 635.990 4.280 ;
        RECT 636.830 3.670 641.050 4.280 ;
        RECT 641.890 3.670 646.110 4.280 ;
        RECT 646.950 3.670 651.170 4.280 ;
        RECT 652.010 3.670 656.230 4.280 ;
        RECT 657.070 3.670 661.290 4.280 ;
        RECT 662.130 3.670 666.350 4.280 ;
        RECT 667.190 3.670 671.410 4.280 ;
        RECT 672.250 3.670 676.470 4.280 ;
        RECT 677.310 3.670 681.530 4.280 ;
        RECT 682.370 3.670 686.590 4.280 ;
        RECT 687.430 3.670 691.650 4.280 ;
        RECT 692.490 3.670 696.710 4.280 ;
        RECT 697.550 3.670 701.770 4.280 ;
        RECT 702.610 3.670 706.830 4.280 ;
        RECT 707.670 3.670 711.890 4.280 ;
        RECT 712.730 3.670 716.950 4.280 ;
        RECT 717.790 3.670 722.010 4.280 ;
        RECT 722.850 3.670 727.070 4.280 ;
        RECT 727.910 3.670 732.130 4.280 ;
        RECT 732.970 3.670 737.190 4.280 ;
        RECT 738.030 3.670 742.250 4.280 ;
        RECT 743.090 3.670 747.310 4.280 ;
        RECT 748.150 3.670 752.370 4.280 ;
        RECT 753.210 3.670 757.430 4.280 ;
        RECT 758.270 3.670 762.490 4.280 ;
        RECT 763.330 3.670 767.550 4.280 ;
        RECT 768.390 3.670 772.610 4.280 ;
        RECT 773.450 3.670 777.670 4.280 ;
        RECT 778.510 3.670 782.730 4.280 ;
        RECT 783.570 3.670 787.790 4.280 ;
        RECT 788.630 3.670 792.850 4.280 ;
        RECT 793.690 3.670 797.910 4.280 ;
        RECT 798.750 3.670 802.970 4.280 ;
        RECT 803.810 3.670 808.030 4.280 ;
        RECT 808.870 3.670 813.090 4.280 ;
        RECT 813.930 3.670 818.150 4.280 ;
        RECT 818.990 3.670 823.210 4.280 ;
        RECT 824.050 3.670 828.270 4.280 ;
        RECT 829.110 3.670 833.330 4.280 ;
        RECT 834.170 3.670 838.390 4.280 ;
        RECT 839.230 3.670 843.450 4.280 ;
        RECT 844.290 3.670 848.510 4.280 ;
        RECT 849.350 3.670 853.570 4.280 ;
        RECT 854.410 3.670 858.630 4.280 ;
        RECT 859.470 3.670 863.690 4.280 ;
        RECT 864.530 3.670 868.750 4.280 ;
        RECT 869.590 3.670 873.810 4.280 ;
        RECT 874.650 3.670 878.870 4.280 ;
        RECT 879.710 3.670 883.930 4.280 ;
        RECT 884.770 3.670 888.990 4.280 ;
        RECT 889.830 3.670 894.050 4.280 ;
        RECT 894.890 3.670 899.110 4.280 ;
        RECT 899.950 3.670 904.170 4.280 ;
        RECT 905.010 3.670 909.230 4.280 ;
        RECT 910.070 3.670 914.290 4.280 ;
        RECT 915.130 3.670 919.350 4.280 ;
        RECT 920.190 3.670 924.410 4.280 ;
        RECT 925.250 3.670 929.470 4.280 ;
        RECT 930.310 3.670 934.530 4.280 ;
        RECT 935.370 3.670 939.590 4.280 ;
        RECT 940.430 3.670 944.650 4.280 ;
        RECT 945.490 3.670 949.710 4.280 ;
        RECT 950.550 3.670 954.770 4.280 ;
        RECT 955.610 3.670 959.830 4.280 ;
        RECT 960.670 3.670 964.890 4.280 ;
        RECT 965.730 3.670 969.950 4.280 ;
        RECT 970.790 3.670 975.010 4.280 ;
        RECT 975.850 3.670 980.070 4.280 ;
        RECT 980.910 3.670 985.130 4.280 ;
        RECT 985.970 3.670 990.190 4.280 ;
        RECT 991.030 3.670 995.250 4.280 ;
        RECT 996.090 3.670 1000.310 4.280 ;
        RECT 1001.150 3.670 1005.370 4.280 ;
        RECT 1006.210 3.670 1010.430 4.280 ;
        RECT 1011.270 3.670 1015.490 4.280 ;
        RECT 1016.330 3.670 1020.550 4.280 ;
        RECT 1021.390 3.670 1025.610 4.280 ;
        RECT 1026.450 3.670 1030.670 4.280 ;
        RECT 1031.510 3.670 1035.730 4.280 ;
        RECT 1036.570 3.670 1040.790 4.280 ;
        RECT 1041.630 3.670 1045.850 4.280 ;
        RECT 1046.690 3.670 1050.910 4.280 ;
        RECT 1051.750 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1061.030 4.280 ;
        RECT 1061.870 3.670 1066.090 4.280 ;
        RECT 1066.930 3.670 1071.150 4.280 ;
        RECT 1071.990 3.670 1076.210 4.280 ;
        RECT 1077.050 3.670 1081.270 4.280 ;
        RECT 1082.110 3.670 1086.330 4.280 ;
        RECT 1087.170 3.670 1091.390 4.280 ;
        RECT 1092.230 3.670 1096.450 4.280 ;
        RECT 1097.290 3.670 1101.510 4.280 ;
        RECT 1102.350 3.670 1106.570 4.280 ;
        RECT 1107.410 3.670 1111.630 4.280 ;
        RECT 1112.470 3.670 1116.690 4.280 ;
        RECT 1117.530 3.670 1121.750 4.280 ;
        RECT 1122.590 3.670 1126.810 4.280 ;
        RECT 1127.650 3.670 1131.870 4.280 ;
        RECT 1132.710 3.670 1136.930 4.280 ;
        RECT 1137.770 3.670 1141.990 4.280 ;
        RECT 1142.830 3.670 1147.050 4.280 ;
        RECT 1147.890 3.670 1152.110 4.280 ;
        RECT 1152.950 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1167.290 4.280 ;
        RECT 1168.130 3.670 1172.350 4.280 ;
        RECT 1173.190 3.670 1177.410 4.280 ;
        RECT 1178.250 3.670 1182.470 4.280 ;
        RECT 1183.310 3.670 1187.530 4.280 ;
        RECT 1188.370 3.670 1192.590 4.280 ;
        RECT 1193.430 3.670 1197.650 4.280 ;
        RECT 1198.490 3.670 1202.710 4.280 ;
        RECT 1203.550 3.670 1207.770 4.280 ;
        RECT 1208.610 3.670 1212.830 4.280 ;
        RECT 1213.670 3.670 1217.890 4.280 ;
        RECT 1218.730 3.670 1222.950 4.280 ;
        RECT 1223.790 3.670 1228.010 4.280 ;
        RECT 1228.850 3.670 1233.070 4.280 ;
        RECT 1233.910 3.670 1238.130 4.280 ;
        RECT 1238.970 3.670 1243.190 4.280 ;
        RECT 1244.030 3.670 1248.250 4.280 ;
        RECT 1249.090 3.670 1253.310 4.280 ;
        RECT 1254.150 3.670 1258.370 4.280 ;
        RECT 1259.210 3.670 1263.430 4.280 ;
        RECT 1264.270 3.670 1268.490 4.280 ;
        RECT 1269.330 3.670 1273.550 4.280 ;
        RECT 1274.390 3.670 1278.610 4.280 ;
        RECT 1279.450 3.670 1283.670 4.280 ;
        RECT 1284.510 3.670 1288.730 4.280 ;
        RECT 1289.570 3.670 1293.790 4.280 ;
        RECT 1294.630 3.670 1298.850 4.280 ;
        RECT 1299.690 3.670 1303.910 4.280 ;
        RECT 1304.750 3.670 1308.970 4.280 ;
        RECT 1309.810 3.670 1314.030 4.280 ;
        RECT 1314.870 3.670 1319.090 4.280 ;
        RECT 1319.930 3.670 1324.150 4.280 ;
        RECT 1324.990 3.670 1329.210 4.280 ;
        RECT 1330.050 3.670 1334.270 4.280 ;
        RECT 1335.110 3.670 1339.330 4.280 ;
        RECT 1340.170 3.670 1344.390 4.280 ;
        RECT 1345.230 3.670 1394.620 4.280 ;
      LAYER met3 ;
        RECT 4.400 128.840 1396.000 129.705 ;
        RECT 4.000 125.480 1396.000 128.840 ;
        RECT 4.400 124.080 1396.000 125.480 ;
        RECT 4.000 120.720 1396.000 124.080 ;
        RECT 4.400 119.320 1396.000 120.720 ;
        RECT 4.000 115.960 1396.000 119.320 ;
        RECT 4.400 114.560 1396.000 115.960 ;
        RECT 4.000 111.200 1396.000 114.560 ;
        RECT 4.400 109.800 1396.000 111.200 ;
        RECT 4.000 106.440 1396.000 109.800 ;
        RECT 4.400 105.040 1396.000 106.440 ;
        RECT 4.000 101.680 1396.000 105.040 ;
        RECT 4.400 100.280 1396.000 101.680 ;
        RECT 4.000 96.920 1396.000 100.280 ;
        RECT 4.400 95.520 1396.000 96.920 ;
        RECT 4.000 92.160 1396.000 95.520 ;
        RECT 4.400 90.760 1396.000 92.160 ;
        RECT 4.000 87.400 1396.000 90.760 ;
        RECT 4.400 86.000 1396.000 87.400 ;
        RECT 4.000 82.640 1396.000 86.000 ;
        RECT 4.400 81.240 1396.000 82.640 ;
        RECT 4.000 77.880 1396.000 81.240 ;
        RECT 4.400 76.480 1396.000 77.880 ;
        RECT 4.000 73.120 1396.000 76.480 ;
        RECT 4.400 71.720 1396.000 73.120 ;
        RECT 4.000 70.400 1396.000 71.720 ;
        RECT 4.000 69.000 1395.600 70.400 ;
        RECT 4.000 68.360 1396.000 69.000 ;
        RECT 4.400 66.960 1396.000 68.360 ;
        RECT 4.000 63.600 1396.000 66.960 ;
        RECT 4.400 62.200 1396.000 63.600 ;
        RECT 4.000 58.840 1396.000 62.200 ;
        RECT 4.400 57.440 1396.000 58.840 ;
        RECT 4.000 54.080 1396.000 57.440 ;
        RECT 4.400 52.680 1396.000 54.080 ;
        RECT 4.000 49.320 1396.000 52.680 ;
        RECT 4.400 47.920 1396.000 49.320 ;
        RECT 4.000 44.560 1396.000 47.920 ;
        RECT 4.400 43.160 1396.000 44.560 ;
        RECT 4.000 39.800 1396.000 43.160 ;
        RECT 4.400 38.400 1396.000 39.800 ;
        RECT 4.000 35.040 1396.000 38.400 ;
        RECT 4.400 33.640 1396.000 35.040 ;
        RECT 4.000 30.280 1396.000 33.640 ;
        RECT 4.400 28.880 1396.000 30.280 ;
        RECT 4.000 25.520 1396.000 28.880 ;
        RECT 4.400 24.120 1396.000 25.520 ;
        RECT 4.000 20.760 1396.000 24.120 ;
        RECT 4.400 19.360 1396.000 20.760 ;
        RECT 4.000 16.000 1396.000 19.360 ;
        RECT 4.400 14.600 1396.000 16.000 ;
        RECT 4.000 11.240 1396.000 14.600 ;
        RECT 4.400 9.840 1396.000 11.240 ;
        RECT 4.000 8.335 1396.000 9.840 ;
      LAYER met4 ;
        RECT 915.695 96.735 917.865 100.465 ;
  END
END controller_unit
END LIBRARY

