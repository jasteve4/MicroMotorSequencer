magic
tech sky130B
magscale 1 2
timestamp 1661137255
<< metal1 >>
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 19242 700992 19248 701004
rect 8168 700964 19248 700992
rect 8168 700952 8174 700964
rect 19242 700952 19248 700964
rect 19300 700992 19306 701004
rect 72970 700992 72976 701004
rect 19300 700964 72976 700992
rect 19300 700952 19306 700964
rect 72970 700952 72976 700964
rect 73028 700952 73034 701004
rect 397454 700952 397460 701004
rect 397512 700992 397518 701004
rect 462314 700992 462320 701004
rect 397512 700964 462320 700992
rect 397512 700952 397518 700964
rect 462314 700952 462320 700964
rect 462372 700952 462378 701004
rect 22002 700340 22008 700392
rect 22060 700380 22066 700392
rect 89162 700380 89168 700392
rect 22060 700352 89168 700380
rect 22060 700340 22066 700352
rect 89162 700340 89168 700352
rect 89220 700340 89226 700392
rect 138014 700340 138020 700392
rect 138072 700380 138078 700392
rect 202782 700380 202788 700392
rect 138072 700352 202788 700380
rect 138072 700340 138078 700352
rect 202782 700340 202788 700352
rect 202840 700340 202846 700392
rect 21910 700272 21916 700324
rect 21968 700312 21974 700324
rect 218974 700312 218980 700324
rect 21968 700284 218980 700312
rect 21968 700272 21974 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 302142 700272 302148 700324
rect 302200 700312 302206 700324
rect 478506 700312 478512 700324
rect 302200 700284 478512 700312
rect 302200 700272 302206 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 543458 700312 543464 700324
rect 527232 700284 543464 700312
rect 527232 700272 527238 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 22094 699660 22100 699712
rect 22152 699700 22158 699712
rect 24302 699700 24308 699712
rect 22152 699672 24308 699700
rect 22152 699660 22158 699672
rect 24302 699660 24308 699672
rect 24360 699660 24366 699712
rect 302234 698912 302240 698964
rect 302292 698952 302298 698964
rect 413646 698952 413652 698964
rect 302292 698924 413652 698952
rect 302292 698912 302298 698924
rect 413646 698912 413652 698924
rect 413704 698912 413710 698964
rect 527266 698232 527272 698284
rect 527324 698272 527330 698284
rect 580166 698272 580172 698284
rect 527324 698244 580172 698272
rect 527324 698232 527330 698244
rect 580166 698232 580172 698244
rect 580224 698232 580230 698284
rect 16482 697620 16488 697672
rect 16540 697660 16546 697672
rect 138014 697660 138020 697672
rect 16540 697632 138020 697660
rect 16540 697620 16546 697632
rect 138014 697620 138020 697632
rect 138072 697620 138078 697672
rect 22186 697552 22192 697604
rect 22244 697592 22250 697604
rect 154114 697592 154120 697604
rect 22244 697564 154120 697592
rect 22244 697552 22250 697564
rect 154114 697552 154120 697564
rect 154172 697552 154178 697604
rect 2774 606432 2780 606484
rect 2832 606472 2838 606484
rect 15838 606472 15844 606484
rect 2832 606444 15844 606472
rect 2832 606432 2838 606444
rect 15838 606432 15844 606444
rect 15896 606432 15902 606484
rect 21910 586440 21916 586492
rect 21968 586480 21974 586492
rect 28166 586480 28172 586492
rect 21968 586452 28172 586480
rect 21968 586440 21974 586452
rect 28166 586440 28172 586452
rect 28224 586440 28230 586492
rect 144822 586440 144828 586492
rect 144880 586480 144886 586492
rect 149974 586480 149980 586492
rect 144880 586452 149980 586480
rect 144880 586440 144886 586452
rect 149974 586440 149980 586452
rect 150032 586440 150038 586492
rect 302142 586440 302148 586492
rect 302200 586480 302206 586492
rect 308490 586480 308496 586492
rect 302200 586452 308496 586480
rect 302200 586440 302206 586452
rect 308490 586440 308496 586452
rect 308548 586440 308554 586492
rect 424870 586440 424876 586492
rect 424928 586480 424934 586492
rect 429930 586480 429936 586492
rect 424928 586452 429936 586480
rect 424928 586440 424934 586452
rect 429930 586440 429936 586452
rect 429988 586440 429994 586492
rect 21818 586100 21824 586152
rect 21876 586140 21882 586152
rect 43346 586140 43352 586152
rect 21876 586112 43352 586140
rect 21876 586100 21882 586112
rect 43346 586100 43352 586112
rect 43404 586100 43410 586152
rect 23290 586032 23296 586084
rect 23348 586072 23354 586084
rect 48498 586072 48504 586084
rect 23348 586044 48504 586072
rect 23348 586032 23354 586044
rect 48498 586032 48504 586044
rect 48556 586032 48562 586084
rect 266262 586032 266268 586084
rect 266320 586072 266326 586084
rect 289998 586072 290004 586084
rect 266320 586044 290004 586072
rect 266320 586032 266326 586044
rect 289998 586032 290004 586044
rect 290056 586032 290062 586084
rect 302050 586032 302056 586084
rect 302108 586072 302114 586084
rect 313550 586072 313556 586084
rect 302108 586044 313556 586072
rect 302108 586032 302114 586044
rect 313550 586032 313556 586044
rect 313608 586032 313614 586084
rect 546310 586032 546316 586084
rect 546368 586072 546374 586084
rect 568850 586072 568856 586084
rect 546368 586044 568856 586072
rect 546368 586032 546374 586044
rect 568850 586032 568856 586044
rect 568908 586032 568914 586084
rect 21726 585964 21732 586016
rect 21784 586004 21790 586016
rect 53466 586004 53472 586016
rect 21784 585976 53472 586004
rect 21784 585964 21790 585976
rect 53466 585964 53472 585976
rect 53524 585964 53530 586016
rect 261570 585964 261576 586016
rect 261628 586004 261634 586016
rect 289906 586004 289912 586016
rect 261628 585976 289912 586004
rect 261628 585964 261634 585976
rect 289906 585964 289912 585976
rect 289964 585964 289970 586016
rect 301866 585964 301872 586016
rect 301924 586004 301930 586016
rect 318610 586004 318616 586016
rect 301924 585976 318616 586004
rect 301924 585964 301930 585976
rect 318610 585964 318616 585976
rect 318668 585964 318674 586016
rect 541250 585964 541256 586016
rect 541308 586004 541314 586016
rect 567470 586004 567476 586016
rect 541308 585976 567476 586004
rect 541308 585964 541314 585976
rect 567470 585964 567476 585976
rect 567528 585964 567534 586016
rect 29638 585896 29644 585948
rect 29696 585936 29702 585948
rect 104066 585936 104072 585948
rect 29696 585908 104072 585936
rect 29696 585896 29702 585908
rect 104066 585896 104072 585908
rect 104124 585896 104130 585948
rect 256510 585896 256516 585948
rect 256568 585936 256574 585948
rect 288526 585936 288532 585948
rect 256568 585908 288532 585936
rect 256568 585896 256574 585908
rect 288526 585896 288532 585908
rect 288584 585896 288590 585948
rect 303154 585896 303160 585948
rect 303212 585936 303218 585948
rect 323670 585936 323676 585948
rect 303212 585908 323676 585936
rect 303212 585896 303218 585908
rect 323670 585896 323676 585908
rect 323728 585896 323734 585948
rect 536190 585896 536196 585948
rect 536248 585936 536254 585948
rect 568666 585936 568672 585948
rect 536248 585908 568672 585936
rect 536248 585896 536254 585908
rect 568666 585896 568672 585908
rect 568724 585896 568730 585948
rect 21910 585828 21916 585880
rect 21968 585868 21974 585880
rect 33226 585868 33232 585880
rect 21968 585840 33232 585868
rect 21968 585828 21974 585840
rect 33226 585828 33232 585840
rect 33284 585828 33290 585880
rect 35158 585828 35164 585880
rect 35216 585868 35222 585880
rect 119246 585868 119252 585880
rect 35216 585840 119252 585868
rect 35216 585828 35222 585840
rect 119246 585828 119252 585840
rect 119304 585828 119310 585880
rect 251082 585828 251088 585880
rect 251140 585868 251146 585880
rect 289814 585868 289820 585880
rect 251140 585840 289820 585868
rect 251140 585828 251146 585840
rect 289814 585828 289820 585840
rect 289872 585828 289878 585880
rect 302142 585828 302148 585880
rect 302200 585868 302206 585880
rect 328730 585868 328736 585880
rect 302200 585840 328736 585868
rect 302200 585828 302206 585840
rect 328730 585828 328736 585840
rect 328788 585828 328794 585880
rect 531130 585828 531136 585880
rect 531188 585868 531194 585880
rect 569954 585868 569960 585880
rect 531188 585840 569960 585868
rect 531188 585828 531194 585840
rect 569954 585828 569960 585840
rect 570012 585828 570018 585880
rect 23106 585760 23112 585812
rect 23164 585800 23170 585812
rect 38286 585800 38292 585812
rect 23164 585772 38292 585800
rect 23164 585760 23170 585772
rect 38286 585760 38292 585772
rect 38344 585760 38350 585812
rect 39298 585760 39304 585812
rect 39356 585800 39362 585812
rect 124306 585800 124312 585812
rect 39356 585772 124312 585800
rect 39356 585760 39362 585772
rect 124306 585760 124312 585772
rect 124364 585760 124370 585812
rect 241330 585760 241336 585812
rect 241388 585800 241394 585812
rect 287606 585800 287612 585812
rect 241388 585772 287612 585800
rect 241388 585760 241394 585772
rect 287606 585760 287612 585772
rect 287664 585760 287670 585812
rect 303246 585760 303252 585812
rect 303304 585800 303310 585812
rect 333790 585800 333796 585812
rect 303304 585772 333796 585800
rect 303304 585760 303310 585772
rect 333790 585760 333796 585772
rect 333848 585760 333854 585812
rect 521010 585760 521016 585812
rect 521068 585800 521074 585812
rect 567562 585800 567568 585812
rect 521068 585772 567568 585800
rect 521068 585760 521074 585772
rect 567562 585760 567568 585772
rect 567620 585760 567626 585812
rect 281442 585148 281448 585200
rect 281500 585188 281506 585200
rect 288618 585188 288624 585200
rect 281500 585160 288624 585188
rect 281500 585148 281506 585160
rect 288618 585148 288624 585160
rect 288676 585148 288682 585200
rect 424318 585148 424324 585200
rect 424376 585188 424382 585200
rect 424870 585188 424876 585200
rect 424376 585160 424876 585188
rect 424376 585148 424382 585160
rect 424870 585148 424876 585160
rect 424928 585148 424934 585200
rect 561490 585148 561496 585200
rect 561548 585188 561554 585200
rect 568758 585188 568764 585200
rect 561548 585160 568764 585188
rect 561548 585148 561554 585160
rect 568758 585148 568764 585160
rect 568816 585148 568822 585200
rect 300670 583312 300676 583364
rect 300728 583352 300734 583364
rect 338850 583352 338856 583364
rect 300728 583324 338856 583352
rect 300728 583312 300734 583324
rect 338850 583312 338856 583324
rect 338908 583312 338914 583364
rect 17862 583244 17868 583296
rect 17920 583284 17926 583296
rect 93946 583284 93952 583296
rect 17920 583256 93952 583284
rect 17920 583244 17926 583256
rect 93946 583244 93952 583256
rect 94004 583244 94010 583296
rect 235902 583244 235908 583296
rect 235960 583284 235966 583296
rect 292574 583284 292580 583296
rect 235960 583256 292580 583284
rect 235960 583244 235966 583256
rect 292574 583244 292580 583256
rect 292632 583244 292638 583296
rect 300486 583244 300492 583296
rect 300544 583284 300550 583296
rect 343910 583284 343916 583296
rect 300544 583256 343916 583284
rect 300544 583244 300550 583256
rect 343910 583244 343916 583256
rect 343968 583244 343974 583296
rect 17770 583176 17776 583228
rect 17828 583216 17834 583228
rect 99006 583216 99012 583228
rect 17828 583188 99012 583216
rect 17828 583176 17834 583188
rect 99006 583176 99012 583188
rect 99064 583176 99070 583228
rect 231210 583176 231216 583228
rect 231268 583216 231274 583228
rect 288802 583216 288808 583228
rect 231268 583188 288808 583216
rect 231268 583176 231274 583188
rect 288802 583176 288808 583188
rect 288860 583176 288866 583228
rect 300762 583176 300768 583228
rect 300820 583216 300826 583228
rect 348970 583216 348976 583228
rect 300820 583188 348976 583216
rect 300820 583176 300826 583188
rect 348970 583176 348976 583188
rect 349028 583176 349034 583228
rect 515950 583176 515956 583228
rect 516008 583216 516014 583228
rect 570322 583216 570328 583228
rect 516008 583188 570328 583216
rect 516008 583176 516014 583188
rect 570322 583176 570328 583188
rect 570380 583176 570386 583228
rect 15102 583108 15108 583160
rect 15160 583148 15166 583160
rect 114186 583148 114192 583160
rect 15160 583120 114192 583148
rect 15160 583108 15166 583120
rect 114186 583108 114192 583120
rect 114244 583108 114250 583160
rect 220722 583108 220728 583160
rect 220780 583148 220786 583160
rect 291470 583148 291476 583160
rect 220780 583120 291476 583148
rect 220780 583108 220786 583120
rect 291470 583108 291476 583120
rect 291528 583108 291534 583160
rect 299290 583108 299296 583160
rect 299348 583148 299354 583160
rect 354030 583148 354036 583160
rect 299348 583120 354036 583148
rect 299348 583108 299354 583120
rect 354030 583108 354036 583120
rect 354088 583108 354094 583160
rect 510890 583108 510896 583160
rect 510948 583148 510954 583160
rect 570138 583148 570144 583160
rect 510948 583120 570144 583148
rect 510948 583108 510954 583120
rect 570138 583108 570144 583120
rect 570196 583108 570202 583160
rect 15010 583040 15016 583092
rect 15068 583080 15074 583092
rect 139486 583080 139492 583092
rect 15068 583052 139492 583080
rect 15068 583040 15074 583052
rect 139486 583040 139492 583052
rect 139544 583040 139550 583092
rect 216030 583040 216036 583092
rect 216088 583080 216094 583092
rect 291194 583080 291200 583092
rect 216088 583052 291200 583080
rect 216088 583040 216094 583052
rect 291194 583040 291200 583052
rect 291252 583040 291258 583092
rect 300578 583040 300584 583092
rect 300636 583080 300642 583092
rect 359090 583080 359096 583092
rect 300636 583052 359096 583080
rect 300636 583040 300642 583052
rect 359090 583040 359096 583052
rect 359148 583040 359154 583092
rect 500770 583040 500776 583092
rect 500828 583080 500834 583092
rect 568942 583080 568948 583092
rect 500828 583052 568948 583080
rect 500828 583040 500834 583052
rect 568942 583040 568948 583052
rect 569000 583040 569006 583092
rect 19150 582972 19156 583024
rect 19208 583012 19214 583024
rect 154758 583012 154764 583024
rect 19208 582984 154764 583012
rect 19208 582972 19214 582984
rect 154758 582972 154764 582984
rect 154816 582972 154822 583024
rect 200850 582972 200856 583024
rect 200908 583012 200914 583024
rect 293218 583012 293224 583024
rect 200908 582984 293224 583012
rect 200908 582972 200914 582984
rect 293218 582972 293224 582984
rect 293276 582972 293282 583024
rect 301958 582972 301964 583024
rect 302016 583012 302022 583024
rect 364150 583012 364156 583024
rect 302016 582984 364156 583012
rect 302016 582972 302022 582984
rect 364150 582972 364156 582984
rect 364208 582972 364214 583024
rect 465350 582972 465356 583024
rect 465408 583012 465414 583024
rect 567654 583012 567660 583024
rect 465408 582984 567660 583012
rect 465408 582972 465414 582984
rect 567654 582972 567660 582984
rect 567712 582972 567718 583024
rect 195790 580524 195796 580576
rect 195848 580564 195854 580576
rect 295334 580564 295340 580576
rect 195848 580536 295340 580564
rect 195848 580524 195854 580536
rect 295334 580524 295340 580536
rect 295392 580524 295398 580576
rect 299198 580524 299204 580576
rect 299256 580564 299262 580576
rect 374270 580564 374276 580576
rect 299256 580536 374276 580564
rect 299256 580524 299262 580536
rect 374270 580524 374276 580536
rect 374328 580524 374334 580576
rect 185670 580456 185676 580508
rect 185728 580496 185734 580508
rect 287790 580496 287796 580508
rect 185728 580468 287796 580496
rect 185728 580456 185734 580468
rect 287790 580456 287796 580468
rect 287848 580456 287854 580508
rect 302970 580456 302976 580508
rect 303028 580496 303034 580508
rect 379330 580496 379336 580508
rect 303028 580468 379336 580496
rect 303028 580456 303034 580468
rect 379330 580456 379336 580468
rect 379388 580456 379394 580508
rect 190362 580388 190368 580440
rect 190420 580428 190426 580440
rect 291838 580428 291844 580440
rect 190420 580400 291844 580428
rect 190420 580388 190426 580400
rect 291838 580388 291844 580400
rect 291896 580388 291902 580440
rect 295150 580388 295156 580440
rect 295208 580428 295214 580440
rect 394510 580428 394516 580440
rect 295208 580400 394516 580428
rect 295208 580388 295214 580400
rect 394510 580388 394516 580400
rect 394568 580388 394574 580440
rect 475470 580388 475476 580440
rect 475528 580428 475534 580440
rect 574186 580428 574192 580440
rect 475528 580400 574192 580428
rect 475528 580388 475534 580400
rect 574186 580388 574192 580400
rect 574244 580388 574250 580440
rect 180610 580320 180616 580372
rect 180668 580360 180674 580372
rect 295426 580360 295432 580372
rect 180668 580332 295432 580360
rect 180668 580320 180674 580332
rect 295426 580320 295432 580332
rect 295484 580320 295490 580372
rect 297818 580320 297824 580372
rect 297876 580360 297882 580372
rect 384390 580360 384396 580372
rect 297876 580332 384396 580360
rect 297876 580320 297882 580332
rect 384390 580320 384396 580332
rect 384448 580320 384454 580372
rect 460290 580320 460296 580372
rect 460348 580360 460354 580372
rect 572714 580360 572720 580372
rect 460348 580332 572720 580360
rect 460348 580320 460354 580332
rect 572714 580320 572720 580332
rect 572772 580320 572778 580372
rect 165430 580252 165436 580304
rect 165488 580292 165494 580304
rect 295518 580292 295524 580304
rect 165488 580264 295524 580292
rect 165488 580252 165494 580264
rect 295518 580252 295524 580264
rect 295576 580252 295582 580304
rect 299382 580252 299388 580304
rect 299440 580292 299446 580304
rect 399570 580292 399576 580304
rect 299440 580264 399576 580292
rect 299440 580252 299446 580264
rect 399570 580252 399576 580264
rect 399628 580252 399634 580304
rect 455230 580252 455236 580304
rect 455288 580292 455294 580304
rect 571426 580292 571432 580304
rect 455288 580264 571432 580292
rect 455288 580252 455294 580264
rect 571426 580252 571432 580264
rect 571484 580252 571490 580304
rect 299106 577600 299112 577652
rect 299164 577640 299170 577652
rect 408494 577640 408500 577652
rect 299164 577612 408500 577640
rect 299164 577600 299170 577612
rect 408494 577600 408500 577612
rect 408552 577600 408558 577652
rect 297910 577532 297916 577584
rect 297968 577572 297974 577584
rect 414014 577572 414020 577584
rect 297968 577544 414020 577572
rect 297968 577532 297974 577544
rect 414014 577532 414020 577544
rect 414072 577532 414078 577584
rect 169754 577464 169760 577516
rect 169812 577504 169818 577516
rect 292666 577504 292672 577516
rect 169812 577476 292672 577504
rect 169812 577464 169818 577476
rect 292666 577464 292672 577476
rect 292724 577464 292730 577516
rect 295242 577464 295248 577516
rect 295300 577504 295306 577516
rect 419534 577504 419540 577516
rect 295300 577476 419540 577504
rect 295300 577464 295306 577476
rect 419534 577464 419540 577476
rect 419592 577464 419598 577516
rect 17678 574812 17684 574864
rect 17736 574852 17742 574864
rect 35158 574852 35164 574864
rect 17736 574824 35164 574852
rect 17736 574812 17742 574824
rect 35158 574812 35164 574824
rect 35216 574812 35222 574864
rect 13722 574744 13728 574796
rect 13780 574784 13786 574796
rect 128354 574784 128360 574796
rect 13780 574756 128360 574784
rect 13780 574744 13786 574756
rect 128354 574744 128360 574756
rect 128412 574744 128418 574796
rect 16390 572296 16396 572348
rect 16448 572336 16454 572348
rect 29638 572336 29644 572348
rect 16448 572308 29644 572336
rect 16448 572296 16454 572308
rect 29638 572296 29644 572308
rect 29696 572296 29702 572348
rect 19058 572228 19064 572280
rect 19116 572268 19122 572280
rect 57974 572268 57980 572280
rect 19116 572240 57980 572268
rect 19116 572228 19122 572240
rect 57974 572228 57980 572240
rect 58032 572228 58038 572280
rect 20530 572160 20536 572212
rect 20588 572200 20594 572212
rect 67634 572200 67640 572212
rect 20588 572172 67640 572200
rect 20588 572160 20594 572172
rect 67634 572160 67640 572172
rect 67692 572160 67698 572212
rect 525794 572160 525800 572212
rect 525852 572200 525858 572212
rect 570230 572200 570236 572212
rect 525852 572172 570236 572200
rect 525852 572160 525858 572172
rect 570230 572160 570236 572172
rect 570288 572160 570294 572212
rect 20622 572092 20628 572144
rect 20680 572132 20686 572144
rect 73154 572132 73160 572144
rect 20680 572104 73160 572132
rect 20680 572092 20686 572104
rect 73154 572092 73160 572104
rect 73212 572092 73218 572144
rect 270494 572092 270500 572144
rect 270552 572132 270558 572144
rect 294598 572132 294604 572144
rect 270552 572104 294604 572132
rect 270552 572092 270558 572104
rect 294598 572092 294604 572104
rect 294656 572092 294662 572144
rect 495434 572092 495440 572144
rect 495492 572132 495498 572144
rect 571518 572132 571524 572144
rect 495492 572104 571524 572132
rect 495492 572092 495498 572104
rect 571518 572092 571524 572104
rect 571576 572092 571582 572144
rect 19242 572024 19248 572076
rect 19300 572064 19306 572076
rect 78674 572064 78680 572076
rect 19300 572036 78680 572064
rect 19300 572024 19306 572036
rect 78674 572024 78680 572036
rect 78732 572024 78738 572076
rect 245654 572024 245660 572076
rect 245712 572064 245718 572076
rect 290090 572064 290096 572076
rect 245712 572036 290096 572064
rect 245712 572024 245718 572036
rect 290090 572024 290096 572036
rect 290148 572024 290154 572076
rect 469214 572024 469220 572076
rect 469272 572064 469278 572076
rect 572806 572064 572812 572076
rect 469272 572036 572812 572064
rect 469272 572024 469278 572036
rect 572806 572024 572812 572036
rect 572864 572024 572870 572076
rect 20438 571956 20444 572008
rect 20496 571996 20502 572008
rect 88334 571996 88340 572008
rect 20496 571968 88340 571996
rect 20496 571956 20502 571968
rect 88334 571956 88340 571968
rect 88392 571956 88398 572008
rect 158714 571956 158720 572008
rect 158772 571996 158778 572008
rect 288710 571996 288716 572008
rect 158772 571968 288716 571996
rect 158772 571956 158778 571968
rect 288710 571956 288716 571968
rect 288768 571956 288774 572008
rect 444374 571956 444380 572008
rect 444432 571996 444438 572008
rect 575474 571996 575480 572008
rect 444432 571968 575480 571996
rect 444432 571956 444438 571968
rect 575474 571956 575480 571968
rect 575532 571956 575538 572008
rect 577682 524424 577688 524476
rect 577740 524464 577746 524476
rect 579614 524464 579620 524476
rect 577740 524436 579620 524464
rect 577740 524424 577746 524436
rect 579614 524424 579620 524436
rect 579672 524424 579678 524476
rect 2866 514768 2872 514820
rect 2924 514808 2930 514820
rect 4798 514808 4804 514820
rect 2924 514780 4804 514808
rect 2924 514768 2930 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 2774 500964 2780 501016
rect 2832 501004 2838 501016
rect 7558 501004 7564 501016
rect 2832 500976 7564 501004
rect 2832 500964 2838 500976
rect 7558 500964 7564 500976
rect 7616 500964 7622 501016
rect 577498 484576 577504 484628
rect 577556 484616 577562 484628
rect 580626 484616 580632 484628
rect 577556 484588 580632 484616
rect 577556 484576 577562 484588
rect 580626 484576 580632 484588
rect 580684 484576 580690 484628
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 13078 462380 13084 462392
rect 3384 462352 13084 462380
rect 3384 462340 3390 462352
rect 13078 462340 13084 462352
rect 13136 462340 13142 462392
rect 285582 461592 285588 461644
rect 285640 461632 285646 461644
rect 292666 461632 292672 461644
rect 285640 461604 292672 461632
rect 285640 461592 285646 461604
rect 292666 461592 292672 461604
rect 292724 461592 292730 461644
rect 296530 461592 296536 461644
rect 296588 461632 296594 461644
rect 299382 461632 299388 461644
rect 296588 461604 299388 461632
rect 296588 461592 296594 461604
rect 299382 461592 299388 461604
rect 299440 461632 299446 461644
rect 399294 461632 399300 461644
rect 299440 461604 399300 461632
rect 299440 461592 299446 461604
rect 399294 461592 399300 461604
rect 399352 461592 399358 461644
rect 24946 461116 24952 461168
rect 25004 461156 25010 461168
rect 99006 461156 99012 461168
rect 25004 461128 99012 461156
rect 25004 461116 25010 461128
rect 99006 461116 99012 461128
rect 99064 461116 99070 461168
rect 22094 461048 22100 461100
rect 22152 461088 22158 461100
rect 23382 461088 23388 461100
rect 22152 461060 23388 461088
rect 22152 461048 22158 461060
rect 23382 461048 23388 461060
rect 23440 461048 23446 461100
rect 104388 461088 104394 461100
rect 23492 461060 104394 461088
rect 16390 460980 16396 461032
rect 16448 461020 16454 461032
rect 17586 461020 17592 461032
rect 16448 460992 17592 461020
rect 16448 460980 16454 460992
rect 17586 460980 17592 460992
rect 17644 461020 17650 461032
rect 23492 461020 23520 461060
rect 104388 461048 104394 461060
rect 104446 461048 104452 461100
rect 109448 461020 109454 461032
rect 17644 460992 23520 461020
rect 23584 460992 109454 461020
rect 17644 460980 17650 460992
rect 20346 460912 20352 460964
rect 20404 460952 20410 460964
rect 23584 460952 23612 460992
rect 109448 460980 109454 460992
rect 109506 460980 109512 461032
rect 391934 461020 391940 461032
rect 296686 460992 391940 461020
rect 296686 460964 296714 460992
rect 391934 460980 391940 460992
rect 391992 460980 391998 461032
rect 20404 460924 23612 460952
rect 20404 460912 20410 460924
rect 24854 460912 24860 460964
rect 24912 460952 24918 460964
rect 139486 460952 139492 460964
rect 24912 460924 139492 460952
rect 24912 460912 24918 460924
rect 139486 460912 139492 460924
rect 139544 460912 139550 460964
rect 296686 460952 296720 460964
rect 296548 460924 296720 460952
rect 17770 460844 17776 460896
rect 17828 460884 17834 460896
rect 24946 460884 24952 460896
rect 17828 460856 24952 460884
rect 17828 460844 17834 460856
rect 24946 460844 24952 460856
rect 25004 460844 25010 460896
rect 119246 460884 119252 460896
rect 26206 460856 119252 460884
rect 15010 460776 15016 460828
rect 15068 460816 15074 460828
rect 24854 460816 24860 460828
rect 15068 460788 24860 460816
rect 15068 460776 15074 460788
rect 24854 460776 24860 460788
rect 24912 460776 24918 460828
rect 17678 460708 17684 460760
rect 17736 460748 17742 460760
rect 26206 460748 26234 460856
rect 119246 460844 119252 460856
rect 119304 460844 119310 460896
rect 241330 460844 241336 460896
rect 241388 460884 241394 460896
rect 287606 460884 287612 460896
rect 241388 460856 287612 460884
rect 241388 460844 241394 460856
rect 287606 460844 287612 460856
rect 287664 460844 287670 460896
rect 295150 460844 295156 460896
rect 295208 460884 295214 460896
rect 296548 460884 296576 460924
rect 296714 460912 296720 460924
rect 296772 460912 296778 460964
rect 305086 460912 305092 460964
rect 305144 460952 305150 460964
rect 404630 460952 404636 460964
rect 305144 460924 404636 460952
rect 305144 460912 305150 460924
rect 404630 460912 404636 460924
rect 404688 460912 404694 460964
rect 575474 460952 575480 460964
rect 447060 460924 575480 460952
rect 295208 460856 296576 460884
rect 295208 460844 295214 460856
rect 296622 460844 296628 460896
rect 296680 460884 296686 460896
rect 297818 460884 297824 460896
rect 296680 460856 297824 460884
rect 296680 460844 296686 460856
rect 297818 460844 297824 460856
rect 297876 460884 297882 460896
rect 384390 460884 384396 460896
rect 297876 460856 384396 460884
rect 297876 460844 297882 460856
rect 384390 460844 384396 460856
rect 384448 460844 384454 460896
rect 391934 460844 391940 460896
rect 391992 460884 391998 460896
rect 394510 460884 394516 460896
rect 391992 460856 394516 460884
rect 391992 460844 391998 460856
rect 394510 460844 394516 460856
rect 394568 460844 394574 460896
rect 445110 460844 445116 460896
rect 445168 460884 445174 460896
rect 447060 460884 447088 460924
rect 575474 460912 575480 460924
rect 575532 460912 575538 460964
rect 445168 460856 447088 460884
rect 445168 460844 445174 460856
rect 470410 460844 470416 460896
rect 470468 460884 470474 460896
rect 572806 460884 572812 460896
rect 470468 460856 572812 460884
rect 470468 460844 470474 460856
rect 572806 460844 572812 460856
rect 572864 460844 572870 460896
rect 246390 460776 246396 460828
rect 246448 460816 246454 460828
rect 290182 460816 290188 460828
rect 246448 460788 290188 460816
rect 246448 460776 246454 460788
rect 290182 460776 290188 460788
rect 290240 460776 290246 460828
rect 300578 460776 300584 460828
rect 300636 460816 300642 460828
rect 359090 460816 359096 460828
rect 300636 460788 359096 460816
rect 300636 460776 300642 460788
rect 359090 460776 359096 460788
rect 359148 460776 359154 460828
rect 495710 460776 495716 460828
rect 495768 460816 495774 460828
rect 571518 460816 571524 460828
rect 495768 460788 571524 460816
rect 495768 460776 495774 460788
rect 571518 460776 571524 460788
rect 571576 460776 571582 460828
rect 17736 460720 26234 460748
rect 17736 460708 17742 460720
rect 256510 460708 256516 460760
rect 256568 460748 256574 460760
rect 286318 460748 286324 460760
rect 256568 460720 286324 460748
rect 256568 460708 256574 460720
rect 286318 460708 286324 460720
rect 286376 460748 286382 460760
rect 288526 460748 288532 460760
rect 286376 460720 288532 460748
rect 286376 460708 286382 460720
rect 288526 460708 288532 460720
rect 288584 460708 288590 460760
rect 521010 460708 521016 460760
rect 521068 460748 521074 460760
rect 567654 460748 567660 460760
rect 521068 460720 567660 460748
rect 521068 460708 521074 460720
rect 567654 460708 567660 460720
rect 567712 460708 567718 460760
rect 526070 460640 526076 460692
rect 526128 460680 526134 460692
rect 570230 460680 570236 460692
rect 526128 460652 570236 460680
rect 526128 460640 526134 460652
rect 570230 460640 570236 460652
rect 570288 460640 570294 460692
rect 536190 460572 536196 460624
rect 536248 460612 536254 460624
rect 568574 460612 568580 460624
rect 536248 460584 568580 460612
rect 536248 460572 536254 460584
rect 568574 460572 568580 460584
rect 568632 460572 568638 460624
rect 285490 460232 285496 460284
rect 285548 460272 285554 460284
rect 295518 460272 295524 460284
rect 285548 460244 295524 460272
rect 285548 460232 285554 460244
rect 295518 460232 295524 460244
rect 295576 460232 295582 460284
rect 14918 460164 14924 460216
rect 14976 460204 14982 460216
rect 129366 460204 129372 460216
rect 14976 460176 129372 460204
rect 14976 460164 14982 460176
rect 129366 460164 129372 460176
rect 129424 460164 129430 460216
rect 190454 460164 190460 460216
rect 190512 460204 190518 460216
rect 291838 460204 291844 460216
rect 190512 460176 291844 460204
rect 190512 460164 190518 460176
rect 291838 460164 291844 460176
rect 291896 460164 291902 460216
rect 343910 460204 343916 460216
rect 306346 460176 343916 460204
rect 287698 460028 287704 460080
rect 287756 460068 287762 460080
rect 288618 460068 288624 460080
rect 287756 460040 288624 460068
rect 287756 460028 287762 460040
rect 288618 460028 288624 460040
rect 288676 460028 288682 460080
rect 300394 460028 300400 460080
rect 300452 460068 300458 460080
rect 301774 460068 301780 460080
rect 300452 460040 301780 460068
rect 300452 460028 300458 460040
rect 301774 460028 301780 460040
rect 301832 460068 301838 460080
rect 306346 460068 306374 460176
rect 343910 460164 343916 460176
rect 343968 460164 343974 460216
rect 301832 460040 306374 460068
rect 301832 460028 301838 460040
rect 13722 459892 13728 459944
rect 13780 459932 13786 459944
rect 14918 459932 14924 459944
rect 13780 459904 14924 459932
rect 13780 459892 13786 459904
rect 14918 459892 14924 459904
rect 14976 459892 14982 459944
rect 301866 459892 301872 459944
rect 301924 459932 301930 459944
rect 303062 459932 303068 459944
rect 301924 459904 303068 459932
rect 301924 459892 301930 459904
rect 303062 459892 303068 459904
rect 303120 459892 303126 459944
rect 570046 459756 570052 459808
rect 570104 459796 570110 459808
rect 570230 459796 570236 459808
rect 570104 459768 570236 459796
rect 570104 459756 570110 459768
rect 570230 459756 570236 459768
rect 570288 459756 570294 459808
rect 572806 459620 572812 459672
rect 572864 459660 572870 459672
rect 574094 459660 574100 459672
rect 572864 459632 574100 459660
rect 572864 459620 572870 459632
rect 574094 459620 574100 459632
rect 574152 459620 574158 459672
rect 291838 459552 291844 459604
rect 291896 459592 291902 459604
rect 293954 459592 293960 459604
rect 291896 459564 293960 459592
rect 291896 459552 291902 459564
rect 293954 459552 293960 459564
rect 294012 459552 294018 459604
rect 298922 459552 298928 459604
rect 298980 459592 298986 459604
rect 300578 459592 300584 459604
rect 298980 459564 300584 459592
rect 298980 459552 298986 459564
rect 300578 459552 300584 459564
rect 300636 459552 300642 459604
rect 434990 459552 434996 459604
rect 435048 459592 435054 459604
rect 438118 459592 438124 459604
rect 435048 459564 438124 459592
rect 435048 459552 435054 459564
rect 438118 459552 438124 459564
rect 438176 459552 438182 459604
rect 571518 459552 571524 459604
rect 571576 459592 571582 459604
rect 572990 459592 572996 459604
rect 571576 459564 572996 459592
rect 571576 459552 571582 459564
rect 572990 459552 572996 459564
rect 573048 459552 573054 459604
rect 22002 459484 22008 459536
rect 22060 459524 22066 459536
rect 28166 459524 28172 459536
rect 22060 459496 28172 459524
rect 22060 459484 22066 459496
rect 28166 459484 28172 459496
rect 28224 459484 28230 459536
rect 144822 459484 144828 459536
rect 144880 459524 144886 459536
rect 149974 459524 149980 459536
rect 144880 459496 149980 459524
rect 144880 459484 144886 459496
rect 149974 459484 149980 459496
rect 150032 459484 150038 459536
rect 195790 459484 195796 459536
rect 195848 459524 195854 459536
rect 295334 459524 295340 459536
rect 195848 459496 295340 459524
rect 195848 459484 195854 459496
rect 295334 459484 295340 459496
rect 295392 459484 295398 459536
rect 302050 459484 302056 459536
rect 302108 459524 302114 459536
rect 313550 459524 313556 459536
rect 302108 459496 313556 459524
rect 302108 459484 302114 459496
rect 313550 459484 313556 459496
rect 313608 459484 313614 459536
rect 424870 459484 424876 459536
rect 424928 459524 424934 459536
rect 429930 459524 429936 459536
rect 424928 459496 429936 459524
rect 424928 459484 424934 459496
rect 429930 459484 429936 459496
rect 429988 459484 429994 459536
rect 546310 459484 546316 459536
rect 546368 459524 546374 459536
rect 556154 459524 556160 459536
rect 546368 459496 556160 459524
rect 546368 459484 546374 459496
rect 556154 459484 556160 459496
rect 556212 459484 556218 459536
rect 20622 459416 20628 459468
rect 20680 459456 20686 459468
rect 73706 459456 73712 459468
rect 20680 459428 73712 459456
rect 20680 459416 20686 459428
rect 73706 459416 73712 459428
rect 73764 459416 73770 459468
rect 185670 459416 185676 459468
rect 185728 459456 185734 459468
rect 285398 459456 285404 459468
rect 185728 459428 285404 459456
rect 185728 459416 185734 459428
rect 285398 459416 285404 459428
rect 285456 459456 285462 459468
rect 287790 459456 287796 459468
rect 285456 459428 287796 459456
rect 285456 459416 285462 459428
rect 287790 459416 287796 459428
rect 287848 459416 287854 459468
rect 301866 459416 301872 459468
rect 301924 459456 301930 459468
rect 389450 459456 389456 459468
rect 301924 459428 389456 459456
rect 301924 459416 301930 459428
rect 389450 459416 389456 459428
rect 389508 459416 389514 459468
rect 450170 459416 450176 459468
rect 450228 459456 450234 459468
rect 564434 459456 564440 459468
rect 450228 459428 564440 459456
rect 450228 459416 450234 459428
rect 564434 459416 564440 459428
rect 564492 459416 564498 459468
rect 19058 459348 19064 459400
rect 19116 459388 19122 459400
rect 58526 459388 58532 459400
rect 19116 459360 58532 459388
rect 19116 459348 19122 459360
rect 58526 459348 58532 459360
rect 58584 459348 58590 459400
rect 266262 459348 266268 459400
rect 266320 459388 266326 459400
rect 289998 459388 290004 459400
rect 266320 459360 290004 459388
rect 266320 459348 266326 459360
rect 289998 459348 290004 459360
rect 290056 459348 290062 459400
rect 299198 459348 299204 459400
rect 299256 459388 299262 459400
rect 374270 459388 374276 459400
rect 299256 459360 374276 459388
rect 299256 459348 299262 459360
rect 374270 459348 374276 459360
rect 374328 459348 374334 459400
rect 460290 459348 460296 459400
rect 460348 459388 460354 459400
rect 572714 459388 572720 459400
rect 460348 459360 572720 459388
rect 460348 459348 460354 459360
rect 572714 459348 572720 459360
rect 572772 459348 572778 459400
rect 20438 459280 20444 459332
rect 20496 459320 20502 459332
rect 88886 459320 88892 459332
rect 20496 459292 88892 459320
rect 20496 459280 20502 459292
rect 88886 459280 88892 459292
rect 88944 459280 88950 459332
rect 299290 459280 299296 459332
rect 299348 459320 299354 459332
rect 354030 459320 354036 459332
rect 299348 459292 354036 459320
rect 299348 459280 299354 459292
rect 354030 459280 354036 459292
rect 354088 459280 354094 459332
rect 465350 459280 465356 459332
rect 465408 459320 465414 459332
rect 567746 459320 567752 459332
rect 465408 459292 567752 459320
rect 465408 459280 465414 459292
rect 567746 459280 567752 459292
rect 567804 459280 567810 459332
rect 303062 459212 303068 459264
rect 303120 459252 303126 459264
rect 318610 459252 318616 459264
rect 303120 459224 318616 459252
rect 303120 459212 303126 459224
rect 318610 459212 318616 459224
rect 318668 459212 318674 459264
rect 531130 459212 531136 459264
rect 531188 459252 531194 459264
rect 569954 459252 569960 459264
rect 531188 459224 569960 459252
rect 531188 459212 531194 459224
rect 569954 459212 569960 459224
rect 570012 459212 570018 459264
rect 313274 459144 313280 459196
rect 313332 459184 313338 459196
rect 323670 459184 323676 459196
rect 313332 459156 323676 459184
rect 313332 459144 313338 459156
rect 323670 459144 323676 459156
rect 323728 459144 323734 459196
rect 308490 459076 308496 459128
rect 308548 459116 308554 459128
rect 580258 459116 580264 459128
rect 308548 459088 580264 459116
rect 308548 459076 308554 459088
rect 580258 459076 580264 459088
rect 580316 459076 580322 459128
rect 20530 458940 20536 458992
rect 20588 458980 20594 458992
rect 21634 458980 21640 458992
rect 20588 458952 21640 458980
rect 20588 458940 20594 458952
rect 21634 458940 21640 458952
rect 21692 458980 21698 458992
rect 21692 458952 26234 458980
rect 21692 458940 21698 458952
rect 26206 458912 26234 458952
rect 34514 458940 34520 458992
rect 34572 458980 34578 458992
rect 38286 458980 38292 458992
rect 34572 458952 38292 458980
rect 34572 458940 34578 458952
rect 38286 458940 38292 458952
rect 38344 458940 38350 458992
rect 216030 458940 216036 458992
rect 216088 458980 216094 458992
rect 288526 458980 288532 458992
rect 216088 458952 288532 458980
rect 216088 458940 216094 458952
rect 288526 458940 288532 458952
rect 288584 458980 288590 458992
rect 291194 458980 291200 458992
rect 288584 458952 291200 458980
rect 288584 458940 288590 458952
rect 291194 458940 291200 458952
rect 291252 458940 291258 458992
rect 68646 458912 68652 458924
rect 26206 458884 68652 458912
rect 68646 458872 68652 458884
rect 68704 458872 68710 458924
rect 180610 458872 180616 458924
rect 180668 458912 180674 458924
rect 292758 458912 292764 458924
rect 180668 458884 292764 458912
rect 180668 458872 180674 458884
rect 292758 458872 292764 458884
rect 292816 458912 292822 458924
rect 295426 458912 295432 458924
rect 292816 458884 295432 458912
rect 292816 458872 292822 458884
rect 295426 458872 295432 458884
rect 295484 458872 295490 458924
rect 17862 458804 17868 458856
rect 17920 458844 17926 458856
rect 18782 458844 18788 458856
rect 17920 458816 18788 458844
rect 17920 458804 17926 458816
rect 18782 458804 18788 458816
rect 18840 458804 18846 458856
rect 19242 458804 19248 458856
rect 19300 458844 19306 458856
rect 20346 458844 20352 458856
rect 19300 458816 20352 458844
rect 19300 458804 19306 458816
rect 20346 458804 20352 458816
rect 20404 458844 20410 458856
rect 78766 458844 78772 458856
rect 20404 458816 78772 458844
rect 20404 458804 20410 458816
rect 78766 458804 78772 458816
rect 78824 458804 78830 458856
rect 149974 458804 149980 458856
rect 150032 458844 150038 458856
rect 288434 458844 288440 458856
rect 150032 458816 288440 458844
rect 150032 458804 150038 458816
rect 288434 458804 288440 458816
rect 288492 458804 288498 458856
rect 556430 458804 556436 458856
rect 556488 458844 556494 458856
rect 571426 458844 571432 458856
rect 556488 458816 571432 458844
rect 556488 458804 556494 458816
rect 571426 458804 571432 458816
rect 571484 458804 571490 458856
rect 27798 458464 27804 458516
rect 27856 458504 27862 458516
rect 33226 458504 33232 458516
rect 27856 458476 33232 458504
rect 27856 458464 27862 458476
rect 33226 458464 33232 458476
rect 33284 458464 33290 458516
rect 110414 458192 110420 458244
rect 110472 458232 110478 458244
rect 114186 458232 114192 458244
rect 110472 458204 114192 458232
rect 110472 458192 110478 458204
rect 114186 458192 114192 458204
rect 114244 458192 114250 458244
rect 289998 458192 290004 458244
rect 290056 458232 290062 458244
rect 290274 458232 290280 458244
rect 290056 458204 290280 458232
rect 290056 458192 290062 458204
rect 290274 458192 290280 458204
rect 290332 458192 290338 458244
rect 369210 458232 369216 458244
rect 367112 458204 369216 458232
rect 23290 458124 23296 458176
rect 23348 458164 23354 458176
rect 30926 458164 30932 458176
rect 23348 458136 30932 458164
rect 23348 458124 23354 458136
rect 30926 458124 30932 458136
rect 30984 458124 30990 458176
rect 63586 458164 63592 458176
rect 31036 458136 63592 458164
rect 21910 458056 21916 458108
rect 21968 458096 21974 458108
rect 23106 458096 23112 458108
rect 21968 458068 23112 458096
rect 21968 458056 21974 458068
rect 23106 458056 23112 458068
rect 23164 458096 23170 458108
rect 27798 458096 27804 458108
rect 23164 458068 27804 458096
rect 23164 458056 23170 458068
rect 27798 458056 27804 458068
rect 27856 458056 27862 458108
rect 31036 458096 31064 458136
rect 63586 458124 63592 458136
rect 63644 458124 63650 458176
rect 226150 458124 226156 458176
rect 226208 458164 226214 458176
rect 287514 458164 287520 458176
rect 226208 458136 287520 458164
rect 226208 458124 226214 458136
rect 287514 458124 287520 458136
rect 287572 458124 287578 458176
rect 298002 458124 298008 458176
rect 298060 458164 298066 458176
rect 367112 458164 367140 458204
rect 369210 458192 369216 458204
rect 369268 458192 369274 458244
rect 424318 458192 424324 458244
rect 424376 458232 424382 458244
rect 424870 458232 424876 458244
rect 424376 458204 424876 458232
rect 424376 458192 424382 458204
rect 424870 458192 424876 458204
rect 424928 458192 424934 458244
rect 500770 458192 500776 458244
rect 500828 458232 500834 458244
rect 500828 458204 502380 458232
rect 500828 458192 500834 458204
rect 298060 458136 367140 458164
rect 502352 458164 502380 458204
rect 569954 458192 569960 458244
rect 570012 458232 570018 458244
rect 571518 458232 571524 458244
rect 570012 458204 571524 458232
rect 570012 458192 570018 458204
rect 571518 458192 571524 458204
rect 571576 458192 571582 458244
rect 572714 458192 572720 458244
rect 572772 458232 572778 458244
rect 575474 458232 575480 458244
rect 572772 458204 575480 458232
rect 572772 458192 572778 458204
rect 575474 458192 575480 458204
rect 575532 458192 575538 458244
rect 568942 458164 568948 458176
rect 502352 458136 568948 458164
rect 298060 458124 298066 458136
rect 568942 458124 568948 458136
rect 569000 458164 569006 458176
rect 570598 458164 570604 458176
rect 569000 458136 570604 458164
rect 569000 458124 569006 458136
rect 570598 458124 570604 458136
rect 570656 458124 570662 458176
rect 53466 458096 53472 458108
rect 30852 458068 31064 458096
rect 31220 458068 53472 458096
rect 23198 457920 23204 457972
rect 23256 457960 23262 457972
rect 30852 457960 30880 458068
rect 23256 457932 30880 457960
rect 23256 457920 23262 457932
rect 21726 457852 21732 457904
rect 21784 457892 21790 457904
rect 31220 457892 31248 458068
rect 53466 458056 53472 458068
rect 53524 458056 53530 458108
rect 231210 458056 231216 458108
rect 231268 458096 231274 458108
rect 288802 458096 288808 458108
rect 231268 458068 288808 458096
rect 231268 458056 231274 458068
rect 288802 458056 288808 458068
rect 288860 458096 288866 458108
rect 291286 458096 291292 458108
rect 288860 458068 291292 458096
rect 288860 458056 288866 458068
rect 291286 458056 291292 458068
rect 291344 458056 291350 458108
rect 300670 458056 300676 458108
rect 300728 458096 300734 458108
rect 338850 458096 338856 458108
rect 300728 458068 338856 458096
rect 300728 458056 300734 458068
rect 338850 458056 338856 458068
rect 338908 458056 338914 458108
rect 505830 458056 505836 458108
rect 505888 458096 505894 458108
rect 565906 458096 565912 458108
rect 505888 458068 565912 458096
rect 505888 458056 505894 458068
rect 565906 458056 565912 458068
rect 565964 458056 565970 458108
rect 48498 458028 48504 458040
rect 21784 457864 31248 457892
rect 35866 458000 48504 458028
rect 21784 457852 21790 457864
rect 30926 457784 30932 457836
rect 30984 457824 30990 457836
rect 35866 457824 35894 458000
rect 48498 457988 48504 458000
rect 48556 457988 48562 458040
rect 251082 457988 251088 458040
rect 251140 458028 251146 458040
rect 289814 458028 289820 458040
rect 251140 458000 289820 458028
rect 251140 457988 251146 458000
rect 289814 457988 289820 458000
rect 289872 457988 289878 458040
rect 303246 457988 303252 458040
rect 303304 458028 303310 458040
rect 333790 458028 333796 458040
rect 303304 458000 333796 458028
rect 303304 457988 303310 458000
rect 333790 457988 333796 458000
rect 333848 457988 333854 458040
rect 510890 457988 510896 458040
rect 510948 458028 510954 458040
rect 570138 458028 570144 458040
rect 510948 458000 570144 458028
rect 510948 457988 510954 458000
rect 570138 457988 570144 458000
rect 570196 457988 570202 458040
rect 302142 457920 302148 457972
rect 302200 457960 302206 457972
rect 328730 457960 328736 457972
rect 302200 457932 328736 457960
rect 302200 457920 302206 457932
rect 328730 457920 328736 457932
rect 328788 457920 328794 457972
rect 515950 457920 515956 457972
rect 516008 457960 516014 457972
rect 570322 457960 570328 457972
rect 516008 457932 570328 457960
rect 516008 457920 516014 457932
rect 570322 457920 570328 457932
rect 570380 457920 570386 457972
rect 541250 457852 541256 457904
rect 541308 457892 541314 457904
rect 567562 457892 567568 457904
rect 541308 457864 567568 457892
rect 541308 457852 541314 457864
rect 567562 457852 567568 457864
rect 567620 457852 567626 457904
rect 30984 457796 35894 457824
rect 30984 457784 30990 457796
rect 300394 457580 300400 457632
rect 300452 457620 300458 457632
rect 303246 457620 303252 457632
rect 300452 457592 303252 457620
rect 300452 457580 300458 457592
rect 303246 457580 303252 457592
rect 303304 457580 303310 457632
rect 261570 457512 261576 457564
rect 261628 457552 261634 457564
rect 289078 457552 289084 457564
rect 261628 457524 289084 457552
rect 261628 457512 261634 457524
rect 289078 457512 289084 457524
rect 289136 457552 289142 457564
rect 289906 457552 289912 457564
rect 289136 457524 289912 457552
rect 289136 457512 289142 457524
rect 289906 457512 289912 457524
rect 289964 457512 289970 457564
rect 21818 457444 21824 457496
rect 21876 457484 21882 457496
rect 23014 457484 23020 457496
rect 21876 457456 23020 457484
rect 21876 457444 21882 457456
rect 23014 457444 23020 457456
rect 23072 457484 23078 457496
rect 43346 457484 43352 457496
rect 23072 457456 43352 457484
rect 23072 457444 23078 457456
rect 43346 457444 43352 457456
rect 43404 457444 43410 457496
rect 235902 457444 235908 457496
rect 235960 457484 235966 457496
rect 291194 457484 291200 457496
rect 235960 457456 291200 457484
rect 235960 457444 235966 457456
rect 291194 457444 291200 457456
rect 291252 457484 291258 457496
rect 292574 457484 292580 457496
rect 291252 457456 292580 457484
rect 291252 457444 291258 457456
rect 292574 457444 292580 457456
rect 292632 457444 292638 457496
rect 301958 457444 301964 457496
rect 302016 457484 302022 457496
rect 303246 457484 303252 457496
rect 302016 457456 303252 457484
rect 302016 457444 302022 457456
rect 303246 457444 303252 457456
rect 303304 457484 303310 457496
rect 364150 457484 364156 457496
rect 303304 457456 364156 457484
rect 303304 457444 303310 457456
rect 364150 457444 364156 457456
rect 364208 457444 364214 457496
rect 21726 456832 21732 456884
rect 21784 456872 21790 456884
rect 23198 456872 23204 456884
rect 21784 456844 23204 456872
rect 21784 456832 21790 456844
rect 23198 456832 23204 456844
rect 23256 456832 23262 456884
rect 22738 456764 22744 456816
rect 22796 456804 22802 456816
rect 23290 456804 23296 456816
rect 22796 456776 23296 456804
rect 22796 456764 22802 456776
rect 23290 456764 23296 456776
rect 23348 456764 23354 456816
rect 570322 456764 570328 456816
rect 570380 456804 570386 456816
rect 572806 456804 572812 456816
rect 570380 456776 572812 456804
rect 570380 456764 570386 456776
rect 572806 456764 572812 456776
rect 572864 456764 572870 456816
rect 299106 456696 299112 456748
rect 299164 456736 299170 456748
rect 409690 456736 409696 456748
rect 299164 456708 409696 456736
rect 299164 456696 299170 456708
rect 409690 456696 409696 456708
rect 409748 456696 409754 456748
rect 301866 456628 301872 456680
rect 301924 456668 301930 456680
rect 302970 456668 302976 456680
rect 301924 456640 302976 456668
rect 301924 456628 301930 456640
rect 302970 456628 302976 456640
rect 303028 456668 303034 456680
rect 379330 456668 379336 456680
rect 303028 456640 379336 456668
rect 303028 456628 303034 456640
rect 379330 456628 379336 456640
rect 379388 456628 379394 456680
rect 304994 456016 305000 456068
rect 305052 456056 305058 456068
rect 419810 456056 419816 456068
rect 305052 456028 419816 456056
rect 305052 456016 305058 456028
rect 419810 456016 419816 456028
rect 419868 456016 419874 456068
rect 15102 455336 15108 455388
rect 15160 455376 15166 455388
rect 17862 455376 17868 455388
rect 15160 455348 17868 455376
rect 15160 455336 15166 455348
rect 17862 455336 17868 455348
rect 17920 455336 17926 455388
rect 19150 455336 19156 455388
rect 19208 455376 19214 455388
rect 154758 455376 154764 455388
rect 19208 455348 154764 455376
rect 19208 455336 19214 455348
rect 154758 455336 154764 455348
rect 154816 455336 154822 455388
rect 295242 455336 295248 455388
rect 295300 455376 295306 455388
rect 304994 455376 305000 455388
rect 295300 455348 305000 455376
rect 295300 455336 295306 455348
rect 304994 455336 305000 455348
rect 305052 455336 305058 455388
rect 440050 455336 440056 455388
rect 440108 455376 440114 455388
rect 564894 455376 564900 455388
rect 440108 455348 564900 455376
rect 440108 455336 440114 455348
rect 564894 455336 564900 455348
rect 564952 455336 564958 455388
rect 17218 454656 17224 454708
rect 17276 454696 17282 454708
rect 17862 454696 17868 454708
rect 17276 454668 17868 454696
rect 17276 454656 17282 454668
rect 17862 454656 17868 454668
rect 17920 454696 17926 454708
rect 110414 454696 110420 454708
rect 17920 454668 110420 454696
rect 17920 454656 17926 454668
rect 110414 454656 110420 454668
rect 110472 454656 110478 454708
rect 564894 454656 564900 454708
rect 564952 454696 564958 454708
rect 571610 454696 571616 454708
rect 564952 454668 571616 454696
rect 564952 454656 564958 454668
rect 571610 454656 571616 454668
rect 571668 454656 571674 454708
rect 21358 444320 21364 444372
rect 21416 444360 21422 444372
rect 24854 444360 24860 444372
rect 21416 444332 24860 444360
rect 21416 444320 21422 444332
rect 24854 444320 24860 444332
rect 24912 444320 24918 444372
rect 219434 444320 219440 444372
rect 219492 444360 219498 444372
rect 291470 444360 291476 444372
rect 219492 444332 291476 444360
rect 219492 444320 219498 444332
rect 291470 444320 291476 444332
rect 291528 444320 291534 444372
rect 300762 444320 300768 444372
rect 300820 444360 300826 444372
rect 347774 444360 347780 444372
rect 300820 444332 347780 444360
rect 300820 444320 300826 444332
rect 347774 444320 347780 444332
rect 347832 444320 347838 444372
rect 438118 444320 438124 444372
rect 438176 444360 438182 444372
rect 565538 444360 565544 444372
rect 438176 444332 565544 444360
rect 438176 444320 438182 444332
rect 565538 444320 565544 444332
rect 565596 444320 565602 444372
rect 270494 444252 270500 444304
rect 270552 444292 270558 444304
rect 297174 444292 297180 444304
rect 270552 444264 297180 444292
rect 270552 444252 270558 444264
rect 297174 444252 297180 444264
rect 297232 444252 297238 444304
rect 474734 444252 474740 444304
rect 474792 444292 474798 444304
rect 574186 444292 574192 444304
rect 474792 444264 574192 444292
rect 474792 444252 474798 444264
rect 574186 444252 574192 444264
rect 574244 444252 574250 444304
rect 291470 443912 291476 443964
rect 291528 443952 291534 443964
rect 292850 443952 292856 443964
rect 291528 443924 292856 443952
rect 291528 443912 291534 443924
rect 292850 443912 292856 443924
rect 292908 443912 292914 443964
rect 23474 443640 23480 443692
rect 23532 443680 23538 443692
rect 200114 443680 200120 443692
rect 23532 443652 200120 443680
rect 23532 443640 23538 443652
rect 200114 443640 200120 443652
rect 200172 443640 200178 443692
rect 300302 443504 300308 443556
rect 300360 443544 300366 443556
rect 300762 443544 300768 443556
rect 300360 443516 300768 443544
rect 300360 443504 300366 443516
rect 300762 443504 300768 443516
rect 300820 443504 300826 443556
rect 565538 442960 565544 443012
rect 565596 443000 565602 443012
rect 568850 443000 568856 443012
rect 565596 442972 568856 443000
rect 565596 442960 565602 442972
rect 568850 442960 568856 442972
rect 568908 442960 568914 443012
rect 164234 442892 164240 442944
rect 164292 442932 164298 442944
rect 284294 442932 284300 442944
rect 164292 442904 284300 442932
rect 164292 442892 164298 442904
rect 284294 442892 284300 442904
rect 284352 442892 284358 442944
rect 169754 442824 169760 442876
rect 169812 442864 169818 442876
rect 284938 442864 284944 442876
rect 169812 442836 284944 442864
rect 169812 442824 169818 442836
rect 284938 442824 284944 442836
rect 284996 442864 285002 442876
rect 285582 442864 285588 442876
rect 284996 442836 285588 442864
rect 284996 442824 285002 442836
rect 285582 442824 285588 442836
rect 285640 442824 285646 442876
rect 13170 442212 13176 442264
rect 13228 442252 13234 442264
rect 23474 442252 23480 442264
rect 13228 442224 23480 442252
rect 13228 442212 13234 442224
rect 23474 442212 23480 442224
rect 23532 442212 23538 442264
rect 284294 442212 284300 442264
rect 284352 442252 284358 442264
rect 285490 442252 285496 442264
rect 284352 442224 285496 442252
rect 284352 442212 284358 442224
rect 285490 442212 285496 442224
rect 285548 442252 285554 442264
rect 296806 442252 296812 442264
rect 285548 442224 296812 442252
rect 285548 442212 285554 442224
rect 296806 442212 296812 442224
rect 296864 442212 296870 442264
rect 284938 441872 284944 441924
rect 284996 441912 285002 441924
rect 288618 441912 288624 441924
rect 284996 441884 288624 441912
rect 284996 441872 285002 441884
rect 288618 441872 288624 441884
rect 288676 441872 288682 441924
rect 3142 410048 3148 410100
rect 3200 410088 3206 410100
rect 6178 410088 6184 410100
rect 3200 410060 6184 410088
rect 3200 410048 3206 410060
rect 6178 410048 6184 410060
rect 6236 410048 6242 410100
rect 2774 398760 2780 398812
rect 2832 398800 2838 398812
rect 7650 398800 7656 398812
rect 2832 398772 7656 398800
rect 2832 398760 2838 398772
rect 7650 398760 7656 398772
rect 7708 398760 7714 398812
rect 577590 364692 577596 364744
rect 577648 364732 577654 364744
rect 580626 364732 580632 364744
rect 577648 364704 580632 364732
rect 577648 364692 577654 364704
rect 580626 364692 580632 364704
rect 580684 364692 580690 364744
rect 2958 357416 2964 357468
rect 3016 357456 3022 357468
rect 6270 357456 6276 357468
rect 3016 357428 6276 357456
rect 3016 357416 3022 357428
rect 6270 357416 6276 357428
rect 6328 357416 6334 357468
rect 3326 345312 3332 345364
rect 3384 345352 3390 345364
rect 8938 345352 8944 345364
rect 3384 345324 8944 345352
rect 3384 345312 3390 345324
rect 8938 345312 8944 345324
rect 8996 345312 9002 345364
rect 17402 333956 17408 334008
rect 17460 333996 17466 334008
rect 21358 333996 21364 334008
rect 17460 333968 21364 333996
rect 17460 333956 17466 333968
rect 21358 333956 21364 333968
rect 21416 333956 21422 334008
rect 570598 333956 570604 334008
rect 570656 333996 570662 334008
rect 574462 333996 574468 334008
rect 570656 333968 574468 333996
rect 570656 333956 570662 333968
rect 574462 333956 574468 333968
rect 574520 333956 574526 334008
rect 300486 333616 300492 333668
rect 300544 333656 300550 333668
rect 304994 333656 305000 333668
rect 300544 333628 305000 333656
rect 300544 333616 300550 333628
rect 304994 333616 305000 333628
rect 305052 333616 305058 333668
rect 285582 333276 285588 333328
rect 285640 333316 285646 333328
rect 292758 333316 292764 333328
rect 285640 333288 292764 333316
rect 285640 333276 285646 333288
rect 292758 333276 292764 333288
rect 292816 333276 292822 333328
rect 295242 333276 295248 333328
rect 295300 333316 295306 333328
rect 305086 333316 305092 333328
rect 295300 333288 305092 333316
rect 295300 333276 295306 333288
rect 305086 333276 305092 333288
rect 305144 333276 305150 333328
rect 501138 333276 501144 333328
rect 501196 333316 501202 333328
rect 570598 333316 570604 333328
rect 501196 333288 570604 333316
rect 501196 333276 501202 333288
rect 570598 333276 570604 333288
rect 570656 333276 570662 333328
rect 20438 333208 20444 333260
rect 20496 333248 20502 333260
rect 88886 333248 88892 333260
rect 20496 333220 88892 333248
rect 20496 333208 20502 333220
rect 88886 333208 88892 333220
rect 88944 333208 88950 333260
rect 284202 333208 284208 333260
rect 284260 333248 284266 333260
rect 296806 333248 296812 333260
rect 284260 333220 296812 333248
rect 284260 333208 284266 333220
rect 296806 333208 296812 333220
rect 296864 333208 296870 333260
rect 475746 333208 475752 333260
rect 475804 333248 475810 333260
rect 574186 333248 574192 333260
rect 475804 333220 574192 333248
rect 475804 333208 475810 333220
rect 574186 333208 574192 333220
rect 574244 333208 574250 333260
rect 18874 332936 18880 332988
rect 18932 332976 18938 332988
rect 20438 332976 20444 332988
rect 18932 332948 20444 332976
rect 18932 332936 18938 332948
rect 20438 332936 20444 332948
rect 20496 332936 20502 332988
rect 20346 332868 20352 332920
rect 20404 332908 20410 332920
rect 78766 332908 78772 332920
rect 20404 332880 78772 332908
rect 20404 332868 20410 332880
rect 78766 332868 78772 332880
rect 78824 332868 78830 332920
rect 20254 332800 20260 332852
rect 20312 332840 20318 332852
rect 109126 332840 109132 332852
rect 20312 332812 109132 332840
rect 20312 332800 20318 332812
rect 109126 332800 109132 332812
rect 109184 332800 109190 332852
rect 20162 332732 20168 332784
rect 20220 332772 20226 332784
rect 20346 332772 20352 332784
rect 20220 332744 20352 332772
rect 20220 332732 20226 332744
rect 20346 332732 20352 332744
rect 20404 332732 20410 332784
rect 21358 332732 21364 332784
rect 21416 332772 21422 332784
rect 124306 332772 124312 332784
rect 21416 332744 124312 332772
rect 21416 332732 21422 332744
rect 124306 332732 124312 332744
rect 124364 332732 124370 332784
rect 299106 332732 299112 332784
rect 299164 332772 299170 332784
rect 303706 332772 303712 332784
rect 299164 332744 303712 332772
rect 299164 332732 299170 332744
rect 303706 332732 303712 332744
rect 303764 332732 303770 332784
rect 14918 332664 14924 332716
rect 14976 332704 14982 332716
rect 15102 332704 15108 332716
rect 14976 332676 15108 332704
rect 14976 332664 14982 332676
rect 15102 332664 15108 332676
rect 15160 332704 15166 332716
rect 129366 332704 129372 332716
rect 15160 332676 129372 332704
rect 15160 332664 15166 332676
rect 129366 332664 129372 332676
rect 129424 332664 129430 332716
rect 231210 332664 231216 332716
rect 231268 332704 231274 332716
rect 291286 332704 291292 332716
rect 231268 332676 291292 332704
rect 231268 332664 231274 332676
rect 291286 332664 291292 332676
rect 291344 332664 291350 332716
rect 296622 332664 296628 332716
rect 296680 332704 296686 332716
rect 384022 332704 384028 332716
rect 296680 332676 384028 332704
rect 296680 332664 296686 332676
rect 384022 332664 384028 332676
rect 384080 332664 384086 332716
rect 574186 332664 574192 332716
rect 574244 332704 574250 332716
rect 575750 332704 575756 332716
rect 574244 332676 575756 332704
rect 574244 332664 574250 332676
rect 575750 332664 575756 332676
rect 575808 332664 575814 332716
rect 15010 332596 15016 332648
rect 15068 332636 15074 332648
rect 139486 332636 139492 332648
rect 15068 332608 139492 332636
rect 15068 332596 15074 332608
rect 139486 332596 139492 332608
rect 139544 332596 139550 332648
rect 210970 332596 210976 332648
rect 211028 332636 211034 332648
rect 287606 332636 287612 332648
rect 211028 332608 287612 332636
rect 211028 332596 211034 332608
rect 287606 332596 287612 332608
rect 287664 332596 287670 332648
rect 305086 332596 305092 332648
rect 305144 332636 305150 332648
rect 419810 332636 419816 332648
rect 305144 332608 419816 332636
rect 305144 332596 305150 332608
rect 419810 332596 419816 332608
rect 419868 332596 419874 332648
rect 575658 332636 575664 332648
rect 447060 332608 575664 332636
rect 22738 332528 22744 332580
rect 22796 332568 22802 332580
rect 22796 332540 23612 332568
rect 22796 332528 22802 332540
rect 3602 332460 3608 332512
rect 3660 332500 3666 332512
rect 23106 332500 23112 332512
rect 3660 332472 23112 332500
rect 3660 332460 3666 332472
rect 23106 332460 23112 332472
rect 23164 332460 23170 332512
rect 23584 332500 23612 332540
rect 23658 332528 23664 332580
rect 23716 332568 23722 332580
rect 63586 332568 63592 332580
rect 23716 332540 63592 332568
rect 23716 332528 23722 332540
rect 63586 332528 63592 332540
rect 63644 332528 63650 332580
rect 144822 332528 144828 332580
rect 144880 332568 144886 332580
rect 149606 332568 149612 332580
rect 144880 332540 149612 332568
rect 144880 332528 144886 332540
rect 149606 332528 149612 332540
rect 149664 332528 149670 332580
rect 246390 332528 246396 332580
rect 246448 332568 246454 332580
rect 290182 332568 290188 332580
rect 246448 332540 290188 332568
rect 246448 332528 246454 332540
rect 290182 332528 290188 332540
rect 290240 332528 290246 332580
rect 301866 332528 301872 332580
rect 301924 332568 301930 332580
rect 306374 332568 306380 332580
rect 301924 332540 306380 332568
rect 301924 332528 301930 332540
rect 306374 332528 306380 332540
rect 306432 332528 306438 332580
rect 318610 332568 318616 332580
rect 311176 332540 318616 332568
rect 48406 332500 48412 332512
rect 23584 332472 48412 332500
rect 48406 332460 48412 332472
rect 48464 332460 48470 332512
rect 251082 332460 251088 332512
rect 251140 332500 251146 332512
rect 289814 332500 289820 332512
rect 251140 332472 289820 332500
rect 251140 332460 251146 332472
rect 289814 332460 289820 332472
rect 289872 332460 289878 332512
rect 303062 332460 303068 332512
rect 303120 332500 303126 332512
rect 311176 332500 311204 332540
rect 318610 332528 318616 332540
rect 318668 332528 318674 332580
rect 424318 332528 424324 332580
rect 424376 332568 424382 332580
rect 424870 332568 424876 332580
rect 424376 332540 424876 332568
rect 424376 332528 424382 332540
rect 424870 332528 424876 332540
rect 424928 332568 424934 332580
rect 429930 332568 429936 332580
rect 424928 332540 429936 332568
rect 424928 332528 424934 332540
rect 429930 332528 429936 332540
rect 429988 332528 429994 332580
rect 445110 332528 445116 332580
rect 445168 332568 445174 332580
rect 447060 332568 447088 332608
rect 575658 332596 575664 332608
rect 575716 332596 575722 332648
rect 445168 332540 447088 332568
rect 445168 332528 445174 332540
rect 303120 332472 311204 332500
rect 303120 332460 303126 332472
rect 311250 332460 311256 332512
rect 311308 332500 311314 332512
rect 333790 332500 333796 332512
rect 311308 332472 333796 332500
rect 311308 332460 311314 332472
rect 333790 332460 333796 332472
rect 333848 332460 333854 332512
rect 536190 332460 536196 332512
rect 536248 332500 536254 332512
rect 568574 332500 568580 332512
rect 536248 332472 568580 332500
rect 536248 332460 536254 332472
rect 568574 332460 568580 332472
rect 568632 332460 568638 332512
rect 22922 332392 22928 332444
rect 22980 332432 22986 332444
rect 43346 332432 43352 332444
rect 22980 332404 43352 332432
rect 22980 332392 22986 332404
rect 43346 332392 43352 332404
rect 43404 332392 43410 332444
rect 256510 332392 256516 332444
rect 256568 332432 256574 332444
rect 281350 332432 281356 332444
rect 256568 332404 281356 332432
rect 256568 332392 256574 332404
rect 281350 332392 281356 332404
rect 281408 332392 281414 332444
rect 281442 332392 281448 332444
rect 281500 332432 281506 332444
rect 287698 332432 287704 332444
rect 281500 332404 287704 332432
rect 281500 332392 281506 332404
rect 287698 332392 287704 332404
rect 287756 332392 287762 332444
rect 302142 332392 302148 332444
rect 302200 332432 302206 332444
rect 328730 332432 328736 332444
rect 302200 332404 328736 332432
rect 302200 332392 302206 332404
rect 328730 332392 328736 332404
rect 328788 332392 328794 332444
rect 541250 332392 541256 332444
rect 541308 332432 541314 332444
rect 567562 332432 567568 332444
rect 541308 332404 567568 332432
rect 541308 332392 541314 332404
rect 567562 332392 567568 332404
rect 567620 332392 567626 332444
rect 22830 332324 22836 332376
rect 22888 332364 22894 332376
rect 38286 332364 38292 332376
rect 22888 332336 38292 332364
rect 22888 332324 22894 332336
rect 38286 332324 38292 332336
rect 38344 332324 38350 332376
rect 261570 332324 261576 332376
rect 261628 332364 261634 332376
rect 282178 332364 282184 332376
rect 261628 332336 282184 332364
rect 261628 332324 261634 332336
rect 282178 332324 282184 332336
rect 282236 332324 282242 332376
rect 303154 332324 303160 332376
rect 303212 332364 303218 332376
rect 323670 332364 323676 332376
rect 303212 332336 323676 332364
rect 303212 332324 303218 332336
rect 323670 332324 323676 332336
rect 323728 332324 323734 332376
rect 546310 332324 546316 332376
rect 546368 332364 546374 332376
rect 568666 332364 568672 332376
rect 546368 332336 568672 332364
rect 546368 332324 546374 332336
rect 568666 332324 568672 332336
rect 568724 332324 568730 332376
rect 23014 332256 23020 332308
rect 23072 332296 23078 332308
rect 33226 332296 33232 332308
rect 23072 332268 33232 332296
rect 23072 332256 23078 332268
rect 33226 332256 33232 332268
rect 33284 332256 33290 332308
rect 266262 332256 266268 332308
rect 266320 332296 266326 332308
rect 290274 332296 290280 332308
rect 266320 332268 290280 332296
rect 266320 332256 266326 332268
rect 290274 332256 290280 332268
rect 290332 332256 290338 332308
rect 302050 332256 302056 332308
rect 302108 332296 302114 332308
rect 313550 332296 313556 332308
rect 302108 332268 313556 332296
rect 302108 332256 302114 332268
rect 313550 332256 313556 332268
rect 313608 332256 313614 332308
rect 21726 332188 21732 332240
rect 21784 332228 21790 332240
rect 23658 332228 23664 332240
rect 21784 332200 23664 332228
rect 21784 332188 21790 332200
rect 23658 332188 23664 332200
rect 23716 332188 23722 332240
rect 281350 332188 281356 332240
rect 281408 332228 281414 332240
rect 285674 332228 285680 332240
rect 281408 332200 285680 332228
rect 281408 332188 281414 332200
rect 285674 332188 285680 332200
rect 285732 332188 285738 332240
rect 308490 332188 308496 332240
rect 308548 332228 308554 332240
rect 580534 332228 580540 332240
rect 308548 332200 580540 332228
rect 308548 332188 308554 332200
rect 580534 332188 580540 332200
rect 580592 332188 580598 332240
rect 300394 332120 300400 332172
rect 300452 332160 300458 332172
rect 311250 332160 311256 332172
rect 300452 332132 311256 332160
rect 300452 332120 300458 332132
rect 311250 332120 311256 332132
rect 311308 332120 311314 332172
rect 21818 331984 21824 332036
rect 21876 332024 21882 332036
rect 22738 332024 22744 332036
rect 21876 331996 22744 332024
rect 21876 331984 21882 331996
rect 22738 331984 22744 331996
rect 22796 331984 22802 332036
rect 190362 331916 190368 331968
rect 190420 331956 190426 331968
rect 192110 331956 192116 331968
rect 190420 331928 192116 331956
rect 190420 331916 190426 331928
rect 192110 331916 192116 331928
rect 192168 331916 192174 331968
rect 561490 331916 561496 331968
rect 561548 331956 561554 331968
rect 568758 331956 568764 331968
rect 561548 331928 568764 331956
rect 561548 331916 561554 331928
rect 568758 331916 568764 331928
rect 568816 331956 568822 331968
rect 570230 331956 570236 331968
rect 568816 331928 570236 331956
rect 568816 331916 568822 331928
rect 570230 331916 570236 331928
rect 570288 331916 570294 331968
rect 22094 331848 22100 331900
rect 22152 331888 22158 331900
rect 22738 331888 22744 331900
rect 22152 331860 22744 331888
rect 22152 331848 22158 331860
rect 22738 331848 22744 331860
rect 22796 331888 22802 331900
rect 53466 331888 53472 331900
rect 22796 331860 53472 331888
rect 22796 331848 22802 331860
rect 53466 331848 53472 331860
rect 53524 331848 53530 331900
rect 185670 331848 185676 331900
rect 185728 331888 185734 331900
rect 187602 331888 187608 331900
rect 185728 331860 187608 331888
rect 185728 331848 185734 331860
rect 187602 331848 187608 331860
rect 187660 331848 187666 331900
rect 282178 331848 282184 331900
rect 282236 331888 282242 331900
rect 289078 331888 289084 331900
rect 282236 331860 289084 331888
rect 282236 331848 282242 331860
rect 289078 331848 289084 331860
rect 289136 331888 289142 331900
rect 292574 331888 292580 331900
rect 289136 331860 292580 331888
rect 289136 331848 289142 331860
rect 292574 331848 292580 331860
rect 292632 331848 292638 331900
rect 556430 331848 556436 331900
rect 556488 331888 556494 331900
rect 569954 331888 569960 331900
rect 556488 331860 569960 331888
rect 556488 331848 556494 331860
rect 569954 331848 569960 331860
rect 570012 331848 570018 331900
rect 299014 331304 299020 331356
rect 299072 331344 299078 331356
rect 302142 331344 302148 331356
rect 299072 331316 302148 331344
rect 299072 331304 299078 331316
rect 302142 331304 302148 331316
rect 302200 331304 302206 331356
rect 21910 331236 21916 331288
rect 21968 331276 21974 331288
rect 22830 331276 22836 331288
rect 21968 331248 22836 331276
rect 21968 331236 21974 331248
rect 22830 331236 22836 331248
rect 22888 331236 22894 331288
rect 134426 331276 134432 331288
rect 132466 331248 134432 331276
rect 16298 331100 16304 331152
rect 16356 331140 16362 331152
rect 132466 331140 132494 331248
rect 134426 331236 134432 331248
rect 134484 331236 134490 331288
rect 170490 331236 170496 331288
rect 170548 331276 170554 331288
rect 171778 331276 171784 331288
rect 170548 331248 171784 331276
rect 170548 331236 170554 331248
rect 171778 331236 171784 331248
rect 171836 331276 171842 331288
rect 172330 331276 172336 331288
rect 171836 331248 172336 331276
rect 171836 331236 171842 331248
rect 172330 331236 172336 331248
rect 172388 331236 172394 331288
rect 173802 331236 173808 331288
rect 173860 331276 173866 331288
rect 174906 331276 174912 331288
rect 173860 331248 174912 331276
rect 173860 331236 173866 331248
rect 174906 331236 174912 331248
rect 174964 331236 174970 331288
rect 290274 331236 290280 331288
rect 290332 331276 290338 331288
rect 292666 331276 292672 331288
rect 290332 331248 292672 331276
rect 290332 331236 290338 331248
rect 292666 331236 292672 331248
rect 292724 331236 292730 331288
rect 301958 331236 301964 331288
rect 302016 331276 302022 331288
rect 303062 331276 303068 331288
rect 302016 331248 303068 331276
rect 302016 331236 302022 331248
rect 303062 331236 303068 331248
rect 303120 331236 303126 331288
rect 352558 331236 352564 331288
rect 352616 331276 352622 331288
rect 354030 331276 354036 331288
rect 352616 331248 354036 331276
rect 352616 331236 352622 331248
rect 354030 331236 354036 331248
rect 354088 331236 354094 331288
rect 404630 331236 404636 331288
rect 404688 331276 404694 331288
rect 405734 331276 405740 331288
rect 404688 331248 405740 331276
rect 404688 331236 404694 331248
rect 405734 331236 405740 331248
rect 405792 331236 405798 331288
rect 465350 331236 465356 331288
rect 465408 331276 465414 331288
rect 467098 331276 467104 331288
rect 465408 331248 467104 331276
rect 465408 331236 465414 331248
rect 467098 331236 467104 331248
rect 467156 331236 467162 331288
rect 160094 331168 160100 331220
rect 160152 331208 160158 331220
rect 291378 331208 291384 331220
rect 160152 331180 291384 331208
rect 160152 331168 160158 331180
rect 291378 331168 291384 331180
rect 291436 331168 291442 331220
rect 293862 331168 293868 331220
rect 293920 331208 293926 331220
rect 296714 331208 296720 331220
rect 293920 331180 296720 331208
rect 293920 331168 293926 331180
rect 296714 331168 296720 331180
rect 296772 331208 296778 331220
rect 394510 331208 394516 331220
rect 296772 331180 394516 331208
rect 296772 331168 296778 331180
rect 394510 331168 394516 331180
rect 394568 331168 394574 331220
rect 434990 331168 434996 331220
rect 435048 331208 435054 331220
rect 565814 331208 565820 331220
rect 435048 331180 565820 331208
rect 435048 331168 435054 331180
rect 565814 331168 565820 331180
rect 565872 331168 565878 331220
rect 16356 331112 132494 331140
rect 16356 331100 16362 331112
rect 172330 331100 172336 331152
rect 172388 331140 172394 331152
rect 285766 331140 285772 331152
rect 172388 331112 285772 331140
rect 172388 331100 172394 331112
rect 285766 331100 285772 331112
rect 285824 331100 285830 331152
rect 17678 331032 17684 331084
rect 17736 331072 17742 331084
rect 119246 331072 119252 331084
rect 17736 331044 119252 331072
rect 17736 331032 17742 331044
rect 119246 331032 119252 331044
rect 119304 331032 119310 331084
rect 220814 331032 220820 331084
rect 220872 331072 220878 331084
rect 292850 331072 292856 331084
rect 220872 331044 292856 331072
rect 220872 331032 220878 331044
rect 292850 331032 292856 331044
rect 292908 331032 292914 331084
rect 23382 330964 23388 331016
rect 23440 331004 23446 331016
rect 99006 331004 99012 331016
rect 23440 330976 99012 331004
rect 23440 330964 23446 330976
rect 99006 330964 99012 330976
rect 99064 330964 99070 331016
rect 19150 330896 19156 330948
rect 19208 330936 19214 330948
rect 154666 330936 154672 330948
rect 19208 330908 154672 330936
rect 19208 330896 19214 330908
rect 154666 330896 154672 330908
rect 154724 330896 154730 330948
rect 112438 330828 112444 330880
rect 112496 330868 112502 330880
rect 114186 330868 114192 330880
rect 112496 330840 114192 330868
rect 112496 330828 112502 330840
rect 114186 330828 114192 330840
rect 114244 330828 114250 330880
rect 292850 330692 292856 330744
rect 292908 330732 292914 330744
rect 294138 330732 294144 330744
rect 292908 330704 294144 330732
rect 292908 330692 292914 330704
rect 294138 330692 294144 330704
rect 294196 330692 294202 330744
rect 18966 330624 18972 330676
rect 19024 330664 19030 330676
rect 19150 330664 19156 330676
rect 19024 330636 19156 330664
rect 19024 330624 19030 330636
rect 19150 330624 19156 330636
rect 19208 330624 19214 330676
rect 187602 330556 187608 330608
rect 187660 330596 187666 330608
rect 285490 330596 285496 330608
rect 187660 330568 285496 330596
rect 187660 330556 187666 330568
rect 285490 330556 285496 330568
rect 285548 330556 285554 330608
rect 192110 330488 192116 330540
rect 192168 330528 192174 330540
rect 291378 330528 291384 330540
rect 192168 330500 291384 330528
rect 192168 330488 192174 330500
rect 291378 330488 291384 330500
rect 291436 330528 291442 330540
rect 293954 330528 293960 330540
rect 291436 330500 293960 330528
rect 291436 330488 291442 330500
rect 293954 330488 293960 330500
rect 294012 330488 294018 330540
rect 303614 330488 303620 330540
rect 303672 330528 303678 330540
rect 414750 330528 414756 330540
rect 303672 330500 414756 330528
rect 303672 330488 303678 330500
rect 414750 330488 414756 330500
rect 414808 330488 414814 330540
rect 565814 330488 565820 330540
rect 565872 330528 565878 330540
rect 568850 330528 568856 330540
rect 565872 330500 568856 330528
rect 565872 330488 565878 330500
rect 568850 330488 568856 330500
rect 568908 330528 568914 330540
rect 572898 330528 572904 330540
rect 568908 330500 572904 330528
rect 568908 330488 568914 330500
rect 572898 330488 572904 330500
rect 572956 330488 572962 330540
rect 285490 329944 285496 329996
rect 285548 329984 285554 329996
rect 286870 329984 286876 329996
rect 285548 329956 286876 329984
rect 285548 329944 285554 329956
rect 286870 329944 286876 329956
rect 286928 329944 286934 329996
rect 17586 329740 17592 329792
rect 17644 329780 17650 329792
rect 17770 329780 17776 329792
rect 17644 329752 17776 329780
rect 17644 329740 17650 329752
rect 17770 329740 17776 329752
rect 17828 329780 17834 329792
rect 104066 329780 104072 329792
rect 17828 329752 104072 329780
rect 17828 329740 17834 329752
rect 104066 329740 104072 329752
rect 104124 329740 104130 329792
rect 294046 329740 294052 329792
rect 294104 329780 294110 329792
rect 295334 329780 295340 329792
rect 294104 329752 295340 329780
rect 294104 329740 294110 329752
rect 295334 329740 295340 329752
rect 295392 329740 295398 329792
rect 296530 329740 296536 329792
rect 296588 329780 296594 329792
rect 297726 329780 297732 329792
rect 296588 329752 297732 329780
rect 296588 329740 296594 329752
rect 297726 329740 297732 329752
rect 297784 329740 297790 329792
rect 299198 329740 299204 329792
rect 299256 329780 299262 329792
rect 300762 329780 300768 329792
rect 299256 329752 300768 329780
rect 299256 329740 299262 329752
rect 300762 329740 300768 329752
rect 300820 329740 300826 329792
rect 301774 329740 301780 329792
rect 301832 329780 301838 329792
rect 302142 329780 302148 329792
rect 301832 329752 302148 329780
rect 301832 329740 301838 329752
rect 302142 329740 302148 329752
rect 302200 329740 302206 329792
rect 302234 329740 302240 329792
rect 302292 329780 302298 329792
rect 373902 329780 373908 329792
rect 302292 329752 373908 329780
rect 302292 329740 302298 329752
rect 373902 329740 373908 329752
rect 373960 329740 373966 329792
rect 440234 329740 440240 329792
rect 440292 329780 440298 329792
rect 571610 329780 571616 329792
rect 440292 329752 571616 329780
rect 440292 329740 440298 329752
rect 571610 329740 571616 329752
rect 571668 329740 571674 329792
rect 19058 329672 19064 329724
rect 19116 329712 19122 329724
rect 58526 329712 58532 329724
rect 19116 329684 58532 329712
rect 19116 329672 19122 329684
rect 58526 329672 58532 329684
rect 58584 329672 58590 329724
rect 300780 329644 300808 329740
rect 302160 329712 302188 329740
rect 343910 329712 343916 329724
rect 302160 329684 343916 329712
rect 343910 329672 343916 329684
rect 343968 329672 343974 329724
rect 338850 329644 338856 329656
rect 300780 329616 338856 329644
rect 338850 329604 338856 329616
rect 338908 329604 338914 329656
rect 299106 329536 299112 329588
rect 299164 329576 299170 329588
rect 302234 329576 302240 329588
rect 299164 329548 302240 329576
rect 299164 329536 299170 329548
rect 302234 329536 302240 329548
rect 302292 329536 302298 329588
rect 195974 329060 195980 329112
rect 196032 329100 196038 329112
rect 294046 329100 294052 329112
rect 196032 329072 294052 329100
rect 196032 329060 196038 329072
rect 294046 329060 294052 329072
rect 294104 329060 294110 329112
rect 297726 329060 297732 329112
rect 297784 329100 297790 329112
rect 297910 329100 297916 329112
rect 297784 329072 297916 329100
rect 297784 329060 297790 329072
rect 297910 329060 297916 329072
rect 297968 329100 297974 329112
rect 399570 329100 399576 329112
rect 297968 329072 399576 329100
rect 297968 329060 297974 329072
rect 399570 329060 399576 329072
rect 399628 329060 399634 329112
rect 289078 319404 289084 319456
rect 289136 319444 289142 319456
rect 424318 319444 424324 319456
rect 289136 319416 424324 319444
rect 289136 319404 289142 319416
rect 424318 319404 424324 319416
rect 424376 319404 424382 319456
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 10318 318832 10324 318844
rect 3384 318804 10324 318832
rect 3384 318792 3390 318804
rect 10318 318792 10324 318804
rect 10376 318792 10382 318844
rect 164234 318724 164240 318776
rect 164292 318764 164298 318776
rect 284202 318764 284208 318776
rect 164292 318736 284208 318764
rect 164292 318724 164298 318736
rect 284202 318724 284208 318736
rect 284260 318724 284266 318776
rect 303062 318724 303068 318776
rect 303120 318764 303126 318776
rect 303706 318764 303712 318776
rect 303120 318736 303712 318764
rect 303120 318724 303126 318736
rect 303706 318724 303712 318736
rect 303764 318764 303770 318776
rect 408494 318764 408500 318776
rect 303764 318736 408500 318764
rect 303764 318724 303770 318736
rect 408494 318724 408500 318736
rect 408552 318724 408558 318776
rect 449894 318724 449900 318776
rect 449952 318764 449958 318776
rect 567654 318764 567660 318776
rect 449952 318736 567660 318764
rect 449952 318724 449958 318736
rect 567654 318724 567660 318736
rect 567712 318724 567718 318776
rect 459554 318656 459560 318708
rect 459612 318696 459618 318708
rect 575474 318696 575480 318708
rect 459612 318668 575480 318696
rect 459612 318656 459618 318668
rect 575474 318656 575480 318668
rect 575532 318656 575538 318708
rect 489914 318588 489920 318640
rect 489972 318628 489978 318640
rect 575566 318628 575572 318640
rect 489972 318600 575572 318628
rect 489972 318588 489978 318600
rect 575566 318588 575572 318600
rect 575624 318588 575630 318640
rect 304258 318044 304264 318096
rect 304316 318084 304322 318096
rect 305178 318084 305184 318096
rect 304316 318056 305184 318084
rect 304316 318044 304322 318056
rect 305178 318044 305184 318056
rect 305236 318084 305242 318096
rect 405734 318084 405740 318096
rect 305236 318056 405740 318084
rect 305236 318044 305242 318056
rect 405734 318044 405740 318056
rect 405792 318044 405798 318096
rect 469214 318044 469220 318096
rect 469272 318084 469278 318096
rect 573358 318084 573364 318096
rect 469272 318056 573364 318084
rect 469272 318044 469278 318056
rect 573358 318044 573364 318056
rect 573416 318044 573422 318096
rect 173802 317364 173808 317416
rect 173860 317404 173866 317416
rect 285398 317404 285404 317416
rect 173860 317376 285404 317404
rect 173860 317364 173866 317376
rect 285398 317364 285404 317376
rect 285456 317364 285462 317416
rect 573358 317364 573364 317416
rect 573416 317404 573422 317416
rect 574094 317404 574100 317416
rect 573416 317376 574100 317404
rect 573416 317364 573422 317376
rect 574094 317364 574100 317376
rect 574152 317364 574158 317416
rect 300578 316004 300584 316056
rect 300636 316044 300642 316056
rect 306374 316044 306380 316056
rect 300636 316016 306380 316044
rect 300636 316004 300642 316016
rect 306374 316004 306380 316016
rect 306432 316004 306438 316056
rect 571518 316004 571524 316056
rect 571576 316004 571582 316056
rect 16390 315936 16396 315988
rect 16448 315976 16454 315988
rect 17218 315976 17224 315988
rect 16448 315948 17224 315976
rect 16448 315936 16454 315948
rect 17218 315936 17224 315948
rect 17276 315976 17282 315988
rect 112438 315976 112444 315988
rect 17276 315948 112444 315976
rect 17276 315936 17282 315948
rect 112438 315936 112444 315948
rect 112496 315936 112502 315988
rect 179414 315936 179420 315988
rect 179472 315976 179478 315988
rect 285582 315976 285588 315988
rect 179472 315948 285588 315976
rect 179472 315936 179478 315948
rect 285582 315936 285588 315948
rect 285640 315936 285646 315988
rect 306392 315976 306420 316004
rect 378134 315976 378140 315988
rect 306392 315948 378140 315976
rect 378134 315936 378140 315948
rect 378192 315936 378198 315988
rect 505094 315936 505100 315988
rect 505152 315976 505158 315988
rect 566366 315976 566372 315988
rect 505152 315948 566372 315976
rect 505152 315936 505158 315948
rect 566366 315936 566372 315948
rect 566424 315976 566430 315988
rect 567102 315976 567108 315988
rect 566424 315948 567108 315976
rect 566424 315936 566430 315948
rect 567102 315936 567108 315948
rect 567160 315936 567166 315988
rect 571536 315976 571564 316004
rect 572806 315976 572812 315988
rect 571536 315948 572812 315976
rect 571536 315920 571564 315948
rect 572806 315936 572812 315948
rect 572864 315936 572870 315988
rect 22002 315868 22008 315920
rect 22060 315908 22066 315920
rect 82814 315908 82820 315920
rect 22060 315880 82820 315908
rect 22060 315868 22066 315880
rect 82814 315868 82820 315880
rect 82872 315868 82878 315920
rect 215202 315868 215208 315920
rect 215260 315908 215266 315920
rect 288526 315908 288532 315920
rect 215260 315880 288532 315908
rect 215260 315868 215266 315880
rect 288526 315868 288532 315880
rect 288584 315868 288590 315920
rect 296530 315868 296536 315920
rect 296588 315908 296594 315920
rect 298002 315908 298008 315920
rect 296588 315880 298008 315908
rect 296588 315868 296594 315880
rect 298002 315868 298008 315880
rect 298060 315908 298066 315920
rect 368474 315908 368480 315920
rect 298060 315880 368480 315908
rect 298060 315868 298066 315880
rect 368474 315868 368480 315880
rect 368532 315868 368538 315920
rect 510614 315868 510620 315920
rect 510672 315908 510678 315920
rect 570138 315908 570144 315920
rect 510672 315880 570144 315908
rect 510672 315868 510678 315880
rect 570138 315868 570144 315880
rect 570196 315868 570202 315920
rect 571518 315868 571524 315920
rect 571576 315868 571582 315920
rect 20622 315800 20628 315852
rect 20680 315840 20686 315852
rect 73154 315840 73160 315852
rect 20680 315812 73160 315840
rect 20680 315800 20686 315812
rect 73154 315800 73160 315812
rect 73212 315800 73218 315852
rect 224954 315800 224960 315852
rect 225012 315840 225018 315852
rect 287514 315840 287520 315852
rect 225012 315812 287520 315840
rect 225012 315800 225018 315812
rect 287514 315800 287520 315812
rect 287572 315800 287578 315852
rect 303246 315800 303252 315852
rect 303304 315840 303310 315852
rect 362954 315840 362960 315852
rect 303304 315812 362960 315840
rect 303304 315800 303310 315812
rect 362954 315800 362960 315812
rect 363012 315800 363018 315852
rect 514754 315800 514760 315852
rect 514812 315840 514818 315852
rect 572714 315840 572720 315852
rect 514812 315812 572720 315840
rect 514812 315800 514818 315812
rect 572714 315800 572720 315812
rect 572772 315800 572778 315852
rect 234614 315732 234620 315784
rect 234672 315772 234678 315784
rect 291194 315772 291200 315784
rect 234672 315744 291200 315772
rect 234672 315732 234678 315744
rect 291194 315732 291200 315744
rect 291252 315732 291258 315784
rect 298922 315732 298928 315784
rect 298980 315772 298986 315784
rect 358814 315772 358820 315784
rect 298980 315744 358820 315772
rect 298980 315732 298986 315744
rect 358814 315732 358820 315744
rect 358872 315732 358878 315784
rect 520274 315732 520280 315784
rect 520332 315772 520338 315784
rect 567746 315772 567752 315784
rect 520332 315744 567752 315772
rect 520332 315732 520338 315744
rect 567746 315732 567752 315744
rect 567804 315732 567810 315784
rect 299382 315664 299388 315716
rect 299440 315704 299446 315716
rect 352558 315704 352564 315716
rect 299440 315676 352564 315704
rect 299440 315664 299446 315676
rect 352558 315664 352564 315676
rect 352616 315664 352622 315716
rect 525794 315664 525800 315716
rect 525852 315704 525858 315716
rect 570046 315704 570052 315716
rect 525852 315676 570052 315704
rect 525852 315664 525858 315676
rect 570046 315664 570052 315676
rect 570104 315664 570110 315716
rect 300302 315596 300308 315648
rect 300360 315636 300366 315648
rect 347774 315636 347780 315648
rect 300360 315608 347780 315636
rect 300360 315596 300366 315608
rect 347774 315596 347780 315608
rect 347832 315596 347838 315648
rect 529934 315596 529940 315648
rect 529992 315636 529998 315648
rect 571518 315636 571524 315648
rect 529992 315608 571524 315636
rect 529992 315596 529998 315608
rect 571518 315596 571524 315608
rect 571576 315596 571582 315648
rect 285582 315392 285588 315444
rect 285640 315432 285646 315444
rect 290090 315432 290096 315444
rect 285640 315404 290096 315432
rect 285640 315392 285646 315404
rect 290090 315392 290096 315404
rect 290148 315392 290154 315444
rect 276014 315324 276020 315376
rect 276072 315364 276078 315376
rect 295978 315364 295984 315376
rect 276072 315336 295984 315364
rect 276072 315324 276078 315336
rect 295978 315324 295984 315336
rect 296036 315324 296042 315376
rect 93854 315296 93860 315308
rect 26206 315268 93860 315296
rect 18782 315188 18788 315240
rect 18840 315228 18846 315240
rect 19334 315228 19340 315240
rect 18840 315200 19340 315228
rect 18840 315188 18846 315200
rect 19334 315188 19340 315200
rect 19392 315228 19398 315240
rect 26206 315228 26234 315268
rect 93854 315256 93860 315268
rect 93912 315256 93918 315308
rect 270494 315256 270500 315308
rect 270552 315296 270558 315308
rect 297358 315296 297364 315308
rect 270552 315268 297364 315296
rect 270552 315256 270558 315268
rect 297358 315256 297364 315268
rect 297416 315256 297422 315308
rect 19392 315200 26234 315228
rect 19392 315188 19398 315200
rect 297818 314644 297824 314696
rect 297876 314684 297882 314696
rect 298922 314684 298928 314696
rect 297876 314656 298928 314684
rect 297876 314644 297882 314656
rect 298922 314644 298928 314656
rect 298980 314644 298986 314696
rect 299106 314644 299112 314696
rect 299164 314684 299170 314696
rect 300302 314684 300308 314696
rect 299164 314656 300308 314684
rect 299164 314644 299170 314656
rect 300302 314644 300308 314656
rect 300360 314644 300366 314696
rect 567746 314644 567752 314696
rect 567804 314684 567810 314696
rect 568758 314684 568764 314696
rect 567804 314656 568764 314684
rect 567804 314644 567810 314656
rect 568758 314644 568764 314656
rect 568816 314644 568822 314696
rect 570138 314644 570144 314696
rect 570196 314684 570202 314696
rect 571518 314684 571524 314696
rect 570196 314656 571524 314684
rect 570196 314644 570202 314656
rect 571518 314644 571524 314656
rect 571576 314644 571582 314696
rect 304994 314576 305000 314628
rect 305052 314616 305058 314628
rect 389174 314616 389180 314628
rect 305052 314588 389180 314616
rect 305052 314576 305058 314588
rect 389174 314576 389180 314588
rect 389232 314576 389238 314628
rect 454034 314576 454040 314628
rect 454092 314616 454098 314628
rect 565722 314616 565728 314628
rect 454092 314588 565728 314616
rect 454092 314576 454098 314588
rect 565722 314576 565728 314588
rect 565780 314576 565786 314628
rect 467098 314508 467104 314560
rect 467156 314548 467162 314560
rect 568850 314548 568856 314560
rect 467156 314520 568856 314548
rect 467156 314508 467162 314520
rect 568850 314508 568856 314520
rect 568908 314548 568914 314560
rect 570322 314548 570328 314560
rect 568908 314520 570328 314548
rect 568908 314508 568914 314520
rect 570322 314508 570328 314520
rect 570380 314508 570386 314560
rect 565722 314168 565728 314220
rect 565780 314208 565786 314220
rect 568850 314208 568856 314220
rect 565780 314180 568856 314208
rect 565780 314168 565786 314180
rect 568850 314168 568856 314180
rect 568908 314168 568914 314220
rect 285490 314032 285496 314084
rect 285548 314072 285554 314084
rect 292758 314072 292764 314084
rect 285548 314044 292764 314072
rect 285548 314032 285554 314044
rect 292758 314032 292764 314044
rect 292816 314032 292822 314084
rect 284294 313964 284300 314016
rect 284352 314004 284358 314016
rect 296714 314004 296720 314016
rect 284352 313976 296720 314004
rect 284352 313964 284358 313976
rect 296714 313964 296720 313976
rect 296772 313964 296778 314016
rect 305086 314004 305092 314016
rect 298848 313976 305092 314004
rect 200114 313896 200120 313948
rect 200172 313936 200178 313948
rect 288618 313936 288624 313948
rect 200172 313908 288624 313936
rect 200172 313896 200178 313908
rect 288618 313896 288624 313908
rect 288676 313896 288682 313948
rect 296438 313896 296444 313948
rect 296496 313936 296502 313948
rect 298848 313936 298876 313976
rect 305086 313964 305092 313976
rect 305144 313964 305150 314016
rect 296496 313908 298876 313936
rect 296496 313896 296502 313908
rect 301866 313896 301872 313948
rect 301924 313936 301930 313948
rect 304994 313936 305000 313948
rect 301924 313908 305000 313936
rect 301924 313896 301930 313908
rect 304994 313896 305000 313908
rect 305052 313896 305058 313948
rect 300670 313828 300676 313880
rect 300728 313868 300734 313880
rect 303614 313868 303620 313880
rect 300728 313840 303620 313868
rect 300728 313828 300734 313840
rect 303614 313828 303620 313840
rect 303672 313828 303678 313880
rect 3326 266364 3332 266416
rect 3384 266404 3390 266416
rect 20898 266404 20904 266416
rect 3384 266376 20904 266404
rect 3384 266364 3390 266376
rect 20898 266364 20904 266376
rect 20956 266364 20962 266416
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 4890 240224 4896 240236
rect 2832 240196 4896 240224
rect 2832 240184 2838 240196
rect 4890 240184 4896 240196
rect 4948 240184 4954 240236
rect 12342 214548 12348 214600
rect 12400 214588 12406 214600
rect 13170 214588 13176 214600
rect 12400 214560 13176 214588
rect 12400 214548 12406 214560
rect 13170 214548 13176 214560
rect 13228 214548 13234 214600
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 13262 213976 13268 213988
rect 3384 213948 13268 213976
rect 3384 213936 3390 213948
rect 13262 213936 13268 213948
rect 13320 213936 13326 213988
rect 296438 206252 296444 206304
rect 296496 206292 296502 206304
rect 296496 206264 296714 206292
rect 296496 206252 296502 206264
rect 285490 205912 285496 205964
rect 285548 205952 285554 205964
rect 288618 205952 288624 205964
rect 285548 205924 288624 205952
rect 285548 205912 285554 205924
rect 288618 205912 288624 205924
rect 288676 205912 288682 205964
rect 296686 205952 296714 206264
rect 303614 205952 303620 205964
rect 296686 205924 303620 205952
rect 303614 205912 303620 205924
rect 303672 205912 303678 205964
rect 568022 205640 568028 205692
rect 568080 205680 568086 205692
rect 578234 205680 578240 205692
rect 568080 205652 578240 205680
rect 568080 205640 568086 205652
rect 578234 205640 578240 205652
rect 578292 205640 578298 205692
rect 285582 204892 285588 204944
rect 285640 204932 285646 204944
rect 291378 204932 291384 204944
rect 285640 204904 291384 204932
rect 285640 204892 285646 204904
rect 291378 204892 291384 204904
rect 291436 204892 291442 204944
rect 293862 204892 293868 204944
rect 293920 204932 293926 204944
rect 305086 204932 305092 204944
rect 293920 204904 305092 204932
rect 293920 204892 293926 204904
rect 305086 204892 305092 204904
rect 305144 204892 305150 204944
rect 526346 204892 526352 204944
rect 526404 204932 526410 204944
rect 570046 204932 570052 204944
rect 526404 204904 570052 204932
rect 526404 204892 526410 204904
rect 570046 204892 570052 204904
rect 570104 204932 570110 204944
rect 572898 204932 572904 204944
rect 570104 204904 572904 204932
rect 570104 204892 570110 204904
rect 572898 204892 572904 204904
rect 572956 204892 572962 204944
rect 297818 204824 297824 204876
rect 297876 204864 297882 204876
rect 301774 204864 301780 204876
rect 297876 204836 301780 204864
rect 297876 204824 297882 204836
rect 301774 204824 301780 204836
rect 301832 204824 301838 204876
rect 298002 204756 298008 204808
rect 298060 204796 298066 204808
rect 299382 204796 299388 204808
rect 298060 204768 299388 204796
rect 298060 204756 298066 204768
rect 299382 204756 299388 204768
rect 299440 204756 299446 204808
rect 572714 204756 572720 204808
rect 572772 204796 572778 204808
rect 574278 204796 574284 204808
rect 572772 204768 574284 204796
rect 572772 204756 572778 204768
rect 574278 204756 574284 204768
rect 574336 204756 574342 204808
rect 17494 204688 17500 204740
rect 17552 204728 17558 204740
rect 18966 204728 18972 204740
rect 17552 204700 18972 204728
rect 17552 204688 17558 204700
rect 18966 204688 18972 204700
rect 19024 204688 19030 204740
rect 14826 204552 14832 204604
rect 14884 204592 14890 204604
rect 180242 204592 180248 204604
rect 14884 204564 180248 204592
rect 14884 204552 14890 204564
rect 180242 204552 180248 204564
rect 180300 204592 180306 204604
rect 180300 204564 180794 204592
rect 180300 204552 180306 204564
rect 16298 204484 16304 204536
rect 16356 204524 16362 204536
rect 18782 204524 18788 204536
rect 16356 204496 18788 204524
rect 16356 204484 16362 204496
rect 18782 204484 18788 204496
rect 18840 204524 18846 204536
rect 134426 204524 134432 204536
rect 18840 204496 134432 204524
rect 18840 204484 18846 204496
rect 134426 204484 134432 204496
rect 134484 204484 134490 204536
rect 17678 204416 17684 204468
rect 17736 204456 17742 204468
rect 119246 204456 119252 204468
rect 17736 204428 119252 204456
rect 17736 204416 17742 204428
rect 119246 204416 119252 204428
rect 119304 204416 119310 204468
rect 18966 204348 18972 204400
rect 19024 204388 19030 204400
rect 154666 204388 154672 204400
rect 19024 204360 154672 204388
rect 19024 204348 19030 204360
rect 154666 204348 154672 204360
rect 154724 204348 154730 204400
rect 180766 204320 180794 204564
rect 246390 204552 246396 204604
rect 246448 204592 246454 204604
rect 290182 204592 290188 204604
rect 246448 204564 290188 204592
rect 246448 204552 246454 204564
rect 290182 204552 290188 204564
rect 290240 204592 290246 204604
rect 292850 204592 292856 204604
rect 290240 204564 292856 204592
rect 290240 204552 290246 204564
rect 292850 204552 292856 204564
rect 292908 204552 292914 204604
rect 299382 204552 299388 204604
rect 299440 204592 299446 204604
rect 354030 204592 354036 204604
rect 299440 204564 354036 204592
rect 299440 204552 299446 204564
rect 354030 204552 354036 204564
rect 354088 204552 354094 204604
rect 531498 204552 531504 204604
rect 531556 204592 531562 204604
rect 572806 204592 572812 204604
rect 531556 204564 572812 204592
rect 531556 204552 531562 204564
rect 572806 204552 572812 204564
rect 572864 204552 572870 204604
rect 241330 204484 241336 204536
rect 241388 204524 241394 204536
rect 289906 204524 289912 204536
rect 241388 204496 289912 204524
rect 241388 204484 241394 204496
rect 289906 204484 289912 204496
rect 289964 204484 289970 204536
rect 301774 204484 301780 204536
rect 301832 204524 301838 204536
rect 359090 204524 359096 204536
rect 301832 204496 359096 204524
rect 301832 204484 301838 204496
rect 359090 204484 359096 204496
rect 359148 204484 359154 204536
rect 521654 204484 521660 204536
rect 521712 204524 521718 204536
rect 567654 204524 567660 204536
rect 521712 204496 567660 204524
rect 521712 204484 521718 204496
rect 567654 204484 567660 204496
rect 567712 204524 567718 204536
rect 568758 204524 568764 204536
rect 567712 204496 568764 204524
rect 567712 204484 567718 204496
rect 568758 204484 568764 204496
rect 568816 204484 568822 204536
rect 235902 204416 235908 204468
rect 235960 204456 235966 204468
rect 287882 204456 287888 204468
rect 235960 204428 287888 204456
rect 235960 204416 235966 204428
rect 287882 204416 287888 204428
rect 287940 204456 287946 204468
rect 291194 204456 291200 204468
rect 287940 204428 291200 204456
rect 287940 204416 287946 204428
rect 291194 204416 291200 204428
rect 291252 204416 291258 204468
rect 300578 204416 300584 204468
rect 300636 204456 300642 204468
rect 303890 204456 303896 204468
rect 300636 204428 303896 204456
rect 300636 204416 300642 204428
rect 303890 204416 303896 204428
rect 303948 204456 303954 204468
rect 379330 204456 379336 204468
rect 303948 204428 379336 204456
rect 303948 204416 303954 204428
rect 379330 204416 379336 204428
rect 379388 204416 379394 204468
rect 515950 204416 515956 204468
rect 516008 204456 516014 204468
rect 572714 204456 572720 204468
rect 516008 204428 572720 204456
rect 516008 204416 516014 204428
rect 572714 204416 572720 204428
rect 572772 204416 572778 204468
rect 220722 204348 220728 204400
rect 220780 204388 220786 204400
rect 293954 204388 293960 204400
rect 220780 204360 293960 204388
rect 220780 204348 220786 204360
rect 293954 204348 293960 204360
rect 294012 204348 294018 204400
rect 300762 204388 300768 204400
rect 300688 204360 300768 204388
rect 290090 204320 290096 204332
rect 180766 204292 290096 204320
rect 290090 204280 290096 204292
rect 290148 204280 290154 204332
rect 20438 204212 20444 204264
rect 20496 204252 20502 204264
rect 20622 204252 20628 204264
rect 20496 204224 20628 204252
rect 20496 204212 20502 204224
rect 20622 204212 20628 204224
rect 20680 204212 20686 204264
rect 88886 204252 88892 204264
rect 21468 204224 88892 204252
rect 18874 204144 18880 204196
rect 18932 204184 18938 204196
rect 21468 204184 21496 204224
rect 88886 204212 88892 204224
rect 88944 204212 88950 204264
rect 144822 204212 144828 204264
rect 144880 204252 144886 204264
rect 149606 204252 149612 204264
rect 144880 204224 149612 204252
rect 144880 204212 144886 204224
rect 149606 204212 149612 204224
rect 149664 204212 149670 204264
rect 173894 204212 173900 204264
rect 173952 204252 173958 204264
rect 175182 204252 175188 204264
rect 173952 204224 175188 204252
rect 173952 204212 173958 204224
rect 175182 204212 175188 204224
rect 175240 204212 175246 204264
rect 251082 204212 251088 204264
rect 251140 204252 251146 204264
rect 251140 204224 287054 204252
rect 251140 204212 251146 204224
rect 18932 204156 21496 204184
rect 18932 204144 18938 204156
rect 22002 204144 22008 204196
rect 22060 204184 22066 204196
rect 83826 204184 83832 204196
rect 22060 204156 83832 204184
rect 22060 204144 22066 204156
rect 83826 204144 83832 204156
rect 83884 204144 83890 204196
rect 256510 204144 256516 204196
rect 256568 204184 256574 204196
rect 285674 204184 285680 204196
rect 256568 204156 285680 204184
rect 256568 204144 256574 204156
rect 285674 204144 285680 204156
rect 285732 204144 285738 204196
rect 20346 204076 20352 204128
rect 20404 204116 20410 204128
rect 78766 204116 78772 204128
rect 20404 204088 78772 204116
rect 20404 204076 20410 204088
rect 78766 204076 78772 204088
rect 78824 204076 78830 204128
rect 190362 204076 190368 204128
rect 190420 204116 190426 204128
rect 192478 204116 192484 204128
rect 190420 204088 192484 204116
rect 190420 204076 190426 204088
rect 192478 204076 192484 204088
rect 192536 204076 192542 204128
rect 287026 204116 287054 204224
rect 291194 204212 291200 204264
rect 291252 204252 291258 204264
rect 292574 204252 292580 204264
rect 291252 204224 292580 204252
rect 291252 204212 291258 204224
rect 292574 204212 292580 204224
rect 292632 204212 292638 204264
rect 299014 204212 299020 204264
rect 299072 204252 299078 204264
rect 299290 204252 299296 204264
rect 299072 204224 299296 204252
rect 299072 204212 299078 204224
rect 299290 204212 299296 204224
rect 299348 204212 299354 204264
rect 299382 204212 299388 204264
rect 299440 204252 299446 204264
rect 300688 204252 300716 204360
rect 300762 204348 300768 204360
rect 300820 204348 300826 204400
rect 301866 204348 301872 204400
rect 301924 204388 301930 204400
rect 304994 204388 305000 204400
rect 301924 204360 305000 204388
rect 301924 204348 301930 204360
rect 304994 204348 305000 204360
rect 305052 204388 305058 204400
rect 389450 204388 389456 204400
rect 305052 204360 389456 204388
rect 305052 204348 305058 204360
rect 389450 204348 389456 204360
rect 389508 204348 389514 204400
rect 510890 204348 510896 204400
rect 510948 204388 510954 204400
rect 571518 204388 571524 204400
rect 510948 204360 571524 204388
rect 510948 204348 510954 204360
rect 571518 204348 571524 204360
rect 571576 204348 571582 204400
rect 302878 204280 302884 204332
rect 302936 204320 302942 204332
rect 302936 204292 404676 204320
rect 302936 204280 302942 204292
rect 404648 204264 404676 204292
rect 505830 204280 505836 204332
rect 505888 204320 505894 204332
rect 567470 204320 567476 204332
rect 505888 204292 567476 204320
rect 505888 204280 505894 204292
rect 567470 204280 567476 204292
rect 567528 204320 567534 204332
rect 567746 204320 567752 204332
rect 567528 204292 567752 204320
rect 567528 204280 567534 204292
rect 567746 204280 567752 204292
rect 567804 204280 567810 204332
rect 299440 204224 300716 204252
rect 299440 204212 299446 204224
rect 291378 204144 291384 204196
rect 291436 204184 291442 204196
rect 292666 204184 292672 204196
rect 291436 204156 292672 204184
rect 291436 204144 291442 204156
rect 292666 204144 292672 204156
rect 292724 204144 292730 204196
rect 300688 204184 300716 204224
rect 300762 204212 300768 204264
rect 300820 204252 300826 204264
rect 302142 204252 302148 204264
rect 300820 204224 302148 204252
rect 300820 204212 300826 204224
rect 302142 204212 302148 204224
rect 302200 204252 302206 204264
rect 343910 204252 343916 204264
rect 302200 204224 343916 204252
rect 302200 204212 302206 204224
rect 343910 204212 343916 204224
rect 343968 204212 343974 204264
rect 404630 204212 404636 204264
rect 404688 204252 404694 204264
rect 405918 204252 405924 204264
rect 404688 204224 405924 204252
rect 404688 204212 404694 204224
rect 405918 204212 405924 204224
rect 405976 204212 405982 204264
rect 424318 204212 424324 204264
rect 424376 204252 424382 204264
rect 424870 204252 424876 204264
rect 424376 204224 424876 204252
rect 424376 204212 424382 204224
rect 424870 204212 424876 204224
rect 424928 204252 424934 204264
rect 429930 204252 429936 204264
rect 424928 204224 429936 204252
rect 424928 204212 424934 204224
rect 429930 204212 429936 204224
rect 429988 204212 429994 204264
rect 541250 204212 541256 204264
rect 541308 204252 541314 204264
rect 567562 204252 567568 204264
rect 541308 204224 567568 204252
rect 541308 204212 541314 204224
rect 567562 204212 567568 204224
rect 567620 204212 567626 204264
rect 333790 204184 333796 204196
rect 300688 204156 333796 204184
rect 333790 204144 333796 204156
rect 333848 204144 333854 204196
rect 546310 204144 546316 204196
rect 546368 204184 546374 204196
rect 568666 204184 568672 204196
rect 546368 204156 568672 204184
rect 546368 204144 546374 204156
rect 568666 204144 568672 204156
rect 568724 204144 568730 204196
rect 289814 204116 289820 204128
rect 287026 204088 289820 204116
rect 289814 204076 289820 204088
rect 289872 204116 289878 204128
rect 294046 204116 294052 204128
rect 289872 204088 294052 204116
rect 289872 204076 289878 204088
rect 294046 204076 294052 204088
rect 294104 204076 294110 204128
rect 299290 204076 299296 204128
rect 299348 204116 299354 204128
rect 328730 204116 328736 204128
rect 299348 204088 328736 204116
rect 299348 204076 299354 204088
rect 328730 204076 328736 204088
rect 328788 204076 328794 204128
rect 382274 204076 382280 204128
rect 382332 204116 382338 204128
rect 384390 204116 384396 204128
rect 382332 204088 384396 204116
rect 382332 204076 382338 204088
rect 384390 204076 384396 204088
rect 384448 204076 384454 204128
rect 470410 204076 470416 204128
rect 470468 204116 470474 204128
rect 471330 204116 471336 204128
rect 470468 204088 471336 204116
rect 470468 204076 470474 204088
rect 471330 204076 471336 204088
rect 471388 204076 471394 204128
rect 561490 204076 561496 204128
rect 561548 204116 561554 204128
rect 570230 204116 570236 204128
rect 561548 204088 570236 204116
rect 561548 204076 561554 204088
rect 570230 204076 570236 204088
rect 570288 204076 570294 204128
rect 20438 204008 20444 204060
rect 20496 204048 20502 204060
rect 73706 204048 73712 204060
rect 20496 204020 73712 204048
rect 20496 204008 20502 204020
rect 73706 204008 73712 204020
rect 73764 204008 73770 204060
rect 303154 204008 303160 204060
rect 303212 204048 303218 204060
rect 323670 204048 323676 204060
rect 303212 204020 323676 204048
rect 303212 204008 303218 204020
rect 323670 204008 323676 204020
rect 323728 204008 323734 204060
rect 4798 203940 4804 203992
rect 4856 203980 4862 203992
rect 4856 203952 20484 203980
rect 4856 203940 4862 203952
rect 19058 203872 19064 203924
rect 19116 203912 19122 203924
rect 20346 203912 20352 203924
rect 19116 203884 20352 203912
rect 19116 203872 19122 203884
rect 20346 203872 20352 203884
rect 20404 203872 20410 203924
rect 20456 203912 20484 203952
rect 23290 203940 23296 203992
rect 23348 203980 23354 203992
rect 33226 203980 33232 203992
rect 23348 203952 33232 203980
rect 23348 203940 23354 203952
rect 33226 203940 33232 203952
rect 33284 203940 33290 203992
rect 33318 203940 33324 203992
rect 33376 203980 33382 203992
rect 38286 203980 38292 203992
rect 33376 203952 38292 203980
rect 33376 203940 33382 203952
rect 38286 203940 38292 203952
rect 38344 203940 38350 203992
rect 301958 203940 301964 203992
rect 302016 203980 302022 203992
rect 318610 203980 318616 203992
rect 302016 203952 318616 203980
rect 302016 203940 302022 203952
rect 318610 203940 318616 203952
rect 318668 203940 318674 203992
rect 23382 203912 23388 203924
rect 20456 203884 23388 203912
rect 23382 203872 23388 203884
rect 23440 203872 23446 203924
rect 281442 203872 281448 203924
rect 281500 203912 281506 203924
rect 287698 203912 287704 203924
rect 281500 203884 287704 203912
rect 281500 203872 281506 203884
rect 287698 203872 287704 203884
rect 287756 203912 287762 203924
rect 291286 203912 291292 203924
rect 287756 203884 291292 203912
rect 287756 203872 287762 203884
rect 291286 203872 291292 203884
rect 291344 203872 291350 203924
rect 302050 203872 302056 203924
rect 302108 203912 302114 203924
rect 313550 203912 313556 203924
rect 302108 203884 313556 203912
rect 302108 203872 302114 203884
rect 313550 203872 313556 203884
rect 313608 203872 313614 203924
rect 286778 203736 286784 203788
rect 286836 203776 286842 203788
rect 293218 203776 293224 203788
rect 286836 203748 293224 203776
rect 286836 203736 286842 203748
rect 293218 203736 293224 203748
rect 293276 203736 293282 203788
rect 266262 203668 266268 203720
rect 266320 203708 266326 203720
rect 291378 203708 291384 203720
rect 266320 203680 291384 203708
rect 266320 203668 266326 203680
rect 291378 203668 291384 203680
rect 291436 203668 291442 203720
rect 261570 203600 261576 203652
rect 261628 203640 261634 203652
rect 291194 203640 291200 203652
rect 261628 203612 291200 203640
rect 261628 203600 261634 203612
rect 291194 203600 291200 203612
rect 291252 203600 291258 203652
rect 556430 203600 556436 203652
rect 556488 203640 556494 203652
rect 568758 203640 568764 203652
rect 556488 203612 568764 203640
rect 556488 203600 556494 203612
rect 568758 203600 568764 203612
rect 568816 203600 568822 203652
rect 20346 203532 20352 203584
rect 20404 203572 20410 203584
rect 58526 203572 58532 203584
rect 20404 203544 58532 203572
rect 20404 203532 20410 203544
rect 58526 203532 58532 203544
rect 58584 203532 58590 203584
rect 149606 203532 149612 203584
rect 149664 203572 149670 203584
rect 289814 203572 289820 203584
rect 149664 203544 289820 203572
rect 149664 203532 149670 203544
rect 289814 203532 289820 203544
rect 289872 203532 289878 203584
rect 551370 203532 551376 203584
rect 551428 203572 551434 203584
rect 570046 203572 570052 203584
rect 551428 203544 570052 203572
rect 551428 203532 551434 203544
rect 570046 203532 570052 203544
rect 570104 203532 570110 203584
rect 96614 203464 96620 203516
rect 96672 203504 96678 203516
rect 99006 203504 99012 203516
rect 96672 203476 99012 203504
rect 96672 203464 96678 203476
rect 99006 203464 99012 203476
rect 99064 203464 99070 203516
rect 566550 203396 566556 203448
rect 566608 203436 566614 203448
rect 568850 203436 568856 203448
rect 566608 203408 568856 203436
rect 566608 203396 566614 203408
rect 568850 203396 568856 203408
rect 568908 203396 568914 203448
rect 465350 203192 465356 203244
rect 465408 203232 465414 203244
rect 467742 203232 467748 203244
rect 465408 203204 467748 203232
rect 465408 203192 465414 203204
rect 467742 203192 467748 203204
rect 467800 203192 467806 203244
rect 170490 203056 170496 203108
rect 170548 203096 170554 203108
rect 171134 203096 171140 203108
rect 170548 203068 171140 203096
rect 170548 203056 170554 203068
rect 171134 203056 171140 203068
rect 171192 203056 171198 203108
rect 500770 203056 500776 203108
rect 500828 203096 500834 203108
rect 503622 203096 503628 203108
rect 500828 203068 503628 203096
rect 500828 203056 500834 203068
rect 503622 203056 503628 203068
rect 503680 203056 503686 203108
rect 103514 202852 103520 202904
rect 103572 202852 103578 202904
rect 165430 202852 165436 202904
rect 165488 202892 165494 202904
rect 166258 202892 166264 202904
rect 165488 202864 166264 202892
rect 165488 202852 165494 202864
rect 166258 202852 166264 202864
rect 166316 202852 166322 202904
rect 413554 202852 413560 202904
rect 413612 202892 413618 202904
rect 414750 202892 414756 202904
rect 413612 202864 414756 202892
rect 413612 202852 413618 202864
rect 414750 202852 414756 202864
rect 414808 202852 414814 202904
rect 440050 202852 440056 202904
rect 440108 202892 440114 202904
rect 440878 202892 440884 202904
rect 440108 202864 440884 202892
rect 440108 202852 440114 202864
rect 440878 202852 440884 202864
rect 440936 202852 440942 202904
rect 445110 202852 445116 202904
rect 445168 202892 445174 202904
rect 446398 202892 446404 202904
rect 445168 202864 446404 202892
rect 445168 202852 445174 202864
rect 446398 202852 446404 202864
rect 446456 202852 446462 202904
rect 495710 202852 495716 202904
rect 495768 202892 495774 202904
rect 498562 202892 498568 202904
rect 495768 202864 498568 202892
rect 495768 202852 495774 202864
rect 498562 202852 498568 202864
rect 498620 202852 498626 202904
rect 21910 202784 21916 202836
rect 21968 202824 21974 202836
rect 23106 202824 23112 202836
rect 21968 202796 23112 202824
rect 21968 202784 21974 202796
rect 23106 202784 23112 202796
rect 23164 202784 23170 202836
rect 23382 202784 23388 202836
rect 23440 202824 23446 202836
rect 63586 202824 63592 202836
rect 23440 202796 63592 202824
rect 23440 202784 23446 202796
rect 63586 202784 63592 202796
rect 63644 202784 63650 202836
rect 103532 202824 103560 202852
rect 104066 202824 104072 202836
rect 103532 202796 104072 202824
rect 104066 202784 104072 202796
rect 104124 202784 104130 202836
rect 166276 202824 166304 202852
rect 296714 202824 296720 202836
rect 166276 202796 296720 202824
rect 296714 202784 296720 202796
rect 296772 202784 296778 202836
rect 303614 202784 303620 202836
rect 303672 202824 303678 202836
rect 419534 202824 419540 202836
rect 303672 202796 419540 202824
rect 303672 202784 303678 202796
rect 419534 202784 419540 202796
rect 419592 202784 419598 202836
rect 22922 202716 22928 202768
rect 22980 202756 22986 202768
rect 53466 202756 53472 202768
rect 22980 202728 53472 202756
rect 22980 202716 22986 202728
rect 53466 202716 53472 202728
rect 53524 202716 53530 202768
rect 175274 202716 175280 202768
rect 175332 202756 175338 202768
rect 285766 202756 285772 202768
rect 175332 202728 285772 202756
rect 175332 202716 175338 202728
rect 285766 202716 285772 202728
rect 285824 202716 285830 202768
rect 303798 202716 303804 202768
rect 303856 202756 303862 202768
rect 408494 202756 408500 202768
rect 303856 202728 408500 202756
rect 303856 202716 303862 202728
rect 408494 202716 408500 202728
rect 408552 202756 408558 202768
rect 409690 202756 409696 202768
rect 408552 202728 409696 202756
rect 408552 202716 408558 202728
rect 409690 202716 409696 202728
rect 409748 202716 409754 202768
rect 21818 202648 21824 202700
rect 21876 202688 21882 202700
rect 48406 202688 48412 202700
rect 21876 202660 48412 202688
rect 21876 202648 21882 202660
rect 48406 202648 48412 202660
rect 48464 202648 48470 202700
rect 195790 202648 195796 202700
rect 195848 202688 195854 202700
rect 284938 202688 284944 202700
rect 195848 202660 284944 202688
rect 195848 202648 195854 202660
rect 284938 202648 284944 202660
rect 284996 202648 285002 202700
rect 21726 202580 21732 202632
rect 21784 202620 21790 202632
rect 23382 202620 23388 202632
rect 21784 202592 23388 202620
rect 21784 202580 21790 202592
rect 23382 202580 23388 202592
rect 23440 202580 23446 202632
rect 226150 202580 226156 202632
rect 226208 202620 226214 202632
rect 287514 202620 287520 202632
rect 226208 202592 287520 202620
rect 226208 202580 226214 202592
rect 287514 202580 287520 202592
rect 287572 202580 287578 202632
rect 23106 202172 23112 202224
rect 23164 202212 23170 202224
rect 33318 202212 33324 202224
rect 23164 202184 33324 202212
rect 23164 202172 23170 202184
rect 33318 202172 33324 202184
rect 33376 202172 33382 202224
rect 455230 202172 455236 202224
rect 455288 202212 455294 202224
rect 564342 202212 564348 202224
rect 455288 202184 564348 202212
rect 455288 202172 455294 202184
rect 564342 202172 564348 202184
rect 564400 202172 564406 202224
rect 405918 202104 405924 202156
rect 405976 202144 405982 202156
rect 560938 202144 560944 202156
rect 405976 202116 560944 202144
rect 405976 202104 405982 202116
rect 560938 202104 560944 202116
rect 560996 202104 561002 202156
rect 185302 201424 185308 201476
rect 185360 201464 185366 201476
rect 292758 201464 292764 201476
rect 185360 201436 292764 201464
rect 185360 201424 185366 201436
rect 292758 201424 292764 201436
rect 292816 201424 292822 201476
rect 300670 201424 300676 201476
rect 300728 201464 300734 201476
rect 413278 201464 413284 201476
rect 300728 201436 413284 201464
rect 300728 201424 300734 201436
rect 413278 201424 413284 201436
rect 413336 201464 413342 201476
rect 413554 201464 413560 201476
rect 413336 201436 413560 201464
rect 413336 201424 413342 201436
rect 413554 201424 413560 201436
rect 413612 201424 413618 201476
rect 467742 201424 467748 201476
rect 467800 201464 467806 201476
rect 570322 201464 570328 201476
rect 467800 201436 570328 201464
rect 467800 201424 467806 201436
rect 570322 201424 570328 201436
rect 570380 201424 570386 201476
rect 572714 201424 572720 201476
rect 572772 201464 572778 201476
rect 573358 201464 573364 201476
rect 572772 201436 573364 201464
rect 572772 201424 572778 201436
rect 573358 201424 573364 201436
rect 573416 201424 573422 201476
rect 574370 201424 574376 201476
rect 574428 201464 574434 201476
rect 575474 201464 575480 201476
rect 574428 201436 575480 201464
rect 574428 201424 574434 201436
rect 575474 201424 575480 201436
rect 575532 201424 575538 201476
rect 216030 201356 216036 201408
rect 216088 201396 216094 201408
rect 288526 201396 288532 201408
rect 216088 201368 288532 201396
rect 216088 201356 216094 201368
rect 288526 201356 288532 201368
rect 288584 201356 288590 201408
rect 296438 201356 296444 201408
rect 296496 201396 296502 201408
rect 299198 201396 299204 201408
rect 296496 201368 299204 201396
rect 296496 201356 296502 201368
rect 299198 201356 299204 201368
rect 299256 201396 299262 201408
rect 338850 201396 338856 201408
rect 299256 201368 338856 201396
rect 299256 201356 299262 201368
rect 338850 201356 338856 201368
rect 338908 201356 338914 201408
rect 471330 201356 471336 201408
rect 471388 201396 471394 201408
rect 572732 201396 572760 201424
rect 471388 201368 572760 201396
rect 471388 201356 471394 201368
rect 231210 201288 231216 201340
rect 231268 201328 231274 201340
rect 231268 201300 277394 201328
rect 231268 201288 231274 201300
rect 277366 201260 277394 201300
rect 476114 201288 476120 201340
rect 476172 201328 476178 201340
rect 575750 201328 575756 201340
rect 476172 201300 575756 201328
rect 476172 201288 476178 201300
rect 575750 201288 575756 201300
rect 575808 201288 575814 201340
rect 291562 201260 291568 201272
rect 277366 201232 291568 201260
rect 291562 201220 291568 201232
rect 291620 201260 291626 201272
rect 292666 201260 292672 201272
rect 291620 201232 292672 201260
rect 291620 201220 291626 201232
rect 292666 201220 292672 201232
rect 292724 201220 292730 201272
rect 498562 201220 498568 201272
rect 498620 201260 498626 201272
rect 574094 201260 574100 201272
rect 498620 201232 574100 201260
rect 498620 201220 498626 201232
rect 574094 201220 574100 201232
rect 574152 201220 574158 201272
rect 503622 201152 503628 201204
rect 503680 201192 503686 201204
rect 574462 201192 574468 201204
rect 503680 201164 574468 201192
rect 503680 201152 503686 201164
rect 574462 201152 574468 201164
rect 574520 201152 574526 201204
rect 574462 201016 574468 201068
rect 574520 201056 574526 201068
rect 575934 201056 575940 201068
rect 574520 201028 575940 201056
rect 574520 201016 574526 201028
rect 575934 201016 575940 201028
rect 575992 201016 575998 201068
rect 299198 200812 299204 200864
rect 299256 200852 299262 200864
rect 374270 200852 374276 200864
rect 299256 200824 374276 200852
rect 299256 200812 299262 200824
rect 374270 200812 374276 200824
rect 374328 200812 374334 200864
rect 24118 200744 24124 200796
rect 24176 200784 24182 200796
rect 185302 200784 185308 200796
rect 24176 200756 185308 200784
rect 24176 200744 24182 200756
rect 185302 200744 185308 200756
rect 185360 200744 185366 200796
rect 210970 200744 210976 200796
rect 211028 200784 211034 200796
rect 285674 200784 285680 200796
rect 211028 200756 285680 200784
rect 211028 200744 211034 200756
rect 285674 200744 285680 200756
rect 285732 200744 285738 200796
rect 296622 200744 296628 200796
rect 296680 200784 296686 200796
rect 302234 200784 302240 200796
rect 296680 200756 302240 200784
rect 296680 200744 296686 200756
rect 302234 200744 302240 200756
rect 302292 200784 302298 200796
rect 382274 200784 382280 200796
rect 302292 200756 382280 200784
rect 302292 200744 302298 200756
rect 382274 200744 382280 200756
rect 382332 200744 382338 200796
rect 460290 200744 460296 200796
rect 460348 200784 460354 200796
rect 574370 200784 574376 200796
rect 460348 200756 574376 200784
rect 460348 200744 460354 200756
rect 574370 200744 574376 200756
rect 574428 200744 574434 200796
rect 285674 200132 285680 200184
rect 285732 200172 285738 200184
rect 286870 200172 286876 200184
rect 285732 200144 286876 200172
rect 285732 200132 285738 200144
rect 286870 200132 286876 200144
rect 286928 200172 286934 200184
rect 287606 200172 287612 200184
rect 286928 200144 287612 200172
rect 286928 200132 286934 200144
rect 287606 200132 287612 200144
rect 287664 200132 287670 200184
rect 23566 200064 23572 200116
rect 23624 200104 23630 200116
rect 158714 200104 158720 200116
rect 23624 200076 158720 200104
rect 23624 200064 23630 200076
rect 158714 200064 158720 200076
rect 158772 200064 158778 200116
rect 15010 199996 15016 200048
rect 15068 200036 15074 200048
rect 139394 200036 139400 200048
rect 15068 200008 139400 200036
rect 15068 199996 15074 200008
rect 139394 199996 139400 200008
rect 139452 199996 139458 200048
rect 15102 199928 15108 199980
rect 15160 199968 15166 199980
rect 17126 199968 17132 199980
rect 15160 199940 17132 199968
rect 15160 199928 15166 199940
rect 17126 199928 17132 199940
rect 17184 199968 17190 199980
rect 128354 199968 128360 199980
rect 17184 199940 128360 199968
rect 17184 199928 17190 199940
rect 128354 199928 128360 199940
rect 128412 199928 128418 199980
rect 17770 199860 17776 199912
rect 17828 199900 17834 199912
rect 103422 199900 103428 199912
rect 17828 199872 103428 199900
rect 17828 199860 17834 199872
rect 103422 199860 103428 199872
rect 103480 199860 103486 199912
rect 14918 199452 14924 199504
rect 14976 199492 14982 199504
rect 23566 199492 23572 199504
rect 14976 199464 23572 199492
rect 14976 199452 14982 199464
rect 23566 199452 23572 199464
rect 23624 199452 23630 199504
rect 22002 199384 22008 199436
rect 22060 199424 22066 199436
rect 109034 199424 109040 199436
rect 22060 199396 109040 199424
rect 22060 199384 22066 199396
rect 109034 199384 109040 199396
rect 109092 199384 109098 199436
rect 20530 199044 20536 199096
rect 20588 199084 20594 199096
rect 22002 199084 22008 199096
rect 20588 199056 22008 199084
rect 20588 199044 20594 199056
rect 22002 199044 22008 199056
rect 22060 199044 22066 199096
rect 17586 198704 17592 198756
rect 17644 198744 17650 198756
rect 17770 198744 17776 198756
rect 17644 198716 17776 198744
rect 17644 198704 17650 198716
rect 17770 198704 17776 198716
rect 17828 198704 17834 198756
rect 440878 198636 440884 198688
rect 440936 198676 440942 198688
rect 571610 198676 571616 198688
rect 440936 198648 571616 198676
rect 440936 198636 440942 198648
rect 571610 198636 571616 198648
rect 571668 198636 571674 198688
rect 446398 198568 446404 198620
rect 446456 198608 446462 198620
rect 575658 198608 575664 198620
rect 446456 198580 575664 198608
rect 446456 198568 446462 198580
rect 575658 198568 575664 198580
rect 575716 198568 575722 198620
rect 20530 197956 20536 198008
rect 20588 197996 20594 198008
rect 166258 197996 166264 198008
rect 20588 197968 166264 197996
rect 20588 197956 20594 197968
rect 166258 197956 166264 197968
rect 166316 197956 166322 198008
rect 408494 197956 408500 198008
rect 408552 197996 408558 198008
rect 574186 197996 574192 198008
rect 408552 197968 574192 197996
rect 408552 197956 408558 197968
rect 574186 197956 574192 197968
rect 574244 197956 574250 198008
rect 287514 189728 287520 189780
rect 287572 189768 287578 189780
rect 424318 189768 424324 189780
rect 287572 189740 424324 189768
rect 287572 189728 287578 189740
rect 424318 189728 424324 189740
rect 424376 189728 424382 189780
rect 23658 188980 23664 189032
rect 23716 189020 23722 189032
rect 171134 189020 171140 189032
rect 23716 188992 171140 189020
rect 23716 188980 23722 188992
rect 171134 188980 171140 188992
rect 171192 188980 171198 189032
rect 434714 188980 434720 189032
rect 434772 189020 434778 189032
rect 565722 189020 565728 189032
rect 434772 188992 565728 189020
rect 434772 188980 434778 188992
rect 565722 188980 565728 188992
rect 565780 188980 565786 189032
rect 16390 188912 16396 188964
rect 16448 188952 16454 188964
rect 113174 188952 113180 188964
rect 16448 188924 113180 188952
rect 16448 188912 16454 188924
rect 113174 188912 113180 188924
rect 113232 188912 113238 188964
rect 489914 188912 489920 188964
rect 489972 188952 489978 188964
rect 575566 188952 575572 188964
rect 489972 188924 575572 188952
rect 489972 188912 489978 188924
rect 575566 188912 575572 188924
rect 575624 188912 575630 188964
rect 565722 188368 565728 188420
rect 565780 188408 565786 188420
rect 572990 188408 572996 188420
rect 565780 188380 572996 188408
rect 565780 188368 565786 188380
rect 572990 188368 572996 188380
rect 573048 188368 573054 188420
rect 296530 188300 296536 188352
rect 296588 188340 296594 188352
rect 300670 188340 300676 188352
rect 296588 188312 300676 188340
rect 296588 188300 296594 188312
rect 300670 188300 300676 188312
rect 300728 188340 300734 188352
rect 368474 188340 368480 188352
rect 300728 188312 368480 188340
rect 300728 188300 300734 188312
rect 368474 188300 368480 188312
rect 368532 188300 368538 188352
rect 560938 188300 560944 188352
rect 560996 188340 561002 188352
rect 578326 188340 578332 188352
rect 560996 188312 578332 188340
rect 560996 188300 561002 188312
rect 578326 188300 578332 188312
rect 578384 188300 578390 188352
rect 2774 187688 2780 187740
rect 2832 187728 2838 187740
rect 4798 187728 4804 187740
rect 2832 187700 4804 187728
rect 2832 187688 2838 187700
rect 4798 187688 4804 187700
rect 4856 187688 4862 187740
rect 18966 187688 18972 187740
rect 19024 187728 19030 187740
rect 23658 187728 23664 187740
rect 19024 187700 23664 187728
rect 19024 187688 19030 187700
rect 23658 187688 23664 187700
rect 23716 187688 23722 187740
rect 575566 187688 575572 187740
rect 575624 187728 575630 187740
rect 575750 187728 575756 187740
rect 575624 187700 575756 187728
rect 575624 187688 575630 187700
rect 575750 187688 575756 187700
rect 575808 187688 575814 187740
rect 305730 187620 305736 187672
rect 305788 187660 305794 187672
rect 398834 187660 398840 187672
rect 305788 187632 398840 187660
rect 305788 187620 305794 187632
rect 398834 187620 398840 187632
rect 398892 187620 398898 187672
rect 297818 187552 297824 187604
rect 297876 187592 297882 187604
rect 305086 187592 305092 187604
rect 297876 187564 305092 187592
rect 297876 187552 297882 187564
rect 305086 187552 305092 187564
rect 305144 187592 305150 187604
rect 393314 187592 393320 187604
rect 305144 187564 393320 187592
rect 305144 187552 305150 187564
rect 393314 187552 393320 187564
rect 393372 187552 393378 187604
rect 303246 187484 303252 187536
rect 303304 187524 303310 187536
rect 362954 187524 362960 187536
rect 303304 187496 362960 187524
rect 303304 187484 303310 187496
rect 362954 187484 362960 187496
rect 363012 187484 363018 187536
rect 296530 187144 296536 187196
rect 296588 187184 296594 187196
rect 302234 187184 302240 187196
rect 296588 187156 302240 187184
rect 296588 187144 296594 187156
rect 302234 187144 302240 187156
rect 302292 187144 302298 187196
rect 285490 187008 285496 187060
rect 285548 187048 285554 187060
rect 294138 187048 294144 187060
rect 285548 187020 294144 187048
rect 285548 187008 285554 187020
rect 294138 187008 294144 187020
rect 294196 187008 294202 187060
rect 276014 186940 276020 186992
rect 276072 186980 276078 186992
rect 298738 186980 298744 186992
rect 276072 186952 298744 186980
rect 276072 186940 276078 186952
rect 298738 186940 298744 186952
rect 298796 186940 298802 186992
rect 299106 186940 299112 186992
rect 299164 186980 299170 186992
rect 303338 186980 303344 186992
rect 299164 186952 303344 186980
rect 299164 186940 299170 186952
rect 303338 186940 303344 186952
rect 303396 186980 303402 186992
rect 347774 186980 347780 186992
rect 303396 186952 347780 186980
rect 303396 186940 303402 186952
rect 347774 186940 347780 186952
rect 347832 186940 347838 186992
rect 413278 186940 413284 186992
rect 413336 186980 413342 186992
rect 579614 186980 579620 186992
rect 413336 186952 579620 186980
rect 413336 186940 413342 186952
rect 579614 186940 579620 186952
rect 579672 186940 579678 186992
rect 297910 186396 297916 186448
rect 297968 186436 297974 186448
rect 303706 186436 303712 186448
rect 297968 186408 303712 186436
rect 297968 186396 297974 186408
rect 303706 186396 303712 186408
rect 303764 186396 303770 186448
rect 303062 186328 303068 186380
rect 303120 186368 303126 186380
rect 303246 186368 303252 186380
rect 303120 186340 303252 186368
rect 303120 186328 303126 186340
rect 303246 186328 303252 186340
rect 303304 186328 303310 186380
rect 192478 186260 192484 186312
rect 192536 186300 192542 186312
rect 285122 186300 285128 186312
rect 192536 186272 285128 186300
rect 192536 186260 192542 186272
rect 285122 186260 285128 186272
rect 285180 186300 285186 186312
rect 285582 186300 285588 186312
rect 285180 186272 285588 186300
rect 285180 186260 285186 186272
rect 285582 186260 285588 186272
rect 285640 186260 285646 186312
rect 17862 185920 17868 185972
rect 17920 185960 17926 185972
rect 17920 185932 26234 185960
rect 17920 185920 17926 185932
rect 23014 185852 23020 185904
rect 23072 185892 23078 185904
rect 24118 185892 24124 185904
rect 23072 185864 24124 185892
rect 23072 185852 23078 185864
rect 24118 185852 24124 185864
rect 24176 185852 24182 185904
rect 26206 185892 26234 185932
rect 286870 185920 286876 185972
rect 286928 185960 286934 185972
rect 292758 185960 292764 185972
rect 286928 185932 292764 185960
rect 286928 185920 286934 185932
rect 292758 185920 292764 185932
rect 292816 185920 292822 185972
rect 173894 185892 173900 185904
rect 26206 185864 173900 185892
rect 173894 185852 173900 185864
rect 173952 185852 173958 185904
rect 200114 185852 200120 185904
rect 200172 185892 200178 185904
rect 290090 185892 290096 185904
rect 200172 185864 290096 185892
rect 200172 185852 200178 185864
rect 290090 185852 290096 185864
rect 290148 185852 290154 185904
rect 300578 185852 300584 185904
rect 300636 185892 300642 185904
rect 304994 185892 305000 185904
rect 300636 185864 305000 185892
rect 300636 185852 300642 185864
rect 304994 185852 305000 185864
rect 305052 185852 305058 185904
rect 419534 185852 419540 185904
rect 419592 185892 419598 185904
rect 570230 185892 570236 185904
rect 419592 185864 570236 185892
rect 419592 185852 419598 185864
rect 570230 185852 570236 185864
rect 570288 185852 570294 185904
rect 2958 149064 2964 149116
rect 3016 149104 3022 149116
rect 6362 149104 6368 149116
rect 3016 149076 6368 149104
rect 3016 149064 3022 149076
rect 6362 149064 6368 149076
rect 6420 149064 6426 149116
rect 2774 136688 2780 136740
rect 2832 136728 2838 136740
rect 4982 136728 4988 136740
rect 2832 136700 4988 136728
rect 2832 136688 2838 136700
rect 4982 136688 4988 136700
rect 5040 136688 5046 136740
rect 3418 110440 3424 110492
rect 3476 110480 3482 110492
rect 9030 110480 9036 110492
rect 3476 110452 9036 110480
rect 3476 110440 3482 110452
rect 9030 110440 9036 110452
rect 9088 110440 9094 110492
rect 2774 84328 2780 84380
rect 2832 84368 2838 84380
rect 5074 84368 5080 84380
rect 2832 84340 5080 84368
rect 2832 84328 2838 84340
rect 5074 84328 5080 84340
rect 5132 84328 5138 84380
rect 574186 79296 574192 79348
rect 574244 79336 574250 79348
rect 574462 79336 574468 79348
rect 574244 79308 574468 79336
rect 574244 79296 574250 79308
rect 574462 79296 574468 79308
rect 574520 79296 574526 79348
rect 288526 78044 288532 78056
rect 240796 78016 288532 78044
rect 16390 77936 16396 77988
rect 16448 77976 16454 77988
rect 16448 77948 103514 77976
rect 16448 77936 16454 77948
rect 23014 77868 23020 77920
rect 23072 77908 23078 77920
rect 25498 77908 25504 77920
rect 23072 77880 25504 77908
rect 23072 77868 23078 77880
rect 25498 77868 25504 77880
rect 25556 77868 25562 77920
rect 103486 77908 103514 77948
rect 193232 77948 219434 77976
rect 193232 77920 193260 77948
rect 114186 77908 114192 77920
rect 103486 77880 114192 77908
rect 114186 77868 114192 77880
rect 114244 77868 114250 77920
rect 193214 77868 193220 77920
rect 193272 77868 193278 77920
rect 219406 77840 219434 77948
rect 240796 77920 240824 78016
rect 288526 78004 288532 78016
rect 288584 78004 288590 78056
rect 300578 78004 300584 78056
rect 300636 78044 300642 78056
rect 300636 78016 332640 78044
rect 300636 78004 300642 78016
rect 290090 77976 290096 77988
rect 248386 77948 290096 77976
rect 240778 77868 240784 77920
rect 240836 77868 240842 77920
rect 248386 77840 248414 77948
rect 290090 77936 290096 77948
rect 290148 77936 290154 77988
rect 297818 77936 297824 77988
rect 297876 77976 297882 77988
rect 297876 77948 316034 77976
rect 297876 77936 297882 77948
rect 284938 77868 284944 77920
rect 284996 77908 285002 77920
rect 294138 77908 294144 77920
rect 284996 77880 294144 77908
rect 284996 77868 285002 77880
rect 294138 77868 294144 77880
rect 294196 77868 294202 77920
rect 219406 77812 248414 77840
rect 316006 77840 316034 77948
rect 332612 77920 332640 78016
rect 332594 77868 332600 77920
rect 332652 77868 332658 77920
rect 335998 77840 336004 77852
rect 316006 77812 336004 77840
rect 335998 77800 336004 77812
rect 336056 77800 336062 77852
rect 20530 77052 20536 77104
rect 20588 77092 20594 77104
rect 23474 77092 23480 77104
rect 20588 77064 23480 77092
rect 20588 77052 20594 77064
rect 23474 77052 23480 77064
rect 23532 77052 23538 77104
rect 299198 76712 299204 76764
rect 299256 76752 299262 76764
rect 329098 76752 329104 76764
rect 299256 76724 329104 76752
rect 299256 76712 299262 76724
rect 329098 76712 329104 76724
rect 329156 76712 329162 76764
rect 293218 76644 293224 76696
rect 293276 76684 293282 76696
rect 418154 76684 418160 76696
rect 293276 76656 418160 76684
rect 293276 76644 293282 76656
rect 418154 76644 418160 76656
rect 418212 76644 418218 76696
rect 430574 76644 430580 76696
rect 430632 76684 430638 76696
rect 568850 76684 568856 76696
rect 430632 76656 568856 76684
rect 430632 76644 430638 76656
rect 568850 76644 568856 76656
rect 568908 76644 568914 76696
rect 222194 76576 222200 76628
rect 222252 76616 222258 76628
rect 300118 76616 300124 76628
rect 222252 76588 300124 76616
rect 222252 76576 222258 76588
rect 300118 76576 300124 76588
rect 300176 76576 300182 76628
rect 301498 76576 301504 76628
rect 301556 76616 301562 76628
rect 376754 76616 376760 76628
rect 301556 76588 376760 76616
rect 301556 76576 301562 76588
rect 376754 76576 376760 76588
rect 376812 76576 376818 76628
rect 404354 76576 404360 76628
rect 404412 76616 404418 76628
rect 571426 76616 571432 76628
rect 404412 76588 571432 76616
rect 404412 76576 404418 76588
rect 571426 76576 571432 76588
rect 571484 76576 571490 76628
rect 153010 76508 153016 76560
rect 153068 76548 153074 76560
rect 580258 76548 580264 76560
rect 153068 76520 580264 76548
rect 153068 76508 153074 76520
rect 580258 76508 580264 76520
rect 580316 76508 580322 76560
rect 13078 76100 13084 76152
rect 13136 76140 13142 76152
rect 28166 76140 28172 76152
rect 13136 76112 28172 76140
rect 13136 76100 13142 76112
rect 28166 76100 28172 76112
rect 28224 76100 28230 76152
rect 17678 76032 17684 76084
rect 17736 76072 17742 76084
rect 119890 76072 119896 76084
rect 17736 76044 119896 76072
rect 17736 76032 17742 76044
rect 119890 76032 119896 76044
rect 119948 76032 119954 76084
rect 219434 76032 219440 76084
rect 219492 76072 219498 76084
rect 297174 76072 297180 76084
rect 219492 76044 297180 76072
rect 219492 76032 219498 76044
rect 297174 76032 297180 76044
rect 297232 76032 297238 76084
rect 18966 75964 18972 76016
rect 19024 76004 19030 76016
rect 169754 76004 169760 76016
rect 19024 75976 169760 76004
rect 19024 75964 19030 75976
rect 169754 75964 169760 75976
rect 169812 75964 169818 76016
rect 200298 75964 200304 76016
rect 200356 76004 200362 76016
rect 291470 76004 291476 76016
rect 200356 75976 291476 76004
rect 200356 75964 200362 75976
rect 291470 75964 291476 75976
rect 291528 75964 291534 76016
rect 385034 75964 385040 76016
rect 385092 76004 385098 76016
rect 571426 76004 571432 76016
rect 385092 75976 571432 76004
rect 385092 75964 385098 75976
rect 571426 75964 571432 75976
rect 571484 75964 571490 76016
rect 18782 75896 18788 75948
rect 18840 75936 18846 75948
rect 134426 75936 134432 75948
rect 18840 75908 134432 75936
rect 18840 75896 18846 75908
rect 134426 75896 134432 75908
rect 134484 75896 134490 75948
rect 153102 75896 153108 75948
rect 153160 75936 153166 75948
rect 574186 75936 574192 75948
rect 153160 75908 574192 75936
rect 153160 75896 153166 75908
rect 574186 75896 574192 75908
rect 574244 75896 574250 75948
rect 19150 75828 19156 75880
rect 19208 75868 19214 75880
rect 88978 75868 88984 75880
rect 19208 75840 88984 75868
rect 19208 75828 19214 75840
rect 88978 75828 88984 75840
rect 89036 75828 89042 75880
rect 144822 75828 144828 75880
rect 144880 75868 144886 75880
rect 149606 75868 149612 75880
rect 144880 75840 149612 75868
rect 144880 75828 144886 75840
rect 149606 75828 149612 75840
rect 149664 75868 149670 75880
rect 149974 75868 149980 75880
rect 149664 75840 149980 75868
rect 149664 75828 149670 75840
rect 149974 75828 149980 75840
rect 150032 75828 150038 75880
rect 188338 75828 188344 75880
rect 188396 75868 188402 75880
rect 190362 75868 190368 75880
rect 188396 75840 190368 75868
rect 188396 75828 188402 75840
rect 190362 75828 190368 75840
rect 190420 75868 190426 75880
rect 284294 75868 284300 75880
rect 190420 75840 284300 75868
rect 190420 75828 190426 75840
rect 284294 75828 284300 75840
rect 284352 75828 284358 75880
rect 301682 75828 301688 75880
rect 301740 75868 301746 75880
rect 301958 75868 301964 75880
rect 301740 75840 301964 75868
rect 301740 75828 301746 75840
rect 301958 75828 301964 75840
rect 302016 75868 302022 75880
rect 318610 75868 318616 75880
rect 302016 75840 318616 75868
rect 302016 75828 302022 75840
rect 318610 75828 318616 75840
rect 318668 75828 318674 75880
rect 332594 75828 332600 75880
rect 332652 75868 332658 75880
rect 389450 75868 389456 75880
rect 332652 75840 389456 75868
rect 332652 75828 332658 75840
rect 389450 75828 389456 75840
rect 389508 75828 389514 75880
rect 423674 75828 423680 75880
rect 423732 75868 423738 75880
rect 424870 75868 424876 75880
rect 423732 75840 424876 75868
rect 423732 75828 423738 75840
rect 424870 75828 424876 75840
rect 424928 75868 424934 75880
rect 429930 75868 429936 75880
rect 424928 75840 429936 75868
rect 424928 75828 424934 75840
rect 429930 75828 429936 75840
rect 429988 75828 429994 75880
rect 505830 75828 505836 75880
rect 505888 75868 505894 75880
rect 567746 75868 567752 75880
rect 505888 75840 567752 75868
rect 505888 75828 505894 75840
rect 567746 75828 567752 75840
rect 567804 75828 567810 75880
rect 20438 75760 20444 75812
rect 20496 75800 20502 75812
rect 73798 75800 73804 75812
rect 20496 75772 73804 75800
rect 20496 75760 20502 75772
rect 73798 75760 73804 75772
rect 73856 75760 73862 75812
rect 216030 75760 216036 75812
rect 216088 75800 216094 75812
rect 217318 75800 217324 75812
rect 216088 75772 217324 75800
rect 216088 75760 216094 75772
rect 217318 75760 217324 75772
rect 217376 75760 217382 75812
rect 261570 75760 261576 75812
rect 261628 75800 261634 75812
rect 264882 75800 264888 75812
rect 261628 75772 264888 75800
rect 261628 75760 261634 75772
rect 264882 75760 264888 75772
rect 264940 75760 264946 75812
rect 511258 75760 511264 75812
rect 511316 75800 511322 75812
rect 571518 75800 571524 75812
rect 511316 75772 571524 75800
rect 511316 75760 511322 75772
rect 571518 75760 571524 75772
rect 571576 75760 571582 75812
rect 20346 75692 20352 75744
rect 20404 75732 20410 75744
rect 59262 75732 59268 75744
rect 20404 75704 59268 75732
rect 20404 75692 20410 75704
rect 59262 75692 59268 75704
rect 59320 75692 59326 75744
rect 515950 75692 515956 75744
rect 516008 75732 516014 75744
rect 574278 75732 574284 75744
rect 516008 75704 574284 75732
rect 516008 75692 516014 75704
rect 574278 75692 574284 75704
rect 574336 75692 574342 75744
rect 21818 75624 21824 75676
rect 21876 75664 21882 75676
rect 49050 75664 49056 75676
rect 21876 75636 49056 75664
rect 21876 75624 21882 75636
rect 49050 75624 49056 75636
rect 49108 75624 49114 75676
rect 520274 75624 520280 75676
rect 520332 75664 520338 75676
rect 521010 75664 521016 75676
rect 520332 75636 521016 75664
rect 520332 75624 520338 75636
rect 521010 75624 521016 75636
rect 521068 75664 521074 75676
rect 567654 75664 567660 75676
rect 521068 75636 567660 75664
rect 521068 75624 521074 75636
rect 567654 75624 567660 75636
rect 567712 75624 567718 75676
rect 6178 75556 6184 75608
rect 6236 75596 6242 75608
rect 23382 75596 23388 75608
rect 6236 75568 23388 75596
rect 6236 75556 6242 75568
rect 23382 75556 23388 75568
rect 23440 75556 23446 75608
rect 526070 75556 526076 75608
rect 526128 75596 526134 75608
rect 572898 75596 572904 75608
rect 526128 75568 572904 75596
rect 526128 75556 526134 75568
rect 572898 75556 572904 75568
rect 572956 75556 572962 75608
rect 266262 75488 266268 75540
rect 266320 75528 266326 75540
rect 270494 75528 270500 75540
rect 266320 75500 270500 75528
rect 266320 75488 266326 75500
rect 270494 75488 270500 75500
rect 270552 75488 270558 75540
rect 529934 75488 529940 75540
rect 529992 75528 529998 75540
rect 531130 75528 531136 75540
rect 529992 75500 531136 75528
rect 529992 75488 529998 75500
rect 531130 75488 531136 75500
rect 531188 75528 531194 75540
rect 572806 75528 572812 75540
rect 531188 75500 572812 75528
rect 531188 75488 531194 75500
rect 572806 75488 572812 75500
rect 572864 75488 572870 75540
rect 241330 75420 241336 75472
rect 241388 75460 241394 75472
rect 248414 75460 248420 75472
rect 241388 75432 248420 75460
rect 241388 75420 241394 75432
rect 248414 75420 248420 75432
rect 248472 75420 248478 75472
rect 251082 75420 251088 75472
rect 251140 75460 251146 75472
rect 261478 75460 261484 75472
rect 251140 75432 261484 75460
rect 251140 75420 251146 75432
rect 261478 75420 261484 75432
rect 261536 75420 261542 75472
rect 286778 75420 286784 75472
rect 286836 75460 286842 75472
rect 308398 75460 308404 75472
rect 286836 75432 308404 75460
rect 286836 75420 286842 75432
rect 308398 75420 308404 75432
rect 308456 75420 308462 75472
rect 246390 75352 246396 75404
rect 246448 75392 246454 75404
rect 263594 75392 263600 75404
rect 246448 75364 263600 75392
rect 246448 75352 246454 75364
rect 263594 75352 263600 75364
rect 263652 75392 263658 75404
rect 292850 75392 292856 75404
rect 263652 75364 292856 75392
rect 263652 75352 263658 75364
rect 292850 75352 292856 75364
rect 292908 75352 292914 75404
rect 235902 75284 235908 75336
rect 235960 75324 235966 75336
rect 240042 75324 240048 75336
rect 235960 75296 240048 75324
rect 235960 75284 235966 75296
rect 240042 75284 240048 75296
rect 240100 75324 240106 75336
rect 287882 75324 287888 75336
rect 240100 75296 287888 75324
rect 240100 75284 240106 75296
rect 287882 75284 287888 75296
rect 287940 75284 287946 75336
rect 319438 75284 319444 75336
rect 319496 75324 319502 75336
rect 333790 75324 333796 75336
rect 319496 75296 333796 75324
rect 319496 75284 319502 75296
rect 333790 75284 333796 75296
rect 333848 75284 333854 75336
rect 292666 75256 292672 75268
rect 238726 75228 292672 75256
rect 49050 75148 49056 75200
rect 49108 75188 49114 75200
rect 116578 75188 116584 75200
rect 49108 75160 116584 75188
rect 49108 75148 49114 75160
rect 116578 75148 116584 75160
rect 116636 75148 116642 75200
rect 191834 75148 191840 75200
rect 191892 75188 191898 75200
rect 200390 75188 200396 75200
rect 191892 75160 200396 75188
rect 191892 75148 191898 75160
rect 200390 75148 200396 75160
rect 200448 75148 200454 75200
rect 226150 75148 226156 75200
rect 226208 75188 226214 75200
rect 234430 75188 234436 75200
rect 226208 75160 234436 75188
rect 226208 75148 226214 75160
rect 234430 75148 234436 75160
rect 234488 75148 234494 75200
rect 231210 75080 231216 75132
rect 231268 75120 231274 75132
rect 235902 75120 235908 75132
rect 231268 75092 235908 75120
rect 231268 75080 231274 75092
rect 235902 75080 235908 75092
rect 235960 75120 235966 75132
rect 238726 75120 238754 75228
rect 292666 75216 292672 75228
rect 292724 75216 292730 75268
rect 292850 75216 292856 75268
rect 292908 75256 292914 75268
rect 301682 75256 301688 75268
rect 292908 75228 301688 75256
rect 292908 75216 292914 75228
rect 301682 75216 301688 75228
rect 301740 75216 301746 75268
rect 307938 75216 307944 75268
rect 307996 75256 308002 75268
rect 323670 75256 323676 75268
rect 307996 75228 323676 75256
rect 307996 75216 308002 75228
rect 323670 75216 323676 75228
rect 323728 75216 323734 75268
rect 239490 75148 239496 75200
rect 239548 75188 239554 75200
rect 515950 75188 515956 75200
rect 239548 75160 515956 75188
rect 239548 75148 239554 75160
rect 515950 75148 515956 75160
rect 516008 75148 516014 75200
rect 235960 75092 238754 75120
rect 235960 75080 235966 75092
rect 271690 74808 271696 74860
rect 271748 74848 271754 74860
rect 276106 74848 276112 74860
rect 271748 74820 276112 74848
rect 271748 74808 271754 74820
rect 276106 74808 276112 74820
rect 276164 74808 276170 74860
rect 270494 74536 270500 74588
rect 270552 74576 270558 74588
rect 271782 74576 271788 74588
rect 270552 74548 271788 74576
rect 270552 74536 270558 74548
rect 271782 74536 271788 74548
rect 271840 74536 271846 74588
rect 414014 74536 414020 74588
rect 414072 74576 414078 74588
rect 414750 74576 414756 74588
rect 414072 74548 414756 74576
rect 414072 74536 414078 74548
rect 414750 74536 414756 74548
rect 414808 74576 414814 74588
rect 507026 74576 507032 74588
rect 414808 74548 507032 74576
rect 414808 74536 414814 74548
rect 507026 74536 507032 74548
rect 507084 74536 507090 74588
rect 19242 74468 19248 74520
rect 19300 74508 19306 74520
rect 94314 74508 94320 74520
rect 19300 74480 94320 74508
rect 19300 74468 19306 74480
rect 94314 74468 94320 74480
rect 94372 74468 94378 74520
rect 256602 74468 256608 74520
rect 256660 74508 256666 74520
rect 289998 74508 290004 74520
rect 256660 74480 290004 74508
rect 256660 74468 256666 74480
rect 289998 74468 290004 74480
rect 290056 74468 290062 74520
rect 302050 74468 302056 74520
rect 302108 74508 302114 74520
rect 313274 74508 313280 74520
rect 302108 74480 313280 74508
rect 302108 74468 302114 74480
rect 313274 74468 313280 74480
rect 313332 74468 313338 74520
rect 536098 74468 536104 74520
rect 536156 74508 536162 74520
rect 568574 74508 568580 74520
rect 536156 74480 568580 74508
rect 536156 74468 536162 74480
rect 568574 74468 568580 74480
rect 568632 74468 568638 74520
rect 20622 74400 20628 74452
rect 20680 74440 20686 74452
rect 68278 74440 68284 74452
rect 20680 74412 68284 74440
rect 20680 74400 20686 74412
rect 68278 74400 68284 74412
rect 68336 74400 68342 74452
rect 271782 74400 271788 74452
rect 271840 74440 271846 74452
rect 291378 74440 291384 74452
rect 271840 74412 291384 74440
rect 271840 74400 271846 74412
rect 291378 74400 291384 74412
rect 291436 74400 291442 74452
rect 303154 74400 303160 74452
rect 303212 74440 303218 74452
rect 307846 74440 307852 74452
rect 303212 74412 307852 74440
rect 303212 74400 303218 74412
rect 307846 74400 307852 74412
rect 307904 74400 307910 74452
rect 541250 74400 541256 74452
rect 541308 74440 541314 74452
rect 567562 74440 567568 74452
rect 541308 74412 567568 74440
rect 541308 74400 541314 74412
rect 567562 74400 567568 74412
rect 567620 74400 567626 74452
rect 21726 74332 21732 74384
rect 21784 74372 21790 74384
rect 64138 74372 64144 74384
rect 21784 74344 64144 74372
rect 21784 74332 21790 74344
rect 64138 74332 64144 74344
rect 64196 74332 64202 74384
rect 281442 74332 281448 74384
rect 281500 74372 281506 74384
rect 291286 74372 291292 74384
rect 281500 74344 291292 74372
rect 281500 74332 281506 74344
rect 291286 74332 291292 74344
rect 291344 74332 291350 74384
rect 545758 74332 545764 74384
rect 545816 74372 545822 74384
rect 568666 74372 568672 74384
rect 545816 74344 568672 74372
rect 545816 74332 545822 74344
rect 568666 74332 568672 74344
rect 568724 74332 568730 74384
rect 23198 74264 23204 74316
rect 23256 74304 23262 74316
rect 43438 74304 43444 74316
rect 23256 74276 43444 74304
rect 23256 74264 23262 74276
rect 43438 74264 43444 74276
rect 43496 74264 43502 74316
rect 560938 74264 560944 74316
rect 560996 74304 561002 74316
rect 570138 74304 570144 74316
rect 560996 74276 570144 74304
rect 560996 74264 561002 74276
rect 570138 74264 570144 74276
rect 570196 74264 570202 74316
rect 23106 74196 23112 74248
rect 23164 74236 23170 74248
rect 37918 74236 37924 74248
rect 23164 74208 37924 74236
rect 23164 74196 23170 74208
rect 37918 74196 37924 74208
rect 37976 74196 37982 74248
rect 23290 74128 23296 74180
rect 23348 74168 23354 74180
rect 33686 74168 33692 74180
rect 23348 74140 33692 74168
rect 23348 74128 23354 74140
rect 33686 74128 33692 74140
rect 33744 74128 33750 74180
rect 342346 73992 342352 74044
rect 342404 74032 342410 74044
rect 414014 74032 414020 74044
rect 342404 74004 414020 74032
rect 342404 73992 342410 74004
rect 414014 73992 414020 74004
rect 414072 73992 414078 74044
rect 79410 73924 79416 73976
rect 79468 73964 79474 73976
rect 322198 73964 322204 73976
rect 79468 73936 322204 73964
rect 79468 73924 79474 73936
rect 322198 73924 322204 73936
rect 322256 73924 322262 73976
rect 322290 73924 322296 73976
rect 322348 73964 322354 73976
rect 359090 73964 359096 73976
rect 322348 73936 359096 73964
rect 322348 73924 322354 73936
rect 359090 73924 359096 73936
rect 359148 73924 359154 73976
rect 408586 73924 408592 73976
rect 408644 73964 408650 73976
rect 568758 73964 568764 73976
rect 408644 73936 568764 73964
rect 408644 73924 408650 73936
rect 568758 73924 568764 73936
rect 568816 73924 568822 73976
rect 119890 73856 119896 73908
rect 119948 73896 119954 73908
rect 366266 73896 366272 73908
rect 119948 73868 366272 73896
rect 119948 73856 119954 73868
rect 366266 73856 366272 73868
rect 366324 73856 366330 73908
rect 390554 73856 390560 73908
rect 390612 73896 390618 73908
rect 570046 73896 570052 73908
rect 390612 73868 570052 73896
rect 390612 73856 390618 73868
rect 570046 73856 570052 73868
rect 570104 73856 570110 73908
rect 226426 73788 226432 73840
rect 226484 73828 226490 73840
rect 485590 73828 485596 73840
rect 226484 73800 485596 73828
rect 226484 73788 226490 73800
rect 485590 73788 485596 73800
rect 485648 73788 485654 73840
rect 507026 73788 507032 73840
rect 507084 73828 507090 73840
rect 534074 73828 534080 73840
rect 507084 73800 534080 73828
rect 507084 73788 507090 73800
rect 534074 73788 534080 73800
rect 534132 73788 534138 73840
rect 14826 73108 14832 73160
rect 14884 73148 14890 73160
rect 180058 73148 180064 73160
rect 14884 73120 180064 73148
rect 14884 73108 14890 73120
rect 180058 73108 180064 73120
rect 180116 73108 180122 73160
rect 301866 73108 301872 73160
rect 301924 73148 301930 73160
rect 322106 73148 322112 73160
rect 301924 73120 322112 73148
rect 301924 73108 301930 73120
rect 322106 73108 322112 73120
rect 322164 73148 322170 73160
rect 322290 73148 322296 73160
rect 322164 73120 322296 73148
rect 322164 73108 322170 73120
rect 322290 73108 322296 73120
rect 322348 73108 322354 73160
rect 435358 73108 435364 73160
rect 435416 73148 435422 73160
rect 572990 73148 572996 73160
rect 435416 73120 572996 73148
rect 435416 73108 435422 73120
rect 572990 73108 572996 73120
rect 573048 73108 573054 73160
rect 17862 73040 17868 73092
rect 17920 73080 17926 73092
rect 174538 73080 174544 73092
rect 17920 73052 174544 73080
rect 17920 73040 17926 73052
rect 174538 73040 174544 73052
rect 174596 73040 174602 73092
rect 445018 73040 445024 73092
rect 445076 73080 445082 73092
rect 575658 73080 575664 73092
rect 445076 73052 575664 73080
rect 445076 73040 445082 73052
rect 575658 73040 575664 73052
rect 575716 73040 575722 73092
rect 14918 72972 14924 73024
rect 14976 73012 14982 73024
rect 159358 73012 159364 73024
rect 14976 72984 159364 73012
rect 14976 72972 14982 72984
rect 159358 72972 159364 72984
rect 159416 72972 159422 73024
rect 450538 72972 450544 73024
rect 450596 73012 450602 73024
rect 578234 73012 578240 73024
rect 450596 72984 578240 73012
rect 450596 72972 450602 72984
rect 578234 72972 578240 72984
rect 578292 72972 578298 73024
rect 23474 72904 23480 72956
rect 23532 72944 23538 72956
rect 164234 72944 164240 72956
rect 23532 72916 164240 72944
rect 23532 72904 23538 72916
rect 164234 72904 164240 72916
rect 164292 72904 164298 72956
rect 459554 72904 459560 72956
rect 459612 72944 459618 72956
rect 460290 72944 460296 72956
rect 459612 72916 460296 72944
rect 459612 72904 459618 72916
rect 460290 72904 460296 72916
rect 460348 72944 460354 72956
rect 574370 72944 574376 72956
rect 460348 72916 574376 72944
rect 460348 72904 460354 72916
rect 574370 72904 574376 72916
rect 574428 72904 574434 72956
rect 17494 72836 17500 72888
rect 17552 72876 17558 72888
rect 155218 72876 155224 72888
rect 17552 72848 155224 72876
rect 17552 72836 17558 72848
rect 155218 72836 155224 72848
rect 155276 72836 155282 72888
rect 490558 72836 490564 72888
rect 490616 72876 490622 72888
rect 575750 72876 575756 72888
rect 490616 72848 575756 72876
rect 490616 72836 490622 72848
rect 575750 72836 575756 72848
rect 575808 72836 575814 72888
rect 534074 72768 534080 72820
rect 534132 72808 534138 72820
rect 579614 72808 579620 72820
rect 534132 72780 579620 72808
rect 534132 72768 534138 72780
rect 579614 72768 579620 72780
rect 579672 72768 579678 72820
rect 211706 72632 211712 72684
rect 211764 72672 211770 72684
rect 288618 72672 288624 72684
rect 211764 72644 288624 72672
rect 211764 72632 211770 72644
rect 288618 72632 288624 72644
rect 288676 72632 288682 72684
rect 134426 72564 134432 72616
rect 134484 72604 134490 72616
rect 371786 72604 371792 72616
rect 134484 72576 371792 72604
rect 134484 72564 134490 72576
rect 371786 72564 371792 72576
rect 371844 72564 371850 72616
rect 254026 72496 254032 72548
rect 254084 72536 254090 72548
rect 529934 72536 529940 72548
rect 254084 72508 529940 72536
rect 254084 72496 254090 72508
rect 529934 72496 529940 72508
rect 529992 72496 529998 72548
rect 164234 72428 164240 72480
rect 164292 72468 164298 72480
rect 164786 72468 164792 72480
rect 164292 72440 164792 72468
rect 164292 72428 164298 72440
rect 164786 72428 164792 72440
rect 164844 72428 164850 72480
rect 169846 72428 169852 72480
rect 169904 72468 169910 72480
rect 459554 72468 459560 72480
rect 169904 72440 459560 72468
rect 169904 72428 169910 72440
rect 459554 72428 459560 72440
rect 459612 72428 459618 72480
rect 15010 71680 15016 71732
rect 15068 71720 15074 71732
rect 140038 71720 140044 71732
rect 15068 71692 140044 71720
rect 15068 71680 15074 71692
rect 140038 71680 140044 71692
rect 140096 71680 140102 71732
rect 439590 71680 439596 71732
rect 439648 71720 439654 71732
rect 571610 71720 571616 71732
rect 439648 71692 571616 71720
rect 439648 71680 439654 71692
rect 571610 71680 571616 71692
rect 571668 71680 571674 71732
rect 25590 71612 25596 71664
rect 25648 71652 25654 71664
rect 124582 71652 124588 71664
rect 25648 71624 124588 71652
rect 25648 71612 25654 71624
rect 124582 71612 124588 71624
rect 124640 71652 124646 71664
rect 125502 71652 125508 71664
rect 124640 71624 125508 71652
rect 124640 71612 124646 71624
rect 125502 71612 125508 71624
rect 125560 71612 125566 71664
rect 469858 71612 469864 71664
rect 469916 71652 469922 71664
rect 470410 71652 470416 71664
rect 469916 71624 470416 71652
rect 469916 71612 469922 71624
rect 470410 71612 470416 71624
rect 470468 71652 470474 71664
rect 572714 71652 572720 71664
rect 470468 71624 572720 71652
rect 470468 71612 470474 71624
rect 572714 71612 572720 71624
rect 572772 71612 572778 71664
rect 22002 71544 22008 71596
rect 22060 71584 22066 71596
rect 109126 71584 109132 71596
rect 22060 71556 109132 71584
rect 22060 71544 22066 71556
rect 109126 71544 109132 71556
rect 109184 71544 109190 71596
rect 475378 71544 475384 71596
rect 475436 71584 475442 71596
rect 575842 71584 575848 71596
rect 475436 71556 575848 71584
rect 475436 71544 475442 71556
rect 575842 71544 575848 71556
rect 575900 71544 575906 71596
rect 496078 71476 496084 71528
rect 496136 71516 496142 71528
rect 574094 71516 574100 71528
rect 496136 71488 574100 71516
rect 496136 71476 496142 71488
rect 574094 71476 574100 71488
rect 574152 71476 574158 71528
rect 500770 71408 500776 71460
rect 500828 71448 500834 71460
rect 575934 71448 575940 71460
rect 500828 71420 575940 71448
rect 500828 71408 500834 71420
rect 575934 71408 575940 71420
rect 575992 71408 575998 71460
rect 262122 71340 262128 71392
rect 262180 71380 262186 71392
rect 289906 71380 289912 71392
rect 262180 71352 289912 71380
rect 262180 71340 262186 71352
rect 289906 71340 289912 71352
rect 289964 71340 289970 71392
rect 239398 71272 239404 71324
rect 239456 71312 239462 71324
rect 292758 71312 292764 71324
rect 239456 71284 292764 71312
rect 239456 71272 239462 71284
rect 292758 71272 292764 71284
rect 292816 71272 292822 71324
rect 248414 71204 248420 71256
rect 248472 71244 248478 71256
rect 261386 71244 261392 71256
rect 248472 71216 261392 71244
rect 248472 71204 248478 71216
rect 261386 71204 261392 71216
rect 261444 71244 261450 71256
rect 262122 71244 262128 71256
rect 261444 71216 262128 71244
rect 261444 71204 261450 71216
rect 262122 71204 262128 71216
rect 262180 71204 262186 71256
rect 288986 71204 288992 71256
rect 289044 71244 289050 71256
rect 423674 71244 423680 71256
rect 289044 71216 423680 71244
rect 289044 71204 289050 71216
rect 423674 71204 423680 71216
rect 423732 71204 423738 71256
rect 114462 71136 114468 71188
rect 114520 71176 114526 71188
rect 364426 71176 364432 71188
rect 114520 71148 364432 71176
rect 114520 71136 114526 71148
rect 364426 71136 364432 71148
rect 364484 71136 364490 71188
rect 94314 71068 94320 71120
rect 94372 71108 94378 71120
rect 357434 71108 357440 71120
rect 94372 71080 357440 71108
rect 94372 71068 94378 71080
rect 357434 71068 357440 71080
rect 357492 71068 357498 71120
rect 33686 71000 33692 71052
rect 33744 71040 33750 71052
rect 303706 71040 303712 71052
rect 33744 71012 303712 71040
rect 33744 71000 33750 71012
rect 303706 71000 303712 71012
rect 303764 71000 303770 71052
rect 331214 71000 331220 71052
rect 331272 71040 331278 71052
rect 384390 71040 384396 71052
rect 331272 71012 384396 71040
rect 331272 71000 331278 71012
rect 384390 71000 384396 71012
rect 384448 71000 384454 71052
rect 109126 70388 109132 70440
rect 109184 70428 109190 70440
rect 109678 70428 109684 70440
rect 109184 70400 109684 70428
rect 109184 70388 109190 70400
rect 109678 70388 109684 70400
rect 109736 70388 109742 70440
rect 296530 70320 296536 70372
rect 296588 70360 296594 70372
rect 331214 70360 331220 70372
rect 296588 70332 331220 70360
rect 296588 70320 296594 70332
rect 331214 70320 331220 70332
rect 331272 70320 331278 70372
rect 405642 70320 405648 70372
rect 405700 70360 405706 70372
rect 578326 70360 578332 70372
rect 405700 70332 578332 70360
rect 405700 70320 405706 70332
rect 578326 70320 578332 70332
rect 578384 70320 578390 70372
rect 237466 69912 237472 69964
rect 237524 69952 237530 69964
rect 239490 69952 239496 69964
rect 237524 69924 239496 69952
rect 237524 69912 237530 69924
rect 239490 69912 239496 69924
rect 239548 69912 239554 69964
rect 264882 69844 264888 69896
rect 264940 69884 264946 69896
rect 269114 69884 269120 69896
rect 264940 69856 269120 69884
rect 264940 69844 264946 69856
rect 269114 69844 269120 69856
rect 269172 69884 269178 69896
rect 291194 69884 291200 69896
rect 269172 69856 291200 69884
rect 269172 69844 269178 69856
rect 291194 69844 291200 69856
rect 291252 69844 291258 69896
rect 317322 69844 317328 69896
rect 317380 69884 317386 69896
rect 343910 69884 343916 69896
rect 317380 69856 343916 69884
rect 317380 69844 317386 69856
rect 343910 69844 343916 69856
rect 343968 69844 343974 69896
rect 125502 69776 125508 69828
rect 125560 69816 125566 69828
rect 368474 69816 368480 69828
rect 125560 69788 368480 69816
rect 125560 69776 125566 69788
rect 368474 69776 368480 69788
rect 368532 69776 368538 69828
rect 59262 69708 59268 69760
rect 59320 69748 59326 69760
rect 313366 69748 313372 69760
rect 59320 69720 313372 69748
rect 59320 69708 59326 69720
rect 313366 69708 313372 69720
rect 313424 69708 313430 69760
rect 338114 69708 338120 69760
rect 338172 69748 338178 69760
rect 404446 69748 404452 69760
rect 338172 69720 404452 69748
rect 338172 69708 338178 69720
rect 404446 69708 404452 69720
rect 404504 69748 404510 69760
rect 405642 69748 405648 69760
rect 404504 69720 405648 69748
rect 404504 69708 404510 69720
rect 405642 69708 405648 69720
rect 405700 69708 405706 69760
rect 410426 69708 410432 69760
rect 410484 69748 410490 69760
rect 556430 69748 556436 69760
rect 410484 69720 556436 69748
rect 410484 69708 410490 69720
rect 556430 69708 556436 69720
rect 556488 69708 556494 69760
rect 12342 69640 12348 69692
rect 12400 69680 12406 69692
rect 40678 69680 40684 69692
rect 12400 69652 40684 69680
rect 12400 69640 12406 69652
rect 40678 69640 40684 69652
rect 40736 69640 40742 69692
rect 252554 69640 252560 69692
rect 252612 69680 252618 69692
rect 526070 69680 526076 69692
rect 252612 69652 526076 69680
rect 252612 69640 252618 69652
rect 526070 69640 526076 69652
rect 526128 69640 526134 69692
rect 25498 68960 25504 69012
rect 25556 69000 25562 69012
rect 184934 69000 184940 69012
rect 25556 68972 184940 69000
rect 25556 68960 25562 68972
rect 184934 68960 184940 68972
rect 184992 68960 184998 69012
rect 300762 68960 300768 69012
rect 300820 69000 300826 69012
rect 316586 69000 316592 69012
rect 300820 68972 316592 69000
rect 300820 68960 300826 68972
rect 316586 68960 316592 68972
rect 316644 69000 316650 69012
rect 317322 69000 317328 69012
rect 316644 68972 317328 69000
rect 316644 68960 316650 68972
rect 317322 68960 317328 68972
rect 317380 68960 317386 69012
rect 409138 68960 409144 69012
rect 409196 69000 409202 69012
rect 574462 69000 574468 69012
rect 409196 68972 574468 69000
rect 409196 68960 409202 68972
rect 574462 68960 574468 68972
rect 574520 68960 574526 69012
rect 195146 68552 195152 68604
rect 195204 68592 195210 68604
rect 284938 68592 284944 68604
rect 195204 68564 284944 68592
rect 195204 68552 195210 68564
rect 284938 68552 284944 68564
rect 284996 68552 285002 68604
rect 149974 68484 149980 68536
rect 150032 68524 150038 68536
rect 272426 68524 272432 68536
rect 150032 68496 272432 68524
rect 150032 68484 150038 68496
rect 272426 68484 272432 68496
rect 272484 68484 272490 68536
rect 276106 68484 276112 68536
rect 276164 68524 276170 68536
rect 375466 68524 375472 68536
rect 276164 68496 375472 68524
rect 276164 68484 276170 68496
rect 375466 68484 375472 68496
rect 375524 68484 375530 68536
rect 265618 68416 265624 68468
rect 265676 68456 265682 68468
rect 520274 68456 520280 68468
rect 265676 68428 520280 68456
rect 265676 68416 265682 68428
rect 520274 68416 520280 68428
rect 520332 68416 520338 68468
rect 84102 68348 84108 68400
rect 84160 68388 84166 68400
rect 353386 68388 353392 68400
rect 84160 68360 353392 68388
rect 84160 68348 84166 68360
rect 353386 68348 353392 68360
rect 353444 68348 353450 68400
rect 234430 68280 234436 68332
rect 234488 68320 234494 68332
rect 244826 68320 244832 68332
rect 234488 68292 244832 68320
rect 234488 68280 234494 68292
rect 244826 68280 244832 68292
rect 244884 68280 244890 68332
rect 258074 68280 258080 68332
rect 258132 68320 258138 68332
rect 541250 68320 541256 68332
rect 258132 68292 541256 68320
rect 258132 68280 258138 68292
rect 541250 68280 541256 68292
rect 541308 68280 541314 68332
rect 217318 67532 217324 67584
rect 217376 67572 217382 67584
rect 240778 67572 240784 67584
rect 217376 67544 240784 67572
rect 217376 67532 217382 67544
rect 240778 67532 240784 67544
rect 240836 67532 240842 67584
rect 244826 67532 244832 67584
rect 244884 67572 244890 67584
rect 287790 67572 287796 67584
rect 244884 67544 287796 67572
rect 244884 67532 244890 67544
rect 287790 67532 287796 67544
rect 287848 67532 287854 67584
rect 335998 67532 336004 67584
rect 336056 67572 336062 67584
rect 393314 67572 393320 67584
rect 336056 67544 393320 67572
rect 336056 67532 336062 67544
rect 393314 67532 393320 67544
rect 393372 67532 393378 67584
rect 261478 67464 261484 67516
rect 261536 67504 261542 67516
rect 265066 67504 265072 67516
rect 261536 67476 265072 67504
rect 261536 67464 261542 67476
rect 265066 67464 265072 67476
rect 265124 67464 265130 67516
rect 265066 67056 265072 67108
rect 265124 67096 265130 67108
rect 294046 67096 294052 67108
rect 265124 67068 294052 67096
rect 265124 67056 265130 67068
rect 294046 67056 294052 67068
rect 294104 67056 294110 67108
rect 231946 66988 231952 67040
rect 232004 67028 232010 67040
rect 500770 67028 500776 67040
rect 232004 67000 500776 67028
rect 232004 66988 232010 67000
rect 500770 66988 500776 67000
rect 500828 66988 500834 67040
rect 73798 66920 73804 66972
rect 73856 66960 73862 66972
rect 349706 66960 349712 66972
rect 73856 66932 349712 66960
rect 73856 66920 73862 66932
rect 349706 66920 349712 66932
rect 349764 66920 349770 66972
rect 255866 66852 255872 66904
rect 255924 66892 255930 66904
rect 536098 66892 536104 66904
rect 255924 66864 536104 66892
rect 255924 66852 255930 66864
rect 536098 66852 536104 66864
rect 536156 66852 536162 66904
rect 335354 66784 335360 66836
rect 335412 66824 335418 66836
rect 335998 66824 336004 66836
rect 335412 66796 336004 66824
rect 335412 66784 335418 66796
rect 335998 66784 336004 66796
rect 336056 66784 336062 66836
rect 219526 65628 219532 65680
rect 219584 65668 219590 65680
rect 242986 65668 242992 65680
rect 219584 65640 242992 65668
rect 219584 65628 219590 65640
rect 242986 65628 242992 65640
rect 243044 65628 243050 65680
rect 271138 65628 271144 65680
rect 271196 65668 271202 65680
rect 480254 65668 480260 65680
rect 271196 65640 480260 65668
rect 271196 65628 271202 65640
rect 480254 65628 480260 65640
rect 480312 65628 480318 65680
rect 228266 65560 228272 65612
rect 228324 65600 228330 65612
rect 490558 65600 490564 65612
rect 228324 65572 490564 65600
rect 228324 65560 228330 65572
rect 490558 65560 490564 65572
rect 490616 65560 490622 65612
rect 187786 65492 187792 65544
rect 187844 65532 187850 65544
rect 194594 65532 194600 65544
rect 187844 65504 194600 65532
rect 187844 65492 187850 65504
rect 194594 65492 194600 65504
rect 194652 65492 194658 65544
rect 209774 65492 209780 65544
rect 209832 65532 209838 65544
rect 226978 65532 226984 65544
rect 209832 65504 226984 65532
rect 209832 65492 209838 65504
rect 226978 65492 226984 65504
rect 227036 65492 227042 65544
rect 230474 65492 230480 65544
rect 230532 65532 230538 65544
rect 496078 65532 496084 65544
rect 230532 65504 496084 65532
rect 230532 65492 230538 65504
rect 496078 65492 496084 65504
rect 496136 65492 496142 65544
rect 242986 64948 242992 65000
rect 243044 64988 243050 65000
rect 243814 64988 243820 65000
rect 243044 64960 243820 64988
rect 243044 64948 243050 64960
rect 243814 64948 243820 64960
rect 243872 64948 243878 65000
rect 243814 64812 243820 64864
rect 243872 64852 243878 64864
rect 293954 64852 293960 64864
rect 243872 64824 293960 64852
rect 243872 64812 243878 64824
rect 293954 64812 293960 64824
rect 294012 64812 294018 64864
rect 40678 64268 40684 64320
rect 40736 64308 40742 64320
rect 178678 64308 178684 64320
rect 40736 64280 178684 64308
rect 40736 64268 40742 64280
rect 178678 64268 178684 64280
rect 178736 64268 178742 64320
rect 206278 64268 206284 64320
rect 206336 64308 206342 64320
rect 465718 64308 465724 64320
rect 206336 64280 465724 64308
rect 206336 64268 206342 64280
rect 465718 64268 465724 64280
rect 465776 64268 465782 64320
rect 173066 64200 173072 64252
rect 173124 64240 173130 64252
rect 469858 64240 469864 64252
rect 173124 64212 469864 64240
rect 173124 64200 173130 64212
rect 469858 64200 469864 64212
rect 469916 64200 469922 64252
rect 175274 64132 175280 64184
rect 175332 64172 175338 64184
rect 475378 64172 475384 64184
rect 175332 64144 475384 64172
rect 175332 64132 175338 64144
rect 475378 64132 475384 64144
rect 475436 64132 475442 64184
rect 297910 63044 297916 63096
rect 297968 63084 297974 63096
rect 329834 63084 329840 63096
rect 297968 63056 329840 63084
rect 297968 63044 297974 63056
rect 329834 63044 329840 63056
rect 329892 63044 329898 63096
rect 303062 62976 303068 63028
rect 303120 63016 303126 63028
rect 324314 63016 324320 63028
rect 303120 62988 324320 63016
rect 303120 62976 303126 62988
rect 324314 62976 324320 62988
rect 324372 63016 324378 63028
rect 362954 63016 362960 63028
rect 324372 62988 362960 63016
rect 324372 62976 324378 62988
rect 362954 62976 362960 62988
rect 363012 62976 363018 63028
rect 203518 62908 203524 62960
rect 203576 62948 203582 62960
rect 445018 62948 445024 62960
rect 203576 62920 445024 62948
rect 203576 62908 203582 62920
rect 445018 62908 445024 62920
rect 445076 62908 445082 62960
rect 154666 62840 154672 62892
rect 154724 62880 154730 62892
rect 435358 62880 435364 62892
rect 154724 62852 435364 62880
rect 154724 62840 154730 62852
rect 435358 62840 435364 62852
rect 435416 62840 435422 62892
rect 156506 62772 156512 62824
rect 156564 62812 156570 62824
rect 439590 62812 439596 62824
rect 156564 62784 439596 62812
rect 156564 62772 156570 62784
rect 439590 62772 439596 62784
rect 439648 62772 439654 62824
rect 299290 62024 299296 62076
rect 299348 62064 299354 62076
rect 328454 62064 328460 62076
rect 299348 62036 328460 62064
rect 299348 62024 299354 62036
rect 328454 62024 328460 62036
rect 328512 62024 328518 62076
rect 329098 62024 329104 62076
rect 329156 62064 329162 62076
rect 373994 62064 374000 62076
rect 329156 62036 374000 62064
rect 329156 62024 329162 62036
rect 373994 62024 374000 62036
rect 374052 62024 374058 62076
rect 300670 61616 300676 61668
rect 300728 61656 300734 61668
rect 325878 61656 325884 61668
rect 300728 61628 325884 61656
rect 300728 61616 300734 61628
rect 325878 61616 325884 61628
rect 325936 61616 325942 61668
rect 308398 61548 308404 61600
rect 308456 61588 308462 61600
rect 415946 61588 415952 61600
rect 308456 61560 415952 61588
rect 308456 61548 308462 61560
rect 415946 61548 415952 61560
rect 416004 61548 416010 61600
rect 116578 61480 116584 61532
rect 116636 61520 116642 61532
rect 309226 61520 309232 61532
rect 116636 61492 309232 61520
rect 116636 61480 116642 61492
rect 309226 61480 309232 61492
rect 309284 61480 309290 61532
rect 309778 61480 309784 61532
rect 309836 61520 309842 61532
rect 338206 61520 338212 61532
rect 309836 61492 338212 61520
rect 309836 61480 309842 61492
rect 338206 61480 338212 61492
rect 338264 61480 338270 61532
rect 52454 61412 52460 61464
rect 52512 61452 52518 61464
rect 311066 61452 311072 61464
rect 52512 61424 311072 61452
rect 52512 61412 52518 61424
rect 311066 61412 311072 61424
rect 311124 61412 311130 61464
rect 3510 61344 3516 61396
rect 3568 61384 3574 61396
rect 13078 61384 13084 61396
rect 3568 61356 13084 61384
rect 3568 61344 3574 61356
rect 13078 61344 13084 61356
rect 13136 61344 13142 61396
rect 43438 61344 43444 61396
rect 43496 61384 43502 61396
rect 307754 61384 307760 61396
rect 43496 61356 307760 61384
rect 43496 61344 43502 61356
rect 307754 61344 307760 61356
rect 307812 61344 307818 61396
rect 325878 61344 325884 61396
rect 325936 61384 325942 61396
rect 368566 61384 368572 61396
rect 325936 61356 368572 61384
rect 325936 61344 325942 61356
rect 368566 61344 368572 61356
rect 368624 61344 368630 61396
rect 412634 61344 412640 61396
rect 412692 61384 412698 61396
rect 560938 61384 560944 61396
rect 412692 61356 560944 61384
rect 412692 61344 412698 61356
rect 560938 61344 560944 61356
rect 560996 61344 561002 61396
rect 298830 60732 298836 60784
rect 298888 60772 298894 60784
rect 299290 60772 299296 60784
rect 298888 60744 299296 60772
rect 298888 60732 298894 60744
rect 299290 60732 299296 60744
rect 299348 60732 299354 60784
rect 297450 60324 297456 60376
rect 297508 60364 297514 60376
rect 313274 60364 313280 60376
rect 297508 60336 313280 60364
rect 297508 60324 297514 60336
rect 313274 60324 313280 60336
rect 313332 60324 313338 60376
rect 340874 60324 340880 60376
rect 340932 60364 340938 60376
rect 409138 60364 409144 60376
rect 340932 60336 409144 60364
rect 340932 60324 340938 60336
rect 409138 60324 409144 60336
rect 409196 60324 409202 60376
rect 298738 60256 298744 60308
rect 298796 60296 298802 60308
rect 396074 60296 396080 60308
rect 298796 60268 396080 60296
rect 298796 60256 298802 60268
rect 396074 60256 396080 60268
rect 396132 60256 396138 60308
rect 295978 60188 295984 60240
rect 296036 60228 296042 60240
rect 397546 60228 397552 60240
rect 296036 60200 397552 60228
rect 296036 60188 296042 60200
rect 397546 60188 397552 60200
rect 397604 60188 397610 60240
rect 109678 60120 109684 60172
rect 109736 60160 109742 60172
rect 362954 60160 362960 60172
rect 109736 60132 362960 60160
rect 109736 60120 109742 60132
rect 362954 60120 362960 60132
rect 363012 60120 363018 60172
rect 104158 60052 104164 60104
rect 104216 60092 104222 60104
rect 360746 60092 360752 60104
rect 104216 60064 360752 60092
rect 104216 60052 104222 60064
rect 360746 60052 360752 60064
rect 360804 60052 360810 60104
rect 98638 59984 98644 60036
rect 98696 60024 98702 60036
rect 358906 60024 358912 60036
rect 98696 59996 358912 60024
rect 98696 59984 98702 59996
rect 358906 59984 358912 59996
rect 358964 59984 358970 60036
rect 336734 59304 336740 59356
rect 336792 59344 336798 59356
rect 398926 59344 398932 59356
rect 336792 59316 398932 59344
rect 336792 59304 336798 59316
rect 398926 59304 398932 59316
rect 398984 59304 398990 59356
rect 140038 58760 140044 58812
rect 140096 58800 140102 58812
rect 373994 58800 374000 58812
rect 140096 58772 374000 58800
rect 140096 58760 140102 58772
rect 373994 58760 374000 58772
rect 374052 58760 374058 58812
rect 432506 58760 432512 58812
rect 432564 58800 432570 58812
rect 565814 58800 565820 58812
rect 432564 58772 565820 58800
rect 432564 58760 432570 58772
rect 565814 58760 565820 58772
rect 565872 58760 565878 58812
rect 88978 58692 88984 58744
rect 89036 58732 89042 58744
rect 355226 58732 355232 58744
rect 89036 58704 355232 58732
rect 89036 58692 89042 58704
rect 355226 58692 355232 58704
rect 355284 58692 355290 58744
rect 355318 58692 355324 58744
rect 355376 58732 355382 58744
rect 511258 58732 511264 58744
rect 355376 58704 511264 58732
rect 355376 58692 355382 58704
rect 511258 58692 511264 58704
rect 511316 58692 511322 58744
rect 68278 58624 68284 58676
rect 68336 58664 68342 58676
rect 347866 58664 347872 58676
rect 68336 58636 347872 58664
rect 68336 58624 68342 58636
rect 347866 58624 347872 58636
rect 347924 58624 347930 58676
rect 392026 58624 392032 58676
rect 392084 58664 392090 58676
rect 550634 58664 550640 58676
rect 392084 58636 550640 58664
rect 392084 58624 392090 58636
rect 550634 58624 550640 58636
rect 550692 58624 550698 58676
rect 329834 57876 329840 57928
rect 329892 57916 329898 57928
rect 378134 57916 378140 57928
rect 329892 57888 378140 57916
rect 329892 57876 329898 57888
rect 378134 57876 378140 57888
rect 378192 57876 378198 57928
rect 294598 57468 294604 57520
rect 294656 57508 294662 57520
rect 383194 57508 383200 57520
rect 294656 57480 383200 57508
rect 294656 57468 294662 57480
rect 383194 57468 383200 57480
rect 383252 57468 383258 57520
rect 128998 57400 129004 57452
rect 129056 57440 129062 57452
rect 370314 57440 370320 57452
rect 129056 57412 370320 57440
rect 129056 57400 129062 57412
rect 370314 57400 370320 57412
rect 370372 57400 370378 57452
rect 37918 57332 37924 57384
rect 37976 57372 37982 57384
rect 305914 57372 305920 57384
rect 37976 57344 305920 57372
rect 37976 57332 37982 57344
rect 305914 57332 305920 57344
rect 305972 57332 305978 57384
rect 64138 57264 64144 57316
rect 64196 57304 64202 57316
rect 346394 57304 346400 57316
rect 64196 57276 346400 57304
rect 64196 57264 64202 57276
rect 346394 57264 346400 57276
rect 346452 57264 346458 57316
rect 259914 57196 259920 57248
rect 259972 57236 259978 57248
rect 545758 57236 545764 57248
rect 259972 57208 545764 57236
rect 259972 57196 259978 57208
rect 545758 57196 545764 57208
rect 545816 57196 545822 57248
rect 299382 56516 299388 56568
rect 299440 56556 299446 56568
rect 319438 56556 319444 56568
rect 299440 56528 319444 56556
rect 299440 56516 299446 56528
rect 319438 56516 319444 56528
rect 319496 56516 319502 56568
rect 298554 56176 298560 56228
rect 298612 56216 298618 56228
rect 299382 56216 299388 56228
rect 298612 56188 299388 56216
rect 298612 56176 298618 56188
rect 299382 56176 299388 56188
rect 299440 56176 299446 56228
rect 294874 56108 294880 56160
rect 294932 56148 294938 56160
rect 307846 56148 307852 56160
rect 294932 56120 307852 56148
rect 294932 56108 294938 56120
rect 307846 56108 307852 56120
rect 307904 56108 307910 56160
rect 318794 56148 318800 56160
rect 316006 56120 318800 56148
rect 303246 56040 303252 56092
rect 303304 56080 303310 56092
rect 316006 56080 316034 56120
rect 318794 56108 318800 56120
rect 318852 56148 318858 56160
rect 347774 56148 347780 56160
rect 318852 56120 347780 56148
rect 318852 56108 318858 56120
rect 347774 56108 347780 56120
rect 347832 56108 347838 56160
rect 303304 56052 316034 56080
rect 303304 56040 303310 56052
rect 320634 56040 320640 56092
rect 320692 56080 320698 56092
rect 353294 56080 353300 56092
rect 320692 56052 353300 56080
rect 320692 56040 320698 56052
rect 353294 56040 353300 56052
rect 353352 56040 353358 56092
rect 169754 55972 169760 56024
rect 169812 56012 169818 56024
rect 178954 56012 178960 56024
rect 169812 55984 178960 56012
rect 169812 55972 169818 55984
rect 178954 55972 178960 55984
rect 179012 55972 179018 56024
rect 235902 55972 235908 56024
rect 235960 56012 235966 56024
rect 247034 56012 247040 56024
rect 235960 55984 247040 56012
rect 235960 55972 235966 55984
rect 247034 55972 247040 55984
rect 247092 55972 247098 56024
rect 256602 55972 256608 56024
rect 256660 56012 256666 56024
rect 267274 56012 267280 56024
rect 256660 55984 267280 56012
rect 256660 55972 256666 55984
rect 267274 55972 267280 55984
rect 267332 55972 267338 56024
rect 281442 55972 281448 56024
rect 281500 56012 281506 56024
rect 294598 56012 294604 56024
rect 281500 55984 294604 56012
rect 281500 55972 281506 55984
rect 294598 55972 294604 55984
rect 294656 55972 294662 56024
rect 298002 55972 298008 56024
rect 298060 56012 298066 56024
rect 320652 56012 320680 56040
rect 298060 55984 320680 56012
rect 298060 55972 298066 55984
rect 344554 55972 344560 56024
rect 344612 56012 344618 56024
rect 420178 56012 420184 56024
rect 344612 55984 420184 56012
rect 344612 55972 344618 55984
rect 420178 55972 420184 55984
rect 420236 55972 420242 56024
rect 166074 55904 166080 55956
rect 166132 55944 166138 55956
rect 450538 55944 450544 55956
rect 166132 55916 450544 55944
rect 166132 55904 166138 55916
rect 450538 55904 450544 55916
rect 450596 55904 450602 55956
rect 167914 55836 167920 55888
rect 167972 55876 167978 55888
rect 454034 55876 454040 55888
rect 167972 55848 454040 55876
rect 167972 55836 167978 55848
rect 454034 55836 454040 55848
rect 454092 55836 454098 55888
rect 226978 55156 226984 55208
rect 227036 55196 227042 55208
rect 239398 55196 239404 55208
rect 227036 55168 239404 55196
rect 227036 55156 227042 55168
rect 239398 55156 239404 55168
rect 239456 55156 239462 55208
rect 278314 54816 278320 54868
rect 278372 54856 278378 54868
rect 288434 54856 288440 54868
rect 278372 54828 288440 54856
rect 278372 54816 278378 54828
rect 288434 54816 288440 54828
rect 288492 54816 288498 54868
rect 296438 54816 296444 54868
rect 296496 54856 296502 54868
rect 296496 54828 300440 54856
rect 296496 54816 296502 54828
rect 300412 54800 300440 54828
rect 178678 54748 178684 54800
rect 178736 54788 178742 54800
rect 178736 54760 190454 54788
rect 178736 54748 178742 54760
rect 174538 54680 174544 54732
rect 174596 54720 174602 54732
rect 180794 54720 180800 54732
rect 174596 54692 180800 54720
rect 174596 54680 174602 54692
rect 180794 54680 180800 54692
rect 180852 54680 180858 54732
rect 180058 54612 180064 54664
rect 180116 54652 180122 54664
rect 182634 54652 182640 54664
rect 180116 54624 182640 54652
rect 180116 54612 180122 54624
rect 182634 54612 182640 54624
rect 182692 54612 182698 54664
rect 190426 54652 190454 54760
rect 281994 54748 282000 54800
rect 282052 54788 282058 54800
rect 287606 54788 287612 54800
rect 282052 54760 287612 54788
rect 282052 54748 282058 54760
rect 287606 54748 287612 54760
rect 287664 54748 287670 54800
rect 297358 54748 297364 54800
rect 297416 54788 297422 54800
rect 297416 54760 297588 54788
rect 297416 54748 297422 54760
rect 240042 54680 240048 54732
rect 240100 54720 240106 54732
rect 248874 54720 248880 54732
rect 240100 54692 248880 54720
rect 240100 54680 240106 54692
rect 248874 54680 248880 54692
rect 248932 54680 248938 54732
rect 250714 54680 250720 54732
rect 250772 54720 250778 54732
rect 265618 54720 265624 54732
rect 250772 54692 265624 54720
rect 250772 54680 250778 54692
rect 265618 54680 265624 54692
rect 265676 54680 265682 54732
rect 274634 54680 274640 54732
rect 274692 54720 274698 54732
rect 289814 54720 289820 54732
rect 274692 54692 289820 54720
rect 274692 54680 274698 54692
rect 289814 54680 289820 54692
rect 289872 54680 289878 54732
rect 291194 54680 291200 54732
rect 291252 54720 291258 54732
rect 297450 54720 297456 54732
rect 291252 54692 297456 54720
rect 291252 54680 291258 54692
rect 297450 54680 297456 54692
rect 297508 54680 297514 54732
rect 297560 54720 297588 54760
rect 300394 54748 300400 54800
rect 300452 54788 300458 54800
rect 309778 54788 309784 54800
rect 300452 54760 309784 54788
rect 300452 54748 300458 54760
rect 309778 54748 309784 54760
rect 309836 54748 309842 54800
rect 322198 54748 322204 54800
rect 322256 54788 322262 54800
rect 351914 54788 351920 54800
rect 322256 54760 351920 54788
rect 322256 54748 322262 54760
rect 351914 54748 351920 54760
rect 351972 54748 351978 54800
rect 379514 54720 379520 54732
rect 297560 54692 379520 54720
rect 379514 54680 379520 54692
rect 379572 54680 379578 54732
rect 197354 54652 197360 54664
rect 190426 54624 197360 54652
rect 197354 54612 197360 54624
rect 197412 54612 197418 54664
rect 208394 54612 208400 54664
rect 208452 54652 208458 54664
rect 271138 54652 271144 54664
rect 208452 54624 271144 54652
rect 208452 54612 208458 54624
rect 271138 54612 271144 54624
rect 271196 54612 271202 54664
rect 276014 54612 276020 54664
rect 276072 54652 276078 54664
rect 394234 54652 394240 54664
rect 276072 54624 394240 54652
rect 276072 54612 276078 54624
rect 394234 54612 394240 54624
rect 394292 54612 394298 54664
rect 171594 54544 171600 54596
rect 171652 54584 171658 54596
rect 206278 54584 206284 54596
rect 171652 54556 206284 54584
rect 171652 54544 171658 54556
rect 206278 54544 206284 54556
rect 206336 54544 206342 54596
rect 235994 54544 236000 54596
rect 236052 54584 236058 54596
rect 355318 54584 355324 54596
rect 236052 54556 355324 54584
rect 236052 54544 236058 54556
rect 355318 54544 355324 54556
rect 355376 54544 355382 54596
rect 429194 54544 429200 54596
rect 429252 54584 429258 54596
rect 439498 54584 439504 54596
rect 429252 54556 439504 54584
rect 429252 54544 429258 54556
rect 439498 54544 439504 54556
rect 439556 54544 439562 54596
rect 158714 54476 158720 54528
rect 158772 54516 158778 54528
rect 203518 54516 203524 54528
rect 158772 54488 203524 54516
rect 158772 54476 158778 54488
rect 203518 54476 203524 54488
rect 203576 54476 203582 54528
rect 204254 54476 204260 54528
rect 204312 54516 204318 54528
rect 210234 54516 210240 54528
rect 204312 54488 210240 54516
rect 204312 54476 204318 54488
rect 210234 54476 210240 54488
rect 210292 54476 210298 54528
rect 282270 54516 282276 54528
rect 219406 54488 282276 54516
rect 159358 54408 159364 54460
rect 159416 54448 159422 54460
rect 162394 54448 162400 54460
rect 159416 54420 162400 54448
rect 159416 54408 159422 54420
rect 162394 54408 162400 54420
rect 162452 54408 162458 54460
rect 206554 54408 206560 54460
rect 206612 54448 206618 54460
rect 219406 54448 219434 54488
rect 282270 54476 282276 54488
rect 282328 54476 282334 54528
rect 294598 54476 294604 54528
rect 294656 54516 294662 54528
rect 414474 54516 414480 54528
rect 294656 54488 414480 54516
rect 294656 54476 294662 54488
rect 414474 54476 414480 54488
rect 414532 54476 414538 54528
rect 427354 54476 427360 54528
rect 427412 54516 427418 54528
rect 558178 54516 558184 54528
rect 427412 54488 558184 54516
rect 427412 54476 427418 54488
rect 558178 54476 558184 54488
rect 558236 54476 558242 54528
rect 206612 54420 219434 54448
rect 206612 54408 206618 54420
rect 285674 54272 285680 54324
rect 285732 54312 285738 54324
rect 289078 54312 289084 54324
rect 285732 54284 289084 54312
rect 285732 54272 285738 54284
rect 289078 54272 289084 54284
rect 289136 54272 289142 54324
rect 240778 53864 240784 53916
rect 240836 53904 240842 53916
rect 241514 53904 241520 53916
rect 240836 53876 241520 53904
rect 240836 53864 240842 53876
rect 241514 53864 241520 53876
rect 241572 53864 241578 53916
rect 155218 53796 155224 53848
rect 155276 53836 155282 53848
rect 160554 53836 160560 53848
rect 155276 53808 160560 53836
rect 155276 53796 155282 53808
rect 160554 53796 160560 53808
rect 160612 53796 160618 53848
rect 186314 53796 186320 53848
rect 186372 53836 186378 53848
rect 188338 53836 188344 53848
rect 186372 53808 188344 53836
rect 186372 53796 186378 53808
rect 188338 53796 188344 53808
rect 188396 53796 188402 53848
rect 221274 53796 221280 53848
rect 221332 53836 221338 53848
rect 285766 53836 285772 53848
rect 221332 53808 285772 53836
rect 221332 53796 221338 53808
rect 285766 53796 285772 53808
rect 285824 53796 285830 53848
rect 296714 53796 296720 53848
rect 296772 53836 296778 53848
rect 298830 53836 298836 53848
rect 296772 53808 298836 53836
rect 296772 53796 296778 53808
rect 298830 53796 298836 53808
rect 298888 53796 298894 53848
rect 327994 53796 328000 53848
rect 328052 53836 328058 53848
rect 329098 53836 329104 53848
rect 328052 53808 329104 53836
rect 328052 53796 328058 53808
rect 329098 53796 329104 53808
rect 329156 53796 329162 53848
rect 13262 53048 13268 53100
rect 13320 53088 13326 53100
rect 151078 53088 151084 53100
rect 13320 53060 151084 53088
rect 13320 53048 13326 53060
rect 151078 53048 151084 53060
rect 151136 53048 151142 53100
rect 151538 53048 151544 53100
rect 151596 53088 151602 53100
rect 577498 53088 577504 53100
rect 151596 53060 577504 53088
rect 151596 53048 151602 53060
rect 577498 53048 577504 53060
rect 577556 53048 577562 53100
rect 4982 51008 4988 51060
rect 5040 51048 5046 51060
rect 150434 51048 150440 51060
rect 5040 51020 150440 51048
rect 5040 51008 5046 51020
rect 150434 51008 150440 51020
rect 150492 51008 150498 51060
rect 6362 49648 6368 49700
rect 6420 49688 6426 49700
rect 150434 49688 150440 49700
rect 6420 49660 150440 49688
rect 6420 49648 6426 49660
rect 150434 49648 150440 49660
rect 150492 49648 150498 49700
rect 4890 48220 4896 48272
rect 4948 48260 4954 48272
rect 150434 48260 150440 48272
rect 4948 48232 150440 48260
rect 4948 48220 4954 48232
rect 150434 48220 150440 48232
rect 150492 48220 150498 48272
rect 21358 48152 21364 48204
rect 21416 48192 21422 48204
rect 150526 48192 150532 48204
rect 21416 48164 150532 48192
rect 21416 48152 21422 48164
rect 150526 48152 150532 48164
rect 150584 48152 150590 48204
rect 4798 46860 4804 46912
rect 4856 46900 4862 46912
rect 150434 46900 150440 46912
rect 4856 46872 150440 46900
rect 4856 46860 4862 46872
rect 150434 46860 150440 46872
rect 150492 46860 150498 46912
rect 13078 45500 13084 45552
rect 13136 45540 13142 45552
rect 150434 45540 150440 45552
rect 13136 45512 150440 45540
rect 13136 45500 13142 45512
rect 150434 45500 150440 45512
rect 150492 45500 150498 45552
rect 10318 44072 10324 44124
rect 10376 44112 10382 44124
rect 150434 44112 150440 44124
rect 10376 44084 150440 44112
rect 10376 44072 10382 44084
rect 150434 44072 150440 44084
rect 150492 44072 150498 44124
rect 8938 42712 8944 42764
rect 8996 42752 9002 42764
rect 150434 42752 150440 42764
rect 8996 42724 150440 42752
rect 8996 42712 9002 42724
rect 150434 42712 150440 42724
rect 150492 42712 150498 42764
rect 6270 41352 6276 41404
rect 6328 41392 6334 41404
rect 150434 41392 150440 41404
rect 6328 41364 150440 41392
rect 6328 41352 6334 41364
rect 150434 41352 150440 41364
rect 150492 41352 150498 41404
rect 7558 39312 7564 39364
rect 7616 39352 7622 39364
rect 151170 39352 151176 39364
rect 7616 39324 151176 39352
rect 7616 39312 7622 39324
rect 151170 39312 151176 39324
rect 151228 39312 151234 39364
rect 437382 37272 437388 37324
rect 437440 37312 437446 37324
rect 565078 37312 565084 37324
rect 437440 37284 565084 37312
rect 437440 37272 437446 37284
rect 565078 37272 565084 37284
rect 565136 37272 565142 37324
rect 9030 36524 9036 36576
rect 9088 36564 9094 36576
rect 151078 36564 151084 36576
rect 9088 36536 151084 36564
rect 9088 36524 9094 36536
rect 151078 36524 151084 36536
rect 151136 36524 151142 36576
rect 16482 35844 16488 35896
rect 16540 35884 16546 35896
rect 150434 35884 150440 35896
rect 16540 35856 150440 35884
rect 16540 35844 16546 35856
rect 150434 35844 150440 35856
rect 150492 35844 150498 35896
rect 15838 34416 15844 34468
rect 15896 34456 15902 34468
rect 150434 34456 150440 34468
rect 15896 34428 150440 34456
rect 15896 34416 15902 34428
rect 150434 34416 150440 34428
rect 150492 34416 150498 34468
rect 7650 33056 7656 33108
rect 7708 33096 7714 33108
rect 150434 33096 150440 33108
rect 7708 33068 150440 33096
rect 7708 33056 7714 33068
rect 150434 33056 150440 33068
rect 150492 33056 150498 33108
rect 3510 31696 3516 31748
rect 3568 31736 3574 31748
rect 150434 31736 150440 31748
rect 3568 31708 150440 31736
rect 3568 31696 3574 31708
rect 150434 31696 150440 31708
rect 150492 31696 150498 31748
rect 3418 30268 3424 30320
rect 3476 30308 3482 30320
rect 150434 30308 150440 30320
rect 3476 30280 150440 30308
rect 3476 30268 3482 30280
rect 150434 30268 150440 30280
rect 150492 30268 150498 30320
rect 5074 28908 5080 28960
rect 5132 28948 5138 28960
rect 150434 28948 150440 28960
rect 5132 28920 150440 28948
rect 5132 28908 5138 28920
rect 150434 28908 150440 28920
rect 150492 28908 150498 28960
rect 3602 26188 3608 26240
rect 3660 26228 3666 26240
rect 150434 26228 150440 26240
rect 3660 26200 150440 26228
rect 3660 26188 3666 26200
rect 150434 26188 150440 26200
rect 150492 26188 150498 26240
rect 214834 23740 214840 23792
rect 214892 23780 214898 23792
rect 299658 23780 299664 23792
rect 214892 23752 299664 23780
rect 214892 23740 214898 23752
rect 299658 23740 299664 23752
rect 299716 23740 299722 23792
rect 244090 23672 244096 23724
rect 244148 23712 244154 23724
rect 335998 23712 336004 23724
rect 244148 23684 336004 23712
rect 244148 23672 244154 23684
rect 335998 23672 336004 23684
rect 336056 23672 336062 23724
rect 266262 23604 266268 23656
rect 266320 23644 266326 23656
rect 480254 23644 480260 23656
rect 266320 23616 480260 23644
rect 266320 23604 266326 23616
rect 480254 23604 480260 23616
rect 480312 23604 480318 23656
rect 267366 23536 267372 23588
rect 267424 23576 267430 23588
rect 483014 23576 483020 23588
rect 267424 23548 483020 23576
rect 267424 23536 267430 23548
rect 483014 23536 483020 23548
rect 483072 23536 483078 23588
rect 269482 23468 269488 23520
rect 269540 23508 269546 23520
rect 489914 23508 489920 23520
rect 269540 23480 489920 23508
rect 269540 23468 269546 23480
rect 489914 23468 489920 23480
rect 489972 23468 489978 23520
rect 215478 22448 215484 22500
rect 215536 22488 215542 22500
rect 301406 22488 301412 22500
rect 215536 22460 301412 22488
rect 215536 22448 215542 22460
rect 301406 22448 301412 22460
rect 301464 22448 301470 22500
rect 217502 22380 217508 22432
rect 217560 22420 217566 22432
rect 309226 22420 309232 22432
rect 217560 22392 309232 22420
rect 217560 22380 217566 22392
rect 309226 22380 309232 22392
rect 309284 22380 309290 22432
rect 220538 22312 220544 22364
rect 220596 22352 220602 22364
rect 320266 22352 320272 22364
rect 220596 22324 320272 22352
rect 220596 22312 220602 22324
rect 320266 22312 320272 22324
rect 320324 22312 320330 22364
rect 228634 22244 228640 22296
rect 228692 22284 228698 22296
rect 349246 22284 349252 22296
rect 228692 22256 349252 22284
rect 228692 22244 228698 22256
rect 349246 22244 349252 22256
rect 349304 22244 349310 22296
rect 241790 22176 241796 22228
rect 241848 22216 241854 22228
rect 394694 22216 394700 22228
rect 241848 22188 394700 22216
rect 241848 22176 241854 22188
rect 394694 22176 394700 22188
rect 394752 22176 394758 22228
rect 275186 22108 275192 22160
rect 275244 22148 275250 22160
rect 511994 22148 512000 22160
rect 275244 22120 512000 22148
rect 275244 22108 275250 22120
rect 511994 22108 512000 22120
rect 512052 22108 512058 22160
rect 297358 21836 297364 21888
rect 297416 21876 297422 21888
rect 297416 21848 306374 21876
rect 297416 21836 297422 21848
rect 291838 21768 291844 21820
rect 291896 21808 291902 21820
rect 291896 21780 301544 21808
rect 291896 21768 291902 21780
rect 250898 21700 250904 21752
rect 250956 21740 250962 21752
rect 276014 21740 276020 21752
rect 250956 21712 276020 21740
rect 250956 21700 250962 21712
rect 276014 21700 276020 21712
rect 276072 21700 276078 21752
rect 278682 21700 278688 21752
rect 278740 21740 278746 21752
rect 297450 21740 297456 21752
rect 278740 21712 297456 21740
rect 278740 21700 278746 21712
rect 297450 21700 297456 21712
rect 297508 21700 297514 21752
rect 226610 21632 226616 21684
rect 226668 21672 226674 21684
rect 246298 21672 246304 21684
rect 226668 21644 246304 21672
rect 226668 21632 226674 21644
rect 246298 21632 246304 21644
rect 246356 21632 246362 21684
rect 254026 21632 254032 21684
rect 254084 21672 254090 21684
rect 301516 21672 301544 21780
rect 306346 21740 306374 21848
rect 383470 21768 383476 21820
rect 383528 21808 383534 21820
rect 388438 21808 388444 21820
rect 383528 21780 388444 21808
rect 383528 21768 383534 21780
rect 388438 21768 388444 21780
rect 388496 21768 388502 21820
rect 307570 21740 307576 21752
rect 306346 21712 307576 21740
rect 307570 21700 307576 21712
rect 307628 21700 307634 21752
rect 315298 21700 315304 21752
rect 315356 21740 315362 21752
rect 322750 21740 322756 21752
rect 315356 21712 322756 21740
rect 315356 21700 315362 21712
rect 322750 21700 322756 21712
rect 322808 21700 322814 21752
rect 350626 21700 350632 21752
rect 350684 21740 350690 21752
rect 358170 21740 358176 21752
rect 350684 21712 358176 21740
rect 350684 21700 350690 21712
rect 358170 21700 358176 21712
rect 358228 21700 358234 21752
rect 385494 21700 385500 21752
rect 385552 21740 385558 21752
rect 394602 21740 394608 21752
rect 385552 21712 394608 21740
rect 385552 21700 385558 21712
rect 394602 21700 394608 21712
rect 394660 21700 394666 21752
rect 398650 21700 398656 21752
rect 398708 21740 398714 21752
rect 437566 21740 437572 21752
rect 398708 21712 437572 21740
rect 398708 21700 398714 21712
rect 437566 21700 437572 21712
rect 437624 21700 437630 21752
rect 254084 21644 277394 21672
rect 301516 21644 306374 21672
rect 254084 21632 254090 21644
rect 230658 21564 230664 21616
rect 230716 21604 230722 21616
rect 262858 21604 262864 21616
rect 230716 21576 262864 21604
rect 230716 21564 230722 21576
rect 262858 21564 262864 21576
rect 262916 21564 262922 21616
rect 277366 21604 277394 21644
rect 298462 21604 298468 21616
rect 277366 21576 298468 21604
rect 298462 21564 298468 21576
rect 298520 21564 298526 21616
rect 306346 21604 306374 21644
rect 323578 21632 323584 21684
rect 323636 21672 323642 21684
rect 342990 21672 342996 21684
rect 323636 21644 342996 21672
rect 323636 21632 323642 21644
rect 342990 21632 342996 21644
rect 343048 21632 343054 21684
rect 369302 21632 369308 21684
rect 369360 21672 369366 21684
rect 371142 21672 371148 21684
rect 369360 21644 371148 21672
rect 369360 21632 369366 21644
rect 371142 21632 371148 21644
rect 371200 21632 371206 21684
rect 386506 21632 386512 21684
rect 386564 21672 386570 21684
rect 426802 21672 426808 21684
rect 386564 21644 426808 21672
rect 386564 21632 386570 21644
rect 426802 21632 426808 21644
rect 426860 21632 426866 21684
rect 338942 21604 338948 21616
rect 306346 21576 338948 21604
rect 338942 21564 338948 21576
rect 339000 21564 339006 21616
rect 342898 21564 342904 21616
rect 342956 21604 342962 21616
rect 354122 21604 354128 21616
rect 342956 21576 354128 21604
rect 342956 21564 342962 21576
rect 354122 21564 354128 21576
rect 354180 21564 354186 21616
rect 388530 21564 388536 21616
rect 388588 21604 388594 21616
rect 440234 21604 440240 21616
rect 388588 21576 440240 21604
rect 388588 21564 388594 21576
rect 440234 21564 440240 21576
rect 440292 21564 440298 21616
rect 164326 21496 164332 21548
rect 164384 21536 164390 21548
rect 176010 21536 176016 21548
rect 164384 21508 176016 21536
rect 164384 21496 164390 21508
rect 176010 21496 176016 21508
rect 176068 21496 176074 21548
rect 193214 21496 193220 21548
rect 193272 21536 193278 21548
rect 210326 21536 210332 21548
rect 193272 21508 210332 21536
rect 193272 21496 193278 21508
rect 210326 21496 210332 21508
rect 210384 21496 210390 21548
rect 211430 21496 211436 21548
rect 211488 21536 211494 21548
rect 249978 21536 249984 21548
rect 211488 21508 249984 21536
rect 211488 21496 211494 21508
rect 249978 21496 249984 21508
rect 250036 21496 250042 21548
rect 263042 21496 263048 21548
rect 263100 21536 263106 21548
rect 278130 21536 278136 21548
rect 263100 21508 278136 21536
rect 263100 21496 263106 21508
rect 278130 21496 278136 21508
rect 278188 21496 278194 21548
rect 279418 21496 279424 21548
rect 279476 21536 279482 21548
rect 279476 21508 318794 21536
rect 279476 21496 279482 21508
rect 199286 21428 199292 21480
rect 199344 21468 199350 21480
rect 228358 21468 228364 21480
rect 199344 21440 228364 21468
rect 199344 21428 199350 21440
rect 228358 21428 228364 21440
rect 228416 21428 228422 21480
rect 242158 21428 242164 21480
rect 242216 21468 242222 21480
rect 301498 21468 301504 21480
rect 242216 21440 301504 21468
rect 242216 21428 242222 21440
rect 301498 21428 301504 21440
rect 301556 21428 301562 21480
rect 304258 21428 304264 21480
rect 304316 21468 304322 21480
rect 312630 21468 312636 21480
rect 304316 21440 312636 21468
rect 304316 21428 304322 21440
rect 312630 21428 312636 21440
rect 312688 21428 312694 21480
rect 127618 21360 127624 21412
rect 127676 21400 127682 21412
rect 164878 21400 164884 21412
rect 127676 21372 164884 21400
rect 127676 21360 127682 21372
rect 164878 21360 164884 21372
rect 164936 21360 164942 21412
rect 206278 21360 206284 21412
rect 206336 21400 206342 21412
rect 303522 21400 303528 21412
rect 206336 21372 303528 21400
rect 206336 21360 206342 21372
rect 303522 21360 303528 21372
rect 303580 21360 303586 21412
rect 311618 21400 311624 21412
rect 306346 21372 311624 21400
rect 302878 21292 302884 21344
rect 302936 21332 302942 21344
rect 306346 21332 306374 21372
rect 311618 21360 311624 21372
rect 311676 21360 311682 21412
rect 302936 21304 306374 21332
rect 302936 21292 302942 21304
rect 311158 21292 311164 21344
rect 311216 21332 311222 21344
rect 316678 21332 316684 21344
rect 311216 21304 316684 21332
rect 311216 21292 311222 21304
rect 316678 21292 316684 21304
rect 316736 21292 316742 21344
rect 318766 21332 318794 21508
rect 320818 21496 320824 21548
rect 320876 21536 320882 21548
rect 320876 21508 328454 21536
rect 320876 21496 320882 21508
rect 328426 21468 328454 21508
rect 333974 21496 333980 21548
rect 334032 21536 334038 21548
rect 340966 21536 340972 21548
rect 334032 21508 340972 21536
rect 334032 21496 334038 21508
rect 340966 21496 340972 21508
rect 341024 21496 341030 21548
rect 343634 21496 343640 21548
rect 343692 21536 343698 21548
rect 356146 21536 356152 21548
rect 343692 21508 356152 21536
rect 343692 21496 343698 21508
rect 356146 21496 356152 21508
rect 356204 21496 356210 21548
rect 371326 21496 371332 21548
rect 371384 21536 371390 21548
rect 377490 21536 377496 21548
rect 371384 21508 377496 21536
rect 371384 21496 371390 21508
rect 377490 21496 377496 21508
rect 377548 21496 377554 21548
rect 381446 21496 381452 21548
rect 381504 21536 381510 21548
rect 387058 21536 387064 21548
rect 381504 21508 387064 21536
rect 381504 21496 381510 21508
rect 387058 21496 387064 21508
rect 387116 21496 387122 21548
rect 392578 21496 392584 21548
rect 392636 21536 392642 21548
rect 456886 21536 456892 21548
rect 392636 21508 456892 21536
rect 392636 21496 392642 21508
rect 456886 21496 456892 21508
rect 456944 21496 456950 21548
rect 345014 21468 345020 21480
rect 328426 21440 345020 21468
rect 345014 21428 345020 21440
rect 345072 21428 345078 21480
rect 390554 21428 390560 21480
rect 390612 21468 390618 21480
rect 465074 21468 465080 21480
rect 390612 21440 465080 21468
rect 390612 21428 390618 21440
rect 465074 21428 465080 21440
rect 465132 21428 465138 21480
rect 334894 21400 334900 21412
rect 321756 21372 334900 21400
rect 321756 21332 321784 21372
rect 334894 21360 334900 21372
rect 334952 21360 334958 21412
rect 351086 21400 351092 21412
rect 335326 21372 351092 21400
rect 318766 21304 321784 21332
rect 325694 21292 325700 21344
rect 325752 21332 325758 21344
rect 335326 21332 335354 21372
rect 351086 21360 351092 21372
rect 351144 21360 351150 21412
rect 368290 21360 368296 21412
rect 368348 21400 368354 21412
rect 378778 21400 378784 21412
rect 368348 21372 378784 21400
rect 368348 21360 368354 21372
rect 378778 21360 378784 21372
rect 378836 21360 378842 21412
rect 394510 21360 394516 21412
rect 394568 21400 394574 21412
rect 478874 21400 478880 21412
rect 394568 21372 478880 21400
rect 394568 21360 394574 21372
rect 478874 21360 478880 21372
rect 478932 21360 478938 21412
rect 325752 21304 335354 21332
rect 325752 21292 325758 21304
rect 312538 21224 312544 21276
rect 312596 21264 312602 21276
rect 319714 21264 319720 21276
rect 312596 21236 319720 21264
rect 312596 21224 312602 21236
rect 319714 21224 319720 21236
rect 319772 21224 319778 21276
rect 309778 21156 309784 21208
rect 309836 21196 309842 21208
rect 318702 21196 318708 21208
rect 309836 21168 318708 21196
rect 309836 21156 309842 21168
rect 318702 21156 318708 21168
rect 318760 21156 318766 21208
rect 322750 21156 322756 21208
rect 322808 21196 322814 21208
rect 325786 21196 325792 21208
rect 322808 21168 325792 21196
rect 322808 21156 322814 21168
rect 325786 21156 325792 21168
rect 325844 21156 325850 21208
rect 300946 21088 300952 21140
rect 301004 21128 301010 21140
rect 306558 21128 306564 21140
rect 301004 21100 306564 21128
rect 301004 21088 301010 21100
rect 306558 21088 306564 21100
rect 306616 21088 306622 21140
rect 375374 21020 375380 21072
rect 375432 21060 375438 21072
rect 382918 21060 382924 21072
rect 375432 21032 382924 21060
rect 375432 21020 375438 21032
rect 382918 21020 382924 21032
rect 382976 21020 382982 21072
rect 306558 20952 306564 21004
rect 306616 20992 306622 21004
rect 308582 20992 308588 21004
rect 306616 20964 308588 20992
rect 306616 20952 306622 20964
rect 308582 20952 308588 20964
rect 308640 20952 308646 21004
rect 347774 20952 347780 21004
rect 347832 20992 347838 21004
rect 357158 20992 357164 21004
rect 347832 20964 357164 20992
rect 347832 20952 347838 20964
rect 357158 20952 357164 20964
rect 357216 20952 357222 21004
rect 363230 20952 363236 21004
rect 363288 20992 363294 21004
rect 366358 20992 366364 21004
rect 363288 20964 366364 20992
rect 363288 20952 363294 20964
rect 366358 20952 366364 20964
rect 366416 20952 366422 21004
rect 174538 20884 174544 20936
rect 174596 20924 174602 20936
rect 178034 20924 178040 20936
rect 174596 20896 178040 20924
rect 174596 20884 174602 20896
rect 178034 20884 178040 20896
rect 178092 20884 178098 20936
rect 184106 20816 184112 20868
rect 184164 20856 184170 20868
rect 185578 20856 185584 20868
rect 184164 20828 185584 20856
rect 184164 20816 184170 20828
rect 185578 20816 185584 20828
rect 185636 20816 185642 20868
rect 234706 20816 234712 20868
rect 234764 20856 234770 20868
rect 240778 20856 240784 20868
rect 234764 20828 240784 20856
rect 234764 20816 234770 20828
rect 240778 20816 240784 20828
rect 240836 20816 240842 20868
rect 380434 20816 380440 20868
rect 380492 20856 380498 20868
rect 384390 20856 384396 20868
rect 380492 20828 384396 20856
rect 380492 20816 380498 20828
rect 384390 20816 384396 20828
rect 384448 20816 384454 20868
rect 178034 20748 178040 20800
rect 178092 20788 178098 20800
rect 180058 20788 180064 20800
rect 178092 20760 180064 20788
rect 178092 20748 178098 20760
rect 180058 20748 180064 20760
rect 180116 20748 180122 20800
rect 182082 20748 182088 20800
rect 182140 20788 182146 20800
rect 184198 20788 184204 20800
rect 182140 20760 184204 20788
rect 182140 20748 182146 20760
rect 184198 20748 184204 20760
rect 184256 20748 184262 20800
rect 317046 20748 317052 20800
rect 317104 20788 317110 20800
rect 323762 20788 323768 20800
rect 317104 20760 323768 20788
rect 317104 20748 317110 20760
rect 323762 20748 323768 20760
rect 323820 20748 323826 20800
rect 366266 20748 366272 20800
rect 366324 20788 366330 20800
rect 367738 20788 367744 20800
rect 366324 20760 367744 20788
rect 366324 20748 366330 20760
rect 367738 20748 367744 20760
rect 367796 20748 367802 20800
rect 171778 20680 171784 20732
rect 171836 20720 171842 20732
rect 177022 20720 177028 20732
rect 171836 20692 177028 20720
rect 171836 20680 171842 20692
rect 177022 20680 177028 20692
rect 177080 20680 177086 20732
rect 177298 20680 177304 20732
rect 177356 20720 177362 20732
rect 179046 20720 179052 20732
rect 177356 20692 179052 20720
rect 177356 20680 177362 20692
rect 179046 20680 179052 20692
rect 179104 20680 179110 20732
rect 181070 20680 181076 20732
rect 181128 20720 181134 20732
rect 182174 20720 182180 20732
rect 181128 20692 182180 20720
rect 181128 20680 181134 20692
rect 182174 20680 182180 20692
rect 182232 20680 182238 20732
rect 183094 20680 183100 20732
rect 183152 20720 183158 20732
rect 184290 20720 184296 20732
rect 183152 20692 184296 20720
rect 183152 20680 183158 20692
rect 184290 20680 184296 20692
rect 184348 20680 184354 20732
rect 210418 20680 210424 20732
rect 210476 20720 210482 20732
rect 211798 20720 211804 20732
rect 210476 20692 211804 20720
rect 210476 20680 210482 20692
rect 211798 20680 211804 20692
rect 211856 20680 211862 20732
rect 298738 20680 298744 20732
rect 298796 20720 298802 20732
rect 304534 20720 304540 20732
rect 298796 20692 304540 20720
rect 298796 20680 298802 20692
rect 304534 20680 304540 20692
rect 304592 20680 304598 20732
rect 307110 20680 307116 20732
rect 307168 20720 307174 20732
rect 309594 20720 309600 20732
rect 307168 20692 309600 20720
rect 307168 20680 307174 20692
rect 309594 20680 309600 20692
rect 309652 20680 309658 20732
rect 311250 20680 311256 20732
rect 311308 20720 311314 20732
rect 314654 20720 314660 20732
rect 311308 20692 314660 20720
rect 311308 20680 311314 20692
rect 314654 20680 314660 20692
rect 314712 20680 314718 20732
rect 318058 20680 318064 20732
rect 318116 20720 318122 20732
rect 320726 20720 320732 20732
rect 318116 20692 320732 20720
rect 318116 20680 318122 20692
rect 320726 20680 320732 20692
rect 320784 20680 320790 20732
rect 356698 20680 356704 20732
rect 356756 20720 356762 20732
rect 359182 20720 359188 20732
rect 356756 20692 359188 20720
rect 356756 20680 356762 20692
rect 359182 20680 359188 20692
rect 359240 20680 359246 20732
rect 359458 20680 359464 20732
rect 359516 20720 359522 20732
rect 360194 20720 360200 20732
rect 359516 20692 360200 20720
rect 359516 20680 359522 20692
rect 360194 20680 360200 20692
rect 360252 20680 360258 20732
rect 362218 20680 362224 20732
rect 362276 20720 362282 20732
rect 363598 20720 363604 20732
rect 362276 20692 363604 20720
rect 362276 20680 362282 20692
rect 363598 20680 363604 20692
rect 363656 20680 363662 20732
rect 365254 20680 365260 20732
rect 365312 20720 365318 20732
rect 366450 20720 366456 20732
rect 365312 20692 366456 20720
rect 365312 20680 365318 20692
rect 366450 20680 366456 20692
rect 366508 20680 366514 20732
rect 378410 20680 378416 20732
rect 378468 20720 378474 20732
rect 380158 20720 380164 20732
rect 378468 20692 380164 20720
rect 378468 20680 378474 20692
rect 380158 20680 380164 20692
rect 380216 20680 380222 20732
rect 384482 20680 384488 20732
rect 384540 20720 384546 20732
rect 392578 20720 392584 20732
rect 384540 20692 392584 20720
rect 384540 20680 384546 20692
rect 392578 20680 392584 20692
rect 392636 20680 392642 20732
rect 249978 20340 249984 20392
rect 250036 20380 250042 20392
rect 288434 20380 288440 20392
rect 250036 20352 288440 20380
rect 250036 20340 250042 20352
rect 288434 20340 288440 20352
rect 288492 20340 288498 20392
rect 301590 20340 301596 20392
rect 301648 20380 301654 20392
rect 331858 20380 331864 20392
rect 301648 20352 331864 20380
rect 301648 20340 301654 20352
rect 331858 20340 331864 20352
rect 331916 20340 331922 20392
rect 237374 20272 237380 20324
rect 237432 20312 237438 20324
rect 322750 20312 322756 20324
rect 237432 20284 322756 20312
rect 237432 20272 237438 20284
rect 322750 20272 322756 20284
rect 322808 20272 322814 20324
rect 201494 20204 201500 20256
rect 201552 20244 201558 20256
rect 315666 20244 315672 20256
rect 201552 20216 315672 20244
rect 201552 20204 201558 20216
rect 315666 20204 315672 20216
rect 315724 20204 315730 20256
rect 334618 20204 334624 20256
rect 334676 20244 334682 20256
rect 350074 20244 350080 20256
rect 334676 20216 350080 20244
rect 334676 20204 334682 20216
rect 350074 20204 350080 20216
rect 350132 20204 350138 20256
rect 394602 20204 394608 20256
rect 394660 20244 394666 20256
rect 447134 20244 447140 20256
rect 394660 20216 447140 20244
rect 394660 20204 394666 20216
rect 447134 20204 447140 20216
rect 447192 20204 447198 20256
rect 176654 20136 176660 20188
rect 176712 20176 176718 20188
rect 306558 20176 306564 20188
rect 176712 20148 306564 20176
rect 176712 20136 176718 20148
rect 306558 20136 306564 20148
rect 306616 20136 306622 20188
rect 330478 20136 330484 20188
rect 330536 20176 330542 20188
rect 347038 20176 347044 20188
rect 330536 20148 347044 20176
rect 330536 20136 330542 20148
rect 347038 20136 347044 20148
rect 347096 20136 347102 20188
rect 378778 20136 378784 20188
rect 378836 20176 378842 20188
rect 386414 20176 386420 20188
rect 378836 20148 386420 20176
rect 378836 20136 378842 20148
rect 386414 20136 386420 20148
rect 386472 20136 386478 20188
rect 396626 20136 396632 20188
rect 396684 20176 396690 20188
rect 485774 20176 485780 20188
rect 396684 20148 485780 20176
rect 396684 20136 396690 20148
rect 485774 20136 485780 20148
rect 485832 20136 485838 20188
rect 169754 20068 169760 20120
rect 169812 20108 169818 20120
rect 300946 20108 300952 20120
rect 169812 20080 300952 20108
rect 169812 20068 169818 20080
rect 300946 20068 300952 20080
rect 301004 20068 301010 20120
rect 319438 20068 319444 20120
rect 319496 20108 319502 20120
rect 339954 20108 339960 20120
rect 319496 20080 339960 20108
rect 319496 20068 319502 20080
rect 339954 20068 339960 20080
rect 340012 20068 340018 20120
rect 371142 20068 371148 20120
rect 371200 20108 371206 20120
rect 390738 20108 390744 20120
rect 371200 20080 390744 20108
rect 371200 20068 371206 20080
rect 390738 20068 390744 20080
rect 390796 20068 390802 20120
rect 397638 20068 397644 20120
rect 397696 20108 397702 20120
rect 490006 20108 490012 20120
rect 397696 20080 490012 20108
rect 397696 20068 397702 20080
rect 490006 20068 490012 20080
rect 490064 20068 490070 20120
rect 138014 20000 138020 20052
rect 138072 20040 138078 20052
rect 278682 20040 278688 20052
rect 138072 20012 278688 20040
rect 138072 20000 138078 20012
rect 278682 20000 278688 20012
rect 278740 20000 278746 20052
rect 291194 20000 291200 20052
rect 291252 20040 291258 20052
rect 333974 20040 333980 20052
rect 291252 20012 333980 20040
rect 291252 20000 291258 20012
rect 333974 20000 333980 20012
rect 334032 20000 334038 20052
rect 367278 20000 367284 20052
rect 367336 20040 367342 20052
rect 382274 20040 382280 20052
rect 367336 20012 382280 20040
rect 367336 20000 367342 20012
rect 382274 20000 382280 20012
rect 382332 20000 382338 20052
rect 382918 20000 382924 20052
rect 382976 20040 382982 20052
rect 411254 20040 411260 20052
rect 382976 20012 411260 20040
rect 382976 20000 382982 20012
rect 411254 20000 411260 20012
rect 411312 20000 411318 20052
rect 411806 20000 411812 20052
rect 411864 20040 411870 20052
rect 539594 20040 539600 20052
rect 411864 20012 539600 20040
rect 411864 20000 411870 20012
rect 539594 20000 539600 20012
rect 539652 20000 539658 20052
rect 165614 19932 165620 19984
rect 165672 19972 165678 19984
rect 166534 19972 166540 19984
rect 165672 19944 166540 19972
rect 165672 19932 165678 19944
rect 166534 19932 166540 19944
rect 166592 19932 166598 19984
rect 169846 19932 169852 19984
rect 169904 19972 169910 19984
rect 170582 19972 170588 19984
rect 169904 19944 170588 19972
rect 169904 19932 169910 19944
rect 170582 19932 170588 19944
rect 170640 19932 170646 19984
rect 173894 19932 173900 19984
rect 173952 19972 173958 19984
rect 174630 19972 174636 19984
rect 173952 19944 174636 19972
rect 173952 19932 173958 19944
rect 174630 19932 174636 19944
rect 174688 19932 174694 19984
rect 189074 19932 189080 19984
rect 189132 19972 189138 19984
rect 189902 19972 189908 19984
rect 189132 19944 189908 19972
rect 189132 19932 189138 19944
rect 189902 19932 189908 19944
rect 189960 19932 189966 19984
rect 195974 19932 195980 19984
rect 196032 19972 196038 19984
rect 196894 19972 196900 19984
rect 196032 19944 196900 19972
rect 196032 19932 196038 19944
rect 196894 19932 196900 19944
rect 196952 19932 196958 19984
rect 208394 19932 208400 19984
rect 208452 19972 208458 19984
rect 209038 19972 209044 19984
rect 208452 19944 209044 19972
rect 208452 19932 208458 19944
rect 209038 19932 209044 19944
rect 209096 19932 209102 19984
rect 245746 19932 245752 19984
rect 245804 19972 245810 19984
rect 246574 19972 246580 19984
rect 245804 19944 246580 19972
rect 245804 19932 245810 19944
rect 246574 19932 246580 19944
rect 246632 19932 246638 19984
rect 271874 19932 271880 19984
rect 271932 19972 271938 19984
rect 272886 19972 272892 19984
rect 271932 19944 272892 19972
rect 271932 19932 271938 19944
rect 272886 19932 272892 19944
rect 272944 19932 272950 19984
rect 278130 19932 278136 19984
rect 278188 19972 278194 19984
rect 469214 19972 469220 19984
rect 278188 19944 469220 19972
rect 278188 19932 278194 19944
rect 469214 19932 469220 19944
rect 469272 19932 469278 19984
rect 287054 19864 287060 19916
rect 287112 19904 287118 19916
rect 287974 19904 287980 19916
rect 287112 19876 287980 19904
rect 287112 19864 287118 19876
rect 287974 19864 287980 19876
rect 288032 19864 288038 19916
rect 332594 19864 332600 19916
rect 332652 19904 332658 19916
rect 333606 19904 333612 19916
rect 332652 19876 333612 19904
rect 332652 19864 332658 19876
rect 333606 19864 333612 19876
rect 333664 19864 333670 19916
rect 336734 19864 336740 19916
rect 336792 19904 336798 19916
rect 337654 19904 337660 19916
rect 336792 19876 337660 19904
rect 336792 19864 336798 19876
rect 337654 19864 337660 19876
rect 337712 19864 337718 19916
rect 401594 19864 401600 19916
rect 401652 19904 401658 19916
rect 402422 19904 402428 19916
rect 401652 19876 402428 19904
rect 401652 19864 401658 19876
rect 402422 19864 402428 19876
rect 402480 19864 402486 19916
rect 408586 19864 408592 19916
rect 408644 19904 408650 19916
rect 409414 19904 409420 19916
rect 408644 19876 409420 19904
rect 408644 19864 408650 19876
rect 409414 19864 409420 19876
rect 409472 19864 409478 19916
rect 412726 19864 412732 19916
rect 412784 19904 412790 19916
rect 413462 19904 413468 19916
rect 412784 19876 413468 19904
rect 412784 19864 412790 19876
rect 413462 19864 413468 19876
rect 413520 19864 413526 19916
rect 389542 19524 389548 19576
rect 389600 19564 389606 19576
rect 393958 19564 393964 19576
rect 389600 19536 393964 19564
rect 389600 19524 389606 19536
rect 393958 19524 393964 19536
rect 394016 19524 394022 19576
rect 185210 18912 185216 18964
rect 185268 18952 185274 18964
rect 310606 18952 310612 18964
rect 185268 18924 310612 18952
rect 185268 18912 185274 18924
rect 310606 18912 310612 18924
rect 310664 18912 310670 18964
rect 420914 18912 420920 18964
rect 420972 18952 420978 18964
rect 421558 18952 421564 18964
rect 420972 18924 421564 18952
rect 420972 18912 420978 18924
rect 421558 18912 421564 18924
rect 421616 18912 421622 18964
rect 135254 18844 135260 18896
rect 135312 18884 135318 18896
rect 296438 18884 296444 18896
rect 135312 18856 296444 18884
rect 135312 18844 135318 18856
rect 296438 18844 296444 18856
rect 296496 18844 296502 18896
rect 298094 18844 298100 18896
rect 298152 18884 298158 18896
rect 323578 18884 323584 18896
rect 298152 18856 323584 18884
rect 298152 18844 298158 18856
rect 323578 18844 323584 18856
rect 323636 18844 323642 18896
rect 257982 18776 257988 18828
rect 258040 18816 258046 18828
rect 451274 18816 451280 18828
rect 258040 18788 451280 18816
rect 258040 18776 258046 18788
rect 451274 18776 451280 18788
rect 451332 18776 451338 18828
rect 258994 18708 259000 18760
rect 259052 18748 259058 18760
rect 455414 18748 455420 18760
rect 259052 18720 455420 18748
rect 259052 18708 259058 18720
rect 455414 18708 455420 18720
rect 455472 18708 455478 18760
rect 202322 18640 202328 18692
rect 202380 18680 202386 18692
rect 256694 18680 256700 18692
rect 202380 18652 256700 18680
rect 202380 18640 202386 18652
rect 256694 18640 256700 18652
rect 256752 18640 256758 18692
rect 260006 18640 260012 18692
rect 260064 18680 260070 18692
rect 458174 18680 458180 18692
rect 260064 18652 458180 18680
rect 260064 18640 260070 18652
rect 458174 18640 458180 18652
rect 458232 18640 458238 18692
rect 203334 18572 203340 18624
rect 203392 18612 203398 18624
rect 259454 18612 259460 18624
rect 203392 18584 259460 18612
rect 203392 18572 203398 18584
rect 259454 18572 259460 18584
rect 259512 18572 259518 18624
rect 261018 18572 261024 18624
rect 261076 18612 261082 18624
rect 462314 18612 462320 18624
rect 261076 18584 462320 18612
rect 261076 18572 261082 18584
rect 462314 18572 462320 18584
rect 462372 18572 462378 18624
rect 230474 17552 230480 17604
rect 230532 17592 230538 17604
rect 317046 17592 317052 17604
rect 230532 17564 317052 17592
rect 230532 17552 230538 17564
rect 317046 17552 317052 17564
rect 317104 17552 317110 17604
rect 142154 17484 142160 17536
rect 142212 17524 142218 17536
rect 254026 17524 254032 17536
rect 142212 17496 254032 17524
rect 142212 17484 142218 17496
rect 254026 17484 254032 17496
rect 254084 17484 254090 17536
rect 276014 17484 276020 17536
rect 276072 17524 276078 17536
rect 426434 17524 426440 17536
rect 276072 17496 426440 17524
rect 276072 17484 276078 17496
rect 426434 17484 426440 17496
rect 426492 17484 426498 17536
rect 426802 17484 426808 17536
rect 426860 17524 426866 17536
rect 449894 17524 449900 17536
rect 426860 17496 449900 17524
rect 426860 17484 426866 17496
rect 449894 17484 449900 17496
rect 449952 17484 449958 17536
rect 131114 17416 131120 17468
rect 131172 17456 131178 17468
rect 295426 17456 295432 17468
rect 131172 17428 295432 17456
rect 131172 17416 131178 17428
rect 295426 17416 295432 17428
rect 295484 17416 295490 17468
rect 416866 17416 416872 17468
rect 416924 17456 416930 17468
rect 556154 17456 556160 17468
rect 416924 17428 556160 17456
rect 416924 17416 416930 17428
rect 556154 17416 556160 17428
rect 556212 17416 556218 17468
rect 251910 17348 251916 17400
rect 251968 17388 251974 17400
rect 430574 17388 430580 17400
rect 251968 17360 430580 17388
rect 251968 17348 251974 17360
rect 430574 17348 430580 17360
rect 430632 17348 430638 17400
rect 198274 17280 198280 17332
rect 198332 17320 198338 17332
rect 242894 17320 242900 17332
rect 198332 17292 242900 17320
rect 198332 17280 198338 17292
rect 242894 17280 242900 17292
rect 242952 17280 242958 17332
rect 252922 17280 252928 17332
rect 252980 17320 252986 17332
rect 433334 17320 433340 17332
rect 252980 17292 433340 17320
rect 252980 17280 252986 17292
rect 433334 17280 433340 17292
rect 433392 17280 433398 17332
rect 440234 17280 440240 17332
rect 440292 17320 440298 17332
rect 456794 17320 456800 17332
rect 440292 17292 456800 17320
rect 440292 17280 440298 17292
rect 456794 17280 456800 17292
rect 456852 17280 456858 17332
rect 456886 17280 456892 17332
rect 456944 17320 456950 17332
rect 471974 17320 471980 17332
rect 456944 17292 471980 17320
rect 456944 17280 456950 17292
rect 471974 17280 471980 17292
rect 472032 17280 472038 17332
rect 201310 17212 201316 17264
rect 201368 17252 201374 17264
rect 252554 17252 252560 17264
rect 201368 17224 252560 17252
rect 201368 17212 201374 17224
rect 252554 17212 252560 17224
rect 252612 17212 252618 17264
rect 253934 17212 253940 17264
rect 253992 17252 253998 17264
rect 437474 17252 437480 17264
rect 253992 17224 437480 17252
rect 253992 17212 253998 17224
rect 437474 17212 437480 17224
rect 437532 17212 437538 17264
rect 437566 17212 437572 17264
rect 437624 17252 437630 17264
rect 492674 17252 492680 17264
rect 437624 17224 492680 17252
rect 437624 17212 437630 17224
rect 492674 17212 492680 17224
rect 492732 17212 492738 17264
rect 204254 16668 204260 16720
rect 204312 16708 204318 16720
rect 204990 16708 204996 16720
rect 204312 16680 204996 16708
rect 204312 16668 204318 16680
rect 204990 16668 204996 16680
rect 205048 16668 205054 16720
rect 145466 16192 145472 16244
rect 145524 16232 145530 16244
rect 247678 16232 247684 16244
rect 145524 16204 247684 16232
rect 145524 16192 145530 16204
rect 247678 16192 247684 16204
rect 247736 16192 247742 16244
rect 273898 16192 273904 16244
rect 273956 16232 273962 16244
rect 304994 16232 305000 16244
rect 273956 16204 305000 16232
rect 273956 16192 273962 16204
rect 304994 16192 305000 16204
rect 305052 16192 305058 16244
rect 307018 16192 307024 16244
rect 307076 16232 307082 16244
rect 329926 16232 329932 16244
rect 307076 16204 329932 16232
rect 307076 16192 307082 16204
rect 329926 16192 329932 16204
rect 329984 16192 329990 16244
rect 401686 16192 401692 16244
rect 401744 16232 401750 16244
rect 503714 16232 503720 16244
rect 401744 16204 503720 16232
rect 401744 16192 401750 16204
rect 503714 16192 503720 16204
rect 503772 16192 503778 16244
rect 198734 16124 198740 16176
rect 198792 16164 198798 16176
rect 311250 16164 311256 16176
rect 198792 16136 311256 16164
rect 198792 16124 198798 16136
rect 311250 16124 311256 16136
rect 311308 16124 311314 16176
rect 402974 16124 402980 16176
rect 403032 16164 403038 16176
rect 511258 16164 511264 16176
rect 403032 16136 511264 16164
rect 403032 16124 403038 16136
rect 511258 16124 511264 16136
rect 511316 16124 511322 16176
rect 244274 16056 244280 16108
rect 244332 16096 244338 16108
rect 406010 16096 406016 16108
rect 244332 16068 406016 16096
rect 244332 16056 244338 16068
rect 406010 16056 406016 16068
rect 406068 16056 406074 16108
rect 409138 16096 409144 16108
rect 406120 16068 409144 16096
rect 228358 15988 228364 16040
rect 228416 16028 228422 16040
rect 228416 16000 245056 16028
rect 228416 15988 228422 16000
rect 196066 15920 196072 15972
rect 196124 15960 196130 15972
rect 234614 15960 234620 15972
rect 196124 15932 234620 15960
rect 196124 15920 196130 15932
rect 234614 15920 234620 15932
rect 234672 15920 234678 15972
rect 200114 15852 200120 15904
rect 200172 15892 200178 15904
rect 244918 15892 244924 15904
rect 200172 15864 244924 15892
rect 200172 15852 200178 15864
rect 244918 15852 244924 15864
rect 244976 15852 244982 15904
rect 245028 15892 245056 16000
rect 245838 15988 245844 16040
rect 245896 16028 245902 16040
rect 406120 16028 406148 16068
rect 409138 16056 409144 16068
rect 409196 16056 409202 16108
rect 245896 16000 406148 16028
rect 245896 15988 245902 16000
rect 408678 15988 408684 16040
rect 408736 16028 408742 16040
rect 528554 16028 528560 16040
rect 408736 16000 528560 16028
rect 408736 15988 408742 16000
rect 528554 15988 528560 16000
rect 528612 15988 528618 16040
rect 245746 15920 245752 15972
rect 245804 15960 245810 15972
rect 412634 15960 412640 15972
rect 245804 15932 412640 15960
rect 245804 15920 245810 15932
rect 412634 15920 412640 15932
rect 412692 15920 412698 15972
rect 412818 15920 412824 15972
rect 412876 15960 412882 15972
rect 542722 15960 542728 15972
rect 412876 15932 542728 15960
rect 412876 15920 412882 15932
rect 542722 15920 542728 15932
rect 542780 15920 542786 15972
rect 245930 15892 245936 15904
rect 245028 15864 245936 15892
rect 245930 15852 245936 15864
rect 245988 15852 245994 15904
rect 247034 15852 247040 15904
rect 247092 15892 247098 15904
rect 415394 15892 415400 15904
rect 247092 15864 415400 15892
rect 247092 15852 247098 15864
rect 415394 15852 415400 15864
rect 415452 15852 415458 15904
rect 260098 14764 260104 14816
rect 260156 14804 260162 14816
rect 330386 14804 330392 14816
rect 260156 14776 330392 14804
rect 260156 14764 260162 14776
rect 330386 14764 330392 14776
rect 330444 14764 330450 14816
rect 380158 14764 380164 14816
rect 380216 14804 380222 14816
rect 422570 14804 422576 14816
rect 380216 14776 422576 14804
rect 380216 14764 380222 14776
rect 422570 14764 422576 14776
rect 422628 14764 422634 14816
rect 213362 14696 213368 14748
rect 213420 14736 213426 14748
rect 309778 14736 309784 14748
rect 213420 14708 309784 14736
rect 213420 14696 213426 14708
rect 309778 14696 309784 14708
rect 309836 14696 309842 14748
rect 384390 14696 384396 14748
rect 384448 14736 384454 14748
rect 429194 14736 429200 14748
rect 384448 14708 429200 14736
rect 384448 14696 384454 14708
rect 429194 14696 429200 14708
rect 429252 14696 429258 14748
rect 235994 14628 236000 14680
rect 236052 14668 236058 14680
rect 347038 14668 347044 14680
rect 236052 14640 347044 14668
rect 236052 14628 236058 14640
rect 347038 14628 347044 14640
rect 347096 14628 347102 14680
rect 388438 14628 388444 14680
rect 388496 14668 388502 14680
rect 440326 14668 440332 14680
rect 388496 14640 440332 14668
rect 388496 14628 388502 14640
rect 440326 14628 440332 14640
rect 440384 14628 440390 14680
rect 190454 14560 190460 14612
rect 190512 14600 190518 14612
rect 218054 14600 218060 14612
rect 190512 14572 218060 14600
rect 190512 14560 190518 14572
rect 218054 14560 218060 14572
rect 218112 14560 218118 14612
rect 237466 14560 237472 14612
rect 237524 14600 237530 14612
rect 370498 14600 370504 14612
rect 237524 14572 370504 14600
rect 237524 14560 237530 14572
rect 370498 14560 370504 14572
rect 370556 14560 370562 14612
rect 376754 14560 376760 14612
rect 376812 14600 376818 14612
rect 418522 14600 418528 14612
rect 376812 14572 418528 14600
rect 376812 14560 376818 14572
rect 418522 14560 418528 14572
rect 418580 14560 418586 14612
rect 419534 14560 419540 14612
rect 419592 14600 419598 14612
rect 567562 14600 567568 14612
rect 419592 14572 567568 14600
rect 419592 14560 419598 14572
rect 567562 14560 567568 14572
rect 567620 14560 567626 14612
rect 194594 14492 194600 14544
rect 194652 14532 194658 14544
rect 231854 14532 231860 14544
rect 194652 14504 231860 14532
rect 194652 14492 194658 14504
rect 231854 14492 231860 14504
rect 231912 14492 231918 14544
rect 238846 14492 238852 14544
rect 238904 14532 238910 14544
rect 377398 14532 377404 14544
rect 238904 14504 377404 14532
rect 238904 14492 238910 14504
rect 377398 14492 377404 14504
rect 377456 14492 377462 14544
rect 421006 14492 421012 14544
rect 421064 14532 421070 14544
rect 571334 14532 571340 14544
rect 421064 14504 571340 14532
rect 421064 14492 421070 14504
rect 571334 14492 571340 14504
rect 571392 14492 571398 14544
rect 195974 14424 195980 14476
rect 196032 14464 196038 14476
rect 196032 14436 238754 14464
rect 196032 14424 196038 14436
rect 238726 14396 238754 14436
rect 238938 14424 238944 14476
rect 238996 14464 239002 14476
rect 381538 14464 381544 14476
rect 238996 14436 381544 14464
rect 238996 14424 239002 14436
rect 381538 14424 381544 14436
rect 381596 14424 381602 14476
rect 420914 14424 420920 14476
rect 420972 14464 420978 14476
rect 575106 14464 575112 14476
rect 420972 14436 575112 14464
rect 420972 14424 420978 14436
rect 575106 14424 575112 14436
rect 575164 14424 575170 14476
rect 239306 14396 239312 14408
rect 238726 14368 239312 14396
rect 239306 14356 239312 14368
rect 239364 14356 239370 14408
rect 262858 13404 262864 13456
rect 262916 13444 262922 13456
rect 356330 13444 356336 13456
rect 262916 13416 356336 13444
rect 262916 13404 262922 13416
rect 356330 13404 356336 13416
rect 356388 13404 356394 13456
rect 219986 13336 219992 13388
rect 220044 13376 220050 13388
rect 318058 13376 318064 13388
rect 220044 13348 318064 13376
rect 220044 13336 220050 13348
rect 318058 13336 318064 13348
rect 318116 13336 318122 13388
rect 378686 13336 378692 13388
rect 378744 13376 378750 13388
rect 425698 13376 425704 13388
rect 378744 13348 425704 13376
rect 378744 13336 378750 13348
rect 425698 13336 425704 13348
rect 425756 13336 425762 13388
rect 229094 13268 229100 13320
rect 229152 13308 229158 13320
rect 337378 13308 337384 13320
rect 229152 13280 337384 13308
rect 229152 13268 229158 13280
rect 337378 13268 337384 13280
rect 337436 13268 337442 13320
rect 381722 13268 381728 13320
rect 381780 13308 381786 13320
rect 515490 13308 515496 13320
rect 381780 13280 515496 13308
rect 381780 13268 381786 13280
rect 515490 13268 515496 13280
rect 515548 13268 515554 13320
rect 230842 13200 230848 13252
rect 230900 13240 230906 13252
rect 359366 13240 359372 13252
rect 230900 13212 359372 13240
rect 230900 13200 230906 13212
rect 359366 13200 359372 13212
rect 359424 13200 359430 13252
rect 375466 13200 375472 13252
rect 375524 13240 375530 13252
rect 375524 13212 383654 13240
rect 375524 13200 375530 13212
rect 231946 13132 231952 13184
rect 232004 13172 232010 13184
rect 363414 13172 363420 13184
rect 232004 13144 363420 13172
rect 232004 13132 232010 13144
rect 363414 13132 363420 13144
rect 363472 13132 363478 13184
rect 369854 13132 369860 13184
rect 369912 13172 369918 13184
rect 381630 13172 381636 13184
rect 369912 13144 381636 13172
rect 369912 13132 369918 13144
rect 381630 13132 381636 13144
rect 381688 13132 381694 13184
rect 193306 13064 193312 13116
rect 193364 13104 193370 13116
rect 228266 13104 228272 13116
rect 193364 13076 228272 13104
rect 193364 13064 193370 13076
rect 228266 13064 228272 13076
rect 228324 13064 228330 13116
rect 233234 13064 233240 13116
rect 233292 13104 233298 13116
rect 365806 13104 365812 13116
rect 233292 13076 365812 13104
rect 233292 13064 233298 13076
rect 365806 13064 365812 13076
rect 365864 13064 365870 13116
rect 366450 13064 366456 13116
rect 366508 13104 366514 13116
rect 376018 13104 376024 13116
rect 366508 13076 376024 13104
rect 366508 13064 366514 13076
rect 376018 13064 376024 13076
rect 376076 13064 376082 13116
rect 383626 13104 383654 13212
rect 412726 13200 412732 13252
rect 412784 13240 412790 13252
rect 546494 13240 546500 13252
rect 412784 13212 546500 13240
rect 412784 13200 412790 13212
rect 546494 13200 546500 13212
rect 546552 13200 546558 13252
rect 386690 13132 386696 13184
rect 386748 13172 386754 13184
rect 413278 13172 413284 13184
rect 386748 13144 413284 13172
rect 386748 13132 386754 13144
rect 413278 13132 413284 13144
rect 413336 13132 413342 13184
rect 414014 13132 414020 13184
rect 414072 13172 414078 13184
rect 550266 13172 550272 13184
rect 414072 13144 550272 13172
rect 414072 13132 414078 13144
rect 550266 13132 550272 13144
rect 550324 13132 550330 13184
rect 415486 13104 415492 13116
rect 383626 13076 415492 13104
rect 415486 13064 415492 13076
rect 415544 13064 415550 13116
rect 415578 13064 415584 13116
rect 415636 13104 415642 13116
rect 553762 13104 553768 13116
rect 415636 13076 553768 13104
rect 415636 13064 415642 13076
rect 553762 13064 553768 13076
rect 553820 13064 553826 13116
rect 276658 12044 276664 12096
rect 276716 12084 276722 12096
rect 336826 12084 336832 12096
rect 276716 12056 336832 12084
rect 276716 12044 276722 12056
rect 336826 12044 336832 12056
rect 336884 12044 336890 12096
rect 210326 11976 210332 12028
rect 210384 12016 210390 12028
rect 225138 12016 225144 12028
rect 210384 11988 225144 12016
rect 210384 11976 210390 11988
rect 225138 11976 225144 11988
rect 225196 11976 225202 12028
rect 227530 11976 227536 12028
rect 227588 12016 227594 12028
rect 315298 12016 315304 12028
rect 227588 11988 315304 12016
rect 227588 11976 227594 11988
rect 315298 11976 315304 11988
rect 315356 11976 315362 12028
rect 387058 11976 387064 12028
rect 387116 12016 387122 12028
rect 431954 12016 431960 12028
rect 387116 11988 431960 12016
rect 387116 11976 387122 11988
rect 431954 11976 431960 11988
rect 432012 11976 432018 12028
rect 151814 11908 151820 11960
rect 151872 11948 151878 11960
rect 242158 11948 242164 11960
rect 151872 11920 242164 11948
rect 151872 11908 151878 11920
rect 242158 11908 242164 11920
rect 242216 11908 242222 11960
rect 246298 11908 246304 11960
rect 246356 11948 246362 11960
rect 340966 11948 340972 11960
rect 246356 11920 340972 11948
rect 246356 11908 246362 11920
rect 340966 11908 340972 11920
rect 341024 11908 341030 11960
rect 405826 11908 405832 11960
rect 405884 11948 405890 11960
rect 494790 11948 494796 11960
rect 405884 11920 494796 11948
rect 405884 11908 405890 11920
rect 494790 11908 494796 11920
rect 494848 11908 494854 11960
rect 223574 11840 223580 11892
rect 223632 11880 223638 11892
rect 331214 11880 331220 11892
rect 223632 11852 331220 11880
rect 223632 11840 223638 11852
rect 331214 11840 331220 11852
rect 331272 11840 331278 11892
rect 405918 11840 405924 11892
rect 405976 11880 405982 11892
rect 521654 11880 521660 11892
rect 405976 11852 521660 11880
rect 405976 11840 405982 11852
rect 521654 11840 521660 11852
rect 521712 11840 521718 11892
rect 189166 11772 189172 11824
rect 189224 11812 189230 11824
rect 209774 11812 209780 11824
rect 189224 11784 209780 11812
rect 189224 11772 189230 11784
rect 209774 11772 209780 11784
rect 209832 11772 209838 11824
rect 223666 11772 223672 11824
rect 223724 11812 223730 11824
rect 334618 11812 334624 11824
rect 223724 11784 334624 11812
rect 223724 11772 223730 11784
rect 334618 11772 334624 11784
rect 334676 11772 334682 11824
rect 337470 11772 337476 11824
rect 337528 11812 337534 11824
rect 352190 11812 352196 11824
rect 337528 11784 352196 11812
rect 337528 11772 337534 11784
rect 352190 11772 352196 11784
rect 352248 11772 352254 11824
rect 372706 11772 372712 11824
rect 372764 11812 372770 11824
rect 404446 11812 404452 11824
rect 372764 11784 404452 11812
rect 372764 11772 372770 11784
rect 404446 11772 404452 11784
rect 404504 11772 404510 11824
rect 407206 11772 407212 11824
rect 407264 11812 407270 11824
rect 525426 11812 525432 11824
rect 407264 11784 525432 11812
rect 407264 11772 407270 11784
rect 525426 11772 525432 11784
rect 525484 11772 525490 11824
rect 157794 11704 157800 11756
rect 157852 11744 157858 11756
rect 173986 11744 173992 11756
rect 157852 11716 173992 11744
rect 157852 11704 157858 11716
rect 173986 11704 173992 11716
rect 174044 11704 174050 11756
rect 189074 11704 189080 11756
rect 189132 11744 189138 11756
rect 214466 11744 214472 11756
rect 189132 11716 214472 11744
rect 189132 11704 189138 11716
rect 214466 11704 214472 11716
rect 214524 11704 214530 11756
rect 225046 11704 225052 11756
rect 225104 11744 225110 11756
rect 338666 11744 338672 11756
rect 225104 11716 338672 11744
rect 225104 11704 225110 11716
rect 338666 11704 338672 11716
rect 338724 11704 338730 11756
rect 338758 11704 338764 11756
rect 338816 11744 338822 11756
rect 351914 11744 351920 11756
rect 338816 11716 351920 11744
rect 338816 11704 338822 11716
rect 351914 11704 351920 11716
rect 351972 11704 351978 11756
rect 363506 11704 363512 11756
rect 363564 11744 363570 11756
rect 372890 11744 372896 11756
rect 363564 11716 372896 11744
rect 363564 11704 363570 11716
rect 372890 11704 372896 11716
rect 372948 11704 372954 11756
rect 373994 11704 374000 11756
rect 374052 11744 374058 11756
rect 407114 11744 407120 11756
rect 374052 11716 407120 11744
rect 374052 11704 374058 11716
rect 407114 11704 407120 11716
rect 407172 11704 407178 11756
rect 408586 11704 408592 11756
rect 408644 11744 408650 11756
rect 532050 11744 532056 11756
rect 408644 11716 532056 11744
rect 408644 11704 408650 11716
rect 532050 11704 532056 11716
rect 532108 11704 532114 11756
rect 393314 10956 393320 11008
rect 393372 10996 393378 11008
rect 399478 10996 399484 11008
rect 393372 10968 399484 10996
rect 393372 10956 393378 10968
rect 399478 10956 399484 10968
rect 399536 10956 399542 11008
rect 280706 10616 280712 10668
rect 280764 10656 280770 10668
rect 336734 10656 336740 10668
rect 280764 10628 336740 10656
rect 280764 10616 280770 10628
rect 336734 10616 336740 10628
rect 336792 10616 336798 10668
rect 262490 10548 262496 10600
rect 262548 10588 262554 10600
rect 332686 10588 332692 10600
rect 262548 10560 332692 10588
rect 262548 10548 262554 10560
rect 332686 10548 332692 10560
rect 332744 10548 332750 10600
rect 382366 10548 382372 10600
rect 382424 10588 382430 10600
rect 436738 10588 436744 10600
rect 382424 10560 436744 10588
rect 382424 10548 382430 10560
rect 436738 10548 436744 10560
rect 436796 10548 436802 10600
rect 191834 10480 191840 10532
rect 191892 10520 191898 10532
rect 221090 10520 221096 10532
rect 191892 10492 221096 10520
rect 191892 10480 191898 10492
rect 221090 10480 221096 10492
rect 221148 10480 221154 10532
rect 241698 10480 241704 10532
rect 241756 10520 241762 10532
rect 325878 10520 325884 10532
rect 241756 10492 325884 10520
rect 241756 10480 241762 10492
rect 325878 10480 325884 10492
rect 325936 10480 325942 10532
rect 398834 10480 398840 10532
rect 398892 10520 398898 10532
rect 497090 10520 497096 10532
rect 398892 10492 497096 10520
rect 398892 10480 398898 10492
rect 497090 10480 497096 10492
rect 497148 10480 497154 10532
rect 218146 10412 218152 10464
rect 218204 10452 218210 10464
rect 305638 10452 305644 10464
rect 218204 10424 305644 10452
rect 218204 10412 218210 10424
rect 305638 10412 305644 10424
rect 305696 10412 305702 10464
rect 330570 10412 330576 10464
rect 330628 10452 330634 10464
rect 345106 10452 345112 10464
rect 330628 10424 345112 10452
rect 330628 10412 330634 10424
rect 345106 10412 345112 10424
rect 345164 10412 345170 10464
rect 345658 10412 345664 10464
rect 345716 10452 345722 10464
rect 354674 10452 354680 10464
rect 345716 10424 354680 10452
rect 345716 10412 345722 10424
rect 354674 10412 354680 10424
rect 354732 10412 354738 10464
rect 367738 10412 367744 10464
rect 367796 10452 367802 10464
rect 379514 10452 379520 10464
rect 367796 10424 379520 10452
rect 367796 10412 367802 10424
rect 379514 10412 379520 10424
rect 379572 10412 379578 10464
rect 400214 10412 400220 10464
rect 400272 10452 400278 10464
rect 500586 10452 500592 10464
rect 400272 10424 500592 10452
rect 400272 10412 400278 10424
rect 500586 10412 500592 10424
rect 500644 10412 500650 10464
rect 143534 10344 143540 10396
rect 143592 10384 143598 10396
rect 169938 10384 169944 10396
rect 143592 10356 169944 10384
rect 143592 10344 143598 10356
rect 169938 10344 169944 10356
rect 169996 10344 170002 10396
rect 186314 10344 186320 10396
rect 186372 10384 186378 10396
rect 203426 10384 203432 10396
rect 186372 10356 203432 10384
rect 186372 10344 186378 10356
rect 203426 10344 203432 10356
rect 203484 10344 203490 10396
rect 219526 10344 219532 10396
rect 219584 10384 219590 10396
rect 316034 10384 316040 10396
rect 219584 10356 316040 10384
rect 219584 10344 219590 10356
rect 316034 10344 316040 10356
rect 316092 10344 316098 10396
rect 316678 10344 316684 10396
rect 316736 10384 316742 10396
rect 335354 10384 335360 10396
rect 316736 10356 335360 10384
rect 316736 10344 316742 10356
rect 335354 10344 335360 10356
rect 335412 10344 335418 10396
rect 337562 10344 337568 10396
rect 337620 10384 337626 10396
rect 348326 10384 348332 10396
rect 337620 10356 348332 10384
rect 337620 10344 337626 10356
rect 348326 10344 348332 10356
rect 348384 10344 348390 10396
rect 377490 10344 377496 10396
rect 377548 10384 377554 10396
rect 397730 10384 397736 10396
rect 377548 10356 397736 10384
rect 377548 10344 377554 10356
rect 397730 10344 397736 10356
rect 397788 10344 397794 10396
rect 401594 10344 401600 10396
rect 401652 10384 401658 10396
rect 507210 10384 507216 10396
rect 401652 10356 507216 10384
rect 401652 10344 401658 10356
rect 507210 10344 507216 10356
rect 507268 10344 507274 10396
rect 141418 10276 141424 10328
rect 141476 10316 141482 10328
rect 168374 10316 168380 10328
rect 141476 10288 168380 10316
rect 141476 10276 141482 10288
rect 168374 10276 168380 10288
rect 168432 10276 168438 10328
rect 187694 10276 187700 10328
rect 187752 10316 187758 10328
rect 207106 10316 207112 10328
rect 187752 10288 207112 10316
rect 187752 10276 187758 10288
rect 207106 10276 207112 10288
rect 207164 10276 207170 10328
rect 209866 10276 209872 10328
rect 209924 10316 209930 10328
rect 317506 10316 317512 10328
rect 209924 10288 317512 10316
rect 209924 10276 209930 10288
rect 317506 10276 317512 10288
rect 317564 10276 317570 10328
rect 336090 10276 336096 10328
rect 336148 10316 336154 10328
rect 347866 10316 347872 10328
rect 336148 10288 347872 10316
rect 336148 10276 336154 10288
rect 347866 10276 347872 10288
rect 347924 10276 347930 10328
rect 371510 10276 371516 10328
rect 371568 10316 371574 10328
rect 400858 10316 400864 10328
rect 371568 10288 400864 10316
rect 371568 10276 371574 10288
rect 400858 10276 400864 10288
rect 400916 10276 400922 10328
rect 409874 10276 409880 10328
rect 409932 10316 409938 10328
rect 536098 10316 536104 10328
rect 409932 10288 536104 10316
rect 409932 10276 409938 10288
rect 536098 10276 536104 10288
rect 536156 10276 536162 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 248782 9324 248788 9376
rect 248840 9364 248846 9376
rect 328454 9364 328460 9376
rect 248840 9336 328460 9364
rect 248840 9324 248846 9336
rect 328454 9324 328460 9336
rect 328512 9324 328518 9376
rect 211614 9256 211620 9308
rect 211672 9296 211678 9308
rect 292574 9296 292580 9308
rect 211672 9268 292580 9296
rect 211672 9256 211678 9268
rect 292574 9256 292580 9268
rect 292632 9256 292638 9308
rect 195606 9188 195612 9240
rect 195664 9228 195670 9240
rect 313274 9228 313280 9240
rect 195664 9200 313280 9228
rect 195664 9188 195670 9200
rect 313274 9188 313280 9200
rect 313332 9188 313338 9240
rect 174262 9120 174268 9172
rect 174320 9160 174326 9172
rect 297358 9160 297364 9172
rect 174320 9132 297364 9160
rect 174320 9120 174326 9132
rect 297358 9120 297364 9132
rect 297416 9120 297422 9172
rect 329650 9120 329656 9172
rect 329708 9160 329714 9172
rect 343726 9160 343732 9172
rect 329708 9132 343732 9160
rect 329708 9120 329714 9132
rect 343726 9120 343732 9132
rect 343784 9120 343790 9172
rect 394786 9120 394792 9172
rect 394844 9160 394850 9172
rect 482830 9160 482836 9172
rect 394844 9132 482836 9160
rect 394844 9120 394850 9132
rect 482830 9120 482836 9132
rect 482888 9120 482894 9172
rect 181438 9052 181444 9104
rect 181496 9092 181502 9104
rect 307110 9092 307116 9104
rect 181496 9064 307116 9092
rect 181496 9052 181502 9064
rect 307110 9052 307116 9064
rect 307168 9052 307174 9104
rect 307754 9052 307760 9104
rect 307812 9092 307818 9104
rect 332594 9092 332600 9104
rect 307812 9064 332600 9092
rect 307812 9052 307818 9064
rect 332594 9052 332600 9064
rect 332652 9052 332658 9104
rect 404354 9052 404360 9104
rect 404412 9092 404418 9104
rect 514754 9092 514760 9104
rect 404412 9064 514760 9092
rect 404412 9052 404418 9064
rect 514754 9052 514760 9064
rect 514812 9052 514818 9104
rect 136450 8984 136456 9036
rect 136508 9024 136514 9036
rect 166994 9024 167000 9036
rect 136508 8996 167000 9024
rect 136508 8984 136514 8996
rect 166994 8984 167000 8996
rect 167052 8984 167058 9036
rect 291286 8984 291292 9036
rect 291344 9024 291350 9036
rect 555418 9024 555424 9036
rect 291344 8996 555424 9024
rect 291344 8984 291350 8996
rect 555418 8984 555424 8996
rect 555476 8984 555482 9036
rect 129366 8916 129372 8968
rect 129424 8956 129430 8968
rect 165706 8956 165712 8968
rect 129424 8928 165712 8956
rect 129424 8916 129430 8928
rect 165706 8916 165712 8928
rect 165764 8916 165770 8968
rect 284386 8916 284392 8968
rect 284444 8956 284450 8968
rect 291838 8956 291844 8968
rect 284444 8928 291844 8956
rect 284444 8916 284450 8928
rect 291838 8916 291844 8928
rect 291896 8916 291902 8968
rect 292666 8916 292672 8968
rect 292724 8956 292730 8968
rect 576302 8956 576308 8968
rect 292724 8928 576308 8956
rect 292724 8916 292730 8928
rect 576302 8916 576308 8928
rect 576360 8916 576366 8968
rect 300486 8168 300492 8220
rect 300544 8208 300550 8220
rect 302326 8208 302332 8220
rect 300544 8180 302332 8208
rect 300544 8168 300550 8180
rect 302326 8168 302332 8180
rect 302384 8168 302390 8220
rect 207014 7896 207020 7948
rect 207072 7936 207078 7948
rect 274818 7936 274824 7948
rect 207072 7908 274824 7936
rect 207072 7896 207078 7908
rect 274818 7896 274824 7908
rect 274876 7896 274882 7948
rect 277486 7896 277492 7948
rect 277544 7936 277550 7948
rect 299566 7936 299572 7948
rect 277544 7908 299572 7936
rect 277544 7896 277550 7908
rect 299566 7896 299572 7908
rect 299624 7896 299630 7948
rect 305546 7896 305552 7948
rect 305604 7936 305610 7948
rect 320818 7936 320824 7948
rect 305604 7908 320824 7936
rect 305604 7896 305610 7908
rect 320818 7896 320824 7908
rect 320876 7896 320882 7948
rect 252462 7828 252468 7880
rect 252520 7868 252526 7880
rect 324314 7868 324320 7880
rect 252520 7840 324320 7868
rect 252520 7828 252526 7840
rect 324314 7828 324320 7840
rect 324372 7828 324378 7880
rect 206186 7760 206192 7812
rect 206244 7800 206250 7812
rect 311158 7800 311164 7812
rect 206244 7772 311164 7800
rect 206244 7760 206250 7772
rect 311158 7760 311164 7772
rect 311216 7760 311222 7812
rect 323578 7760 323584 7812
rect 323636 7800 323642 7812
rect 341058 7800 341064 7812
rect 323636 7772 341064 7800
rect 323636 7760 323642 7772
rect 341058 7760 341064 7772
rect 341116 7760 341122 7812
rect 392578 7760 392584 7812
rect 392636 7800 392642 7812
rect 443822 7800 443828 7812
rect 392636 7772 443828 7800
rect 392636 7760 392642 7772
rect 443822 7760 443828 7772
rect 443880 7760 443886 7812
rect 234890 7692 234896 7744
rect 234948 7732 234954 7744
rect 348510 7732 348516 7744
rect 234948 7704 348516 7732
rect 234948 7692 234954 7704
rect 348510 7692 348516 7704
rect 348568 7692 348574 7744
rect 417050 7692 417056 7744
rect 417108 7732 417114 7744
rect 560846 7732 560852 7744
rect 417108 7704 560852 7732
rect 417108 7692 417114 7704
rect 560846 7692 560852 7704
rect 560904 7692 560910 7744
rect 154206 7624 154212 7676
rect 154264 7664 154270 7676
rect 172514 7664 172520 7676
rect 154264 7636 172520 7664
rect 154264 7624 154270 7636
rect 172514 7624 172520 7636
rect 172572 7624 172578 7676
rect 185026 7624 185032 7676
rect 185084 7664 185090 7676
rect 196802 7664 196808 7676
rect 185084 7636 196808 7664
rect 185084 7624 185090 7636
rect 196802 7624 196808 7636
rect 196860 7624 196866 7676
rect 208486 7624 208492 7676
rect 208544 7664 208550 7676
rect 278314 7664 278320 7676
rect 208544 7636 278320 7664
rect 208544 7624 208550 7636
rect 278314 7624 278320 7636
rect 278372 7624 278378 7676
rect 284478 7624 284484 7676
rect 284536 7664 284542 7676
rect 547874 7664 547880 7676
rect 284536 7636 547880 7664
rect 284536 7624 284542 7636
rect 547874 7624 547880 7636
rect 547932 7624 547938 7676
rect 132954 7556 132960 7608
rect 133012 7596 133018 7608
rect 165614 7596 165620 7608
rect 133012 7568 165620 7596
rect 133012 7556 133018 7568
rect 165614 7556 165620 7568
rect 165672 7556 165678 7608
rect 185118 7556 185124 7608
rect 185176 7596 185182 7608
rect 200298 7596 200304 7608
rect 185176 7568 200304 7596
rect 185176 7556 185182 7568
rect 200298 7556 200304 7568
rect 200356 7556 200362 7608
rect 208394 7556 208400 7608
rect 208452 7596 208458 7608
rect 281902 7596 281908 7608
rect 208452 7568 281908 7596
rect 208452 7556 208458 7568
rect 281902 7556 281908 7568
rect 281960 7556 281966 7608
rect 285674 7556 285680 7608
rect 285732 7596 285738 7608
rect 551462 7596 551468 7608
rect 285732 7568 551468 7596
rect 285732 7556 285738 7568
rect 551462 7556 551468 7568
rect 551520 7556 551526 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 151078 6848 151084 6860
rect 3476 6820 151084 6848
rect 3476 6808 3482 6820
rect 151078 6808 151084 6820
rect 151136 6808 151142 6860
rect 270034 6536 270040 6588
rect 270092 6576 270098 6588
rect 279418 6576 279424 6588
rect 270092 6548 279424 6576
rect 270092 6536 270098 6548
rect 279418 6536 279424 6548
rect 279476 6536 279482 6588
rect 245194 6468 245200 6520
rect 245252 6508 245258 6520
rect 327074 6508 327080 6520
rect 245252 6480 327080 6508
rect 245252 6468 245258 6480
rect 327074 6468 327080 6480
rect 327132 6468 327138 6520
rect 216858 6400 216864 6452
rect 216916 6440 216922 6452
rect 312538 6440 312544 6452
rect 216916 6412 312544 6440
rect 216916 6400 216922 6412
rect 312538 6400 312544 6412
rect 312596 6400 312602 6452
rect 188522 6332 188528 6384
rect 188580 6372 188586 6384
rect 302878 6372 302884 6384
rect 188580 6344 302884 6372
rect 188580 6332 188586 6344
rect 302878 6332 302884 6344
rect 302936 6332 302942 6384
rect 422294 6332 422300 6384
rect 422352 6372 422358 6384
rect 468754 6372 468760 6384
rect 422352 6344 468760 6372
rect 422352 6332 422358 6344
rect 468754 6332 468760 6344
rect 468812 6332 468818 6384
rect 277394 6264 277400 6316
rect 277452 6304 277458 6316
rect 523034 6304 523040 6316
rect 277452 6276 523040 6304
rect 277452 6264 277458 6276
rect 523034 6264 523040 6276
rect 523092 6264 523098 6316
rect 150618 6196 150624 6248
rect 150676 6236 150682 6248
rect 171134 6236 171140 6248
rect 150676 6208 171140 6236
rect 150676 6196 150682 6208
rect 171134 6196 171140 6208
rect 171192 6196 171198 6248
rect 205634 6196 205640 6248
rect 205692 6236 205698 6248
rect 271230 6236 271236 6248
rect 205692 6208 271236 6236
rect 205692 6196 205698 6208
rect 271230 6196 271236 6208
rect 271288 6196 271294 6248
rect 278774 6196 278780 6248
rect 278832 6236 278838 6248
rect 526622 6236 526628 6248
rect 278832 6208 526628 6236
rect 278832 6196 278838 6208
rect 526622 6196 526628 6208
rect 526680 6196 526686 6248
rect 160094 6128 160100 6180
rect 160152 6168 160158 6180
rect 206278 6168 206284 6180
rect 160152 6140 206284 6168
rect 160152 6128 160158 6140
rect 206278 6128 206284 6140
rect 206336 6128 206342 6180
rect 212534 6128 212540 6180
rect 212592 6168 212598 6180
rect 280062 6168 280068 6180
rect 212592 6140 280068 6168
rect 212592 6128 212598 6140
rect 280062 6128 280068 6140
rect 280120 6128 280126 6180
rect 284294 6128 284300 6180
rect 284352 6168 284358 6180
rect 544378 6168 544384 6180
rect 284352 6140 544384 6168
rect 284352 6128 284358 6140
rect 544378 6128 544384 6140
rect 544436 6128 544442 6180
rect 211798 5108 211804 5160
rect 211856 5148 211862 5160
rect 285398 5148 285404 5160
rect 211856 5120 285404 5148
rect 211856 5108 211862 5120
rect 285398 5108 285404 5120
rect 285456 5108 285462 5160
rect 223942 5040 223948 5092
rect 224000 5080 224006 5092
rect 321646 5080 321652 5092
rect 224000 5052 321652 5080
rect 224000 5040 224006 5052
rect 321646 5040 321652 5052
rect 321704 5040 321710 5092
rect 192018 4972 192024 5024
rect 192076 5012 192082 5024
rect 304258 5012 304264 5024
rect 192076 4984 304264 5012
rect 192076 4972 192082 4984
rect 304258 4972 304264 4984
rect 304316 4972 304322 5024
rect 240778 4904 240784 4956
rect 240836 4944 240842 4956
rect 370590 4944 370596 4956
rect 240836 4916 370596 4944
rect 240836 4904 240842 4916
rect 370590 4904 370596 4916
rect 370648 4904 370654 4956
rect 418154 4904 418160 4956
rect 418212 4944 418218 4956
rect 564434 4944 564440 4956
rect 418212 4916 564440 4944
rect 418212 4904 418218 4916
rect 564434 4904 564440 4916
rect 564492 4904 564498 4956
rect 161290 4836 161296 4888
rect 161348 4876 161354 4888
rect 173894 4876 173900 4888
rect 161348 4848 173900 4876
rect 161348 4836 161354 4848
rect 173894 4836 173900 4848
rect 173952 4836 173958 4888
rect 204346 4836 204352 4888
rect 204404 4876 204410 4888
rect 264146 4876 264152 4888
rect 204404 4848 264152 4876
rect 204404 4836 204410 4848
rect 264146 4836 264152 4848
rect 264204 4836 264210 4888
rect 269114 4836 269120 4888
rect 269172 4876 269178 4888
rect 487154 4876 487160 4888
rect 269172 4848 487160 4876
rect 269172 4836 269178 4848
rect 487154 4836 487160 4848
rect 487212 4836 487218 4888
rect 147674 4768 147680 4820
rect 147732 4808 147738 4820
rect 169846 4808 169852 4820
rect 147732 4780 169852 4808
rect 147732 4768 147738 4780
rect 169846 4768 169852 4780
rect 169904 4768 169910 4820
rect 185578 4768 185584 4820
rect 185636 4808 185642 4820
rect 193214 4808 193220 4820
rect 185636 4780 193220 4808
rect 185636 4768 185642 4780
rect 193214 4768 193220 4780
rect 193272 4768 193278 4820
rect 204254 4768 204260 4820
rect 204312 4808 204318 4820
rect 267734 4808 267740 4820
rect 204312 4780 267740 4808
rect 204312 4768 204318 4780
rect 267734 4768 267740 4780
rect 267792 4768 267798 4820
rect 270494 4768 270500 4820
rect 270552 4808 270558 4820
rect 498194 4808 498200 4820
rect 270552 4780 498200 4808
rect 270552 4768 270558 4780
rect 498194 4768 498200 4780
rect 498252 4768 498258 4820
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 337470 3992 337476 4004
rect 333940 3964 337476 3992
rect 333940 3952 333946 3964
rect 337470 3952 337476 3964
rect 337528 3952 337534 4004
rect 168374 3884 168380 3936
rect 168432 3924 168438 3936
rect 171778 3924 171784 3936
rect 168432 3896 171784 3924
rect 168432 3884 168438 3896
rect 171778 3884 171784 3896
rect 171836 3884 171842 3936
rect 319714 3884 319720 3936
rect 319772 3924 319778 3936
rect 337562 3924 337568 3936
rect 319772 3896 337568 3924
rect 319772 3884 319778 3896
rect 337562 3884 337568 3896
rect 337620 3884 337626 3936
rect 301958 3816 301964 3868
rect 302016 3856 302022 3868
rect 329650 3856 329656 3868
rect 302016 3828 329656 3856
rect 302016 3816 302022 3828
rect 329650 3816 329656 3828
rect 329708 3816 329714 3868
rect 266538 3748 266544 3800
rect 266596 3788 266602 3800
rect 307754 3788 307760 3800
rect 266596 3760 307760 3788
rect 266596 3748 266602 3760
rect 307754 3748 307760 3760
rect 307812 3748 307818 3800
rect 316218 3748 316224 3800
rect 316276 3788 316282 3800
rect 336090 3788 336096 3800
rect 316276 3760 336096 3788
rect 316276 3748 316282 3760
rect 336090 3748 336096 3760
rect 336148 3748 336154 3800
rect 234706 3680 234712 3732
rect 234764 3720 234770 3732
rect 252462 3720 252468 3732
rect 234764 3692 252468 3720
rect 234764 3680 234770 3692
rect 252462 3680 252468 3692
rect 252520 3680 252526 3732
rect 259546 3680 259552 3732
rect 259604 3720 259610 3732
rect 301590 3720 301596 3732
rect 259604 3692 301596 3720
rect 259604 3680 259610 3692
rect 301590 3680 301596 3692
rect 301648 3680 301654 3732
rect 312630 3680 312636 3732
rect 312688 3720 312694 3732
rect 330478 3720 330484 3732
rect 312688 3692 330484 3720
rect 312688 3680 312694 3692
rect 330478 3680 330484 3692
rect 330536 3680 330542 3732
rect 335998 3680 336004 3732
rect 336056 3720 336062 3732
rect 402514 3720 402520 3732
rect 336056 3692 402520 3720
rect 336056 3680 336062 3692
rect 402514 3680 402520 3692
rect 402572 3680 402578 3732
rect 413278 3680 413284 3732
rect 413336 3720 413342 3732
rect 454494 3720 454500 3732
rect 413336 3692 454500 3720
rect 413336 3680 413342 3692
rect 454494 3680 454500 3692
rect 454552 3680 454558 3732
rect 175458 3612 175464 3664
rect 175516 3652 175522 3664
rect 177298 3652 177304 3664
rect 175516 3624 177304 3652
rect 175516 3612 175522 3624
rect 177298 3612 177304 3624
rect 177356 3612 177362 3664
rect 252370 3612 252376 3664
rect 252428 3652 252434 3664
rect 307018 3652 307024 3664
rect 252428 3624 307024 3652
rect 252428 3612 252434 3624
rect 307018 3612 307024 3624
rect 307076 3612 307082 3664
rect 309042 3612 309048 3664
rect 309100 3652 309106 3664
rect 330570 3652 330576 3664
rect 309100 3624 330576 3652
rect 309100 3612 309106 3624
rect 330570 3612 330576 3624
rect 330628 3612 330634 3664
rect 337378 3612 337384 3664
rect 337436 3652 337442 3664
rect 352834 3652 352840 3664
rect 337436 3624 352840 3652
rect 337436 3612 337442 3624
rect 352834 3612 352840 3624
rect 352892 3612 352898 3664
rect 370498 3612 370504 3664
rect 370556 3652 370562 3664
rect 381170 3652 381176 3664
rect 370556 3624 381176 3652
rect 370556 3612 370562 3624
rect 381170 3612 381176 3624
rect 381228 3612 381234 3664
rect 381538 3612 381544 3664
rect 381596 3652 381602 3664
rect 388254 3652 388260 3664
rect 381596 3624 388260 3652
rect 381596 3612 381602 3624
rect 388254 3612 388260 3624
rect 388312 3612 388318 3664
rect 390554 3612 390560 3664
rect 390612 3652 390618 3664
rect 390612 3624 392072 3652
rect 390612 3612 390618 3624
rect 151814 3544 151820 3596
rect 151872 3584 151878 3596
rect 153010 3584 153016 3596
rect 151872 3556 153016 3584
rect 151872 3544 151878 3556
rect 153010 3544 153016 3556
rect 153068 3544 153074 3596
rect 167178 3544 167184 3596
rect 167236 3584 167242 3596
rect 273898 3584 273904 3596
rect 167236 3556 273904 3584
rect 167236 3544 167242 3556
rect 273898 3544 273904 3556
rect 273956 3544 273962 3596
rect 294874 3544 294880 3596
rect 294932 3584 294938 3596
rect 323578 3584 323584 3596
rect 294932 3556 323584 3584
rect 294932 3544 294938 3556
rect 323578 3544 323584 3556
rect 323636 3544 323642 3596
rect 330386 3544 330392 3596
rect 330444 3584 330450 3596
rect 338758 3584 338764 3596
rect 330444 3556 338764 3584
rect 330444 3544 330450 3556
rect 338758 3544 338764 3556
rect 338816 3544 338822 3596
rect 348510 3544 348516 3596
rect 348568 3584 348574 3596
rect 374086 3584 374092 3596
rect 348568 3556 374092 3584
rect 348568 3544 348574 3556
rect 374086 3544 374092 3556
rect 374144 3544 374150 3596
rect 381630 3544 381636 3596
rect 381688 3584 381694 3596
rect 390278 3584 390284 3596
rect 381688 3556 390284 3584
rect 381688 3544 381694 3556
rect 390278 3544 390284 3556
rect 390336 3544 390342 3596
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141418 3516 141424 3528
rect 140096 3488 141424 3516
rect 140096 3476 140102 3488
rect 141418 3476 141424 3488
rect 141476 3476 141482 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 277486 3516 277492 3528
rect 149572 3488 277492 3516
rect 149572 3476 149578 3488
rect 277486 3476 277492 3488
rect 277544 3476 277550 3528
rect 287790 3476 287796 3528
rect 287848 3516 287854 3528
rect 319438 3516 319444 3528
rect 287848 3488 319444 3516
rect 287848 3476 287854 3488
rect 319438 3476 319444 3488
rect 319496 3476 319502 3528
rect 323302 3476 323308 3528
rect 323360 3516 323366 3528
rect 334710 3516 334716 3528
rect 323360 3488 334716 3516
rect 323360 3476 323366 3488
rect 334710 3476 334716 3488
rect 334768 3476 334774 3528
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 342162 3516 342168 3528
rect 341024 3488 342168 3516
rect 341024 3476 341030 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 347038 3476 347044 3528
rect 347096 3516 347102 3528
rect 377674 3516 377680 3528
rect 347096 3488 377680 3516
rect 347096 3476 347102 3488
rect 377674 3476 377680 3488
rect 377732 3476 377738 3528
rect 382274 3476 382280 3528
rect 382332 3516 382338 3528
rect 383562 3516 383568 3528
rect 382332 3488 383568 3516
rect 382332 3476 382338 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 384298 3476 384304 3528
rect 384356 3516 384362 3528
rect 391842 3516 391848 3528
rect 384356 3488 391848 3516
rect 384356 3476 384362 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 392044 3516 392072 3624
rect 393958 3612 393964 3664
rect 394016 3652 394022 3664
rect 461578 3652 461584 3664
rect 394016 3624 461584 3652
rect 394016 3612 394022 3624
rect 461578 3612 461584 3624
rect 461636 3612 461642 3664
rect 487154 3612 487160 3664
rect 487212 3652 487218 3664
rect 494698 3652 494704 3664
rect 487212 3624 494704 3652
rect 487212 3612 487218 3624
rect 494698 3612 494704 3624
rect 494756 3612 494762 3664
rect 494790 3612 494796 3664
rect 494848 3652 494854 3664
rect 518342 3652 518348 3664
rect 494848 3624 518348 3652
rect 494848 3612 494854 3624
rect 518342 3612 518348 3624
rect 518400 3612 518406 3664
rect 399478 3544 399484 3596
rect 399536 3584 399542 3596
rect 475746 3584 475752 3596
rect 399536 3556 475752 3584
rect 399536 3544 399542 3556
rect 475746 3544 475752 3556
rect 475804 3544 475810 3596
rect 480254 3544 480260 3596
rect 480312 3584 480318 3596
rect 554958 3584 554964 3596
rect 480312 3556 554964 3584
rect 480312 3544 480318 3556
rect 554958 3544 554964 3556
rect 555016 3544 555022 3596
rect 555418 3544 555424 3596
rect 555476 3584 555482 3596
rect 569126 3584 569132 3596
rect 555476 3556 569132 3584
rect 555476 3544 555482 3556
rect 569126 3544 569132 3556
rect 569184 3544 569190 3596
rect 468662 3516 468668 3528
rect 392044 3488 468668 3516
rect 468662 3476 468668 3488
rect 468720 3476 468726 3528
rect 468754 3476 468760 3528
rect 468812 3516 468818 3528
rect 578602 3516 578608 3528
rect 468812 3488 578608 3516
rect 468812 3476 468818 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 128170 3408 128176 3460
rect 128228 3448 128234 3460
rect 269206 3448 269212 3460
rect 128228 3420 269212 3448
rect 128228 3408 128234 3420
rect 269206 3408 269212 3420
rect 269264 3408 269270 3460
rect 273622 3408 273628 3460
rect 273680 3448 273686 3460
rect 316678 3448 316684 3460
rect 273680 3420 316684 3448
rect 273680 3408 273686 3420
rect 316678 3408 316684 3420
rect 316736 3408 316742 3460
rect 329098 3408 329104 3460
rect 329156 3448 329162 3460
rect 562042 3448 562048 3460
rect 329156 3420 562048 3448
rect 329156 3408 329162 3420
rect 562042 3408 562048 3420
rect 562100 3408 562106 3460
rect 565078 3408 565084 3460
rect 565136 3448 565142 3460
rect 579798 3448 579804 3460
rect 565136 3420 579804 3448
rect 565136 3408 565142 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 177850 3380 177856 3392
rect 176712 3352 177856 3380
rect 176712 3340 176718 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 201494 3340 201500 3392
rect 201552 3380 201558 3392
rect 202690 3380 202696 3392
rect 201552 3352 202696 3380
rect 201552 3340 201558 3352
rect 202690 3340 202696 3352
rect 202748 3340 202754 3392
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 235810 3380 235816 3392
rect 234672 3352 235816 3380
rect 234672 3340 234678 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 355226 3340 355232 3392
rect 355284 3380 355290 3392
rect 356698 3380 356704 3392
rect 355284 3352 356704 3380
rect 355284 3340 355290 3352
rect 356698 3340 356704 3352
rect 356756 3340 356762 3392
rect 358722 3340 358728 3392
rect 358780 3380 358786 3392
rect 359458 3380 359464 3392
rect 358780 3352 359464 3380
rect 358780 3340 358786 3352
rect 359458 3340 359464 3352
rect 359516 3340 359522 3392
rect 365806 3340 365812 3392
rect 365864 3380 365870 3392
rect 367002 3380 367008 3392
rect 365864 3352 367008 3380
rect 365864 3340 365870 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 377398 3340 377404 3392
rect 377456 3380 377462 3392
rect 384758 3380 384764 3392
rect 377456 3352 384764 3380
rect 377456 3340 377462 3352
rect 384758 3340 384764 3352
rect 384816 3340 384822 3392
rect 390278 3340 390284 3392
rect 390336 3380 390342 3392
rect 394234 3380 394240 3392
rect 390336 3352 394240 3380
rect 390336 3340 390342 3352
rect 394234 3340 394240 3352
rect 394292 3340 394298 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 490742 3380 490748 3392
rect 489972 3352 490748 3380
rect 489972 3340 489978 3352
rect 490742 3340 490748 3352
rect 490800 3340 490806 3392
rect 184290 3272 184296 3324
rect 184348 3312 184354 3324
rect 189718 3312 189724 3324
rect 184348 3284 189724 3312
rect 184348 3272 184354 3284
rect 189718 3272 189724 3284
rect 189776 3272 189782 3324
rect 363598 3136 363604 3188
rect 363656 3176 363662 3188
rect 365806 3176 365812 3188
rect 363656 3148 365812 3176
rect 363656 3136 363662 3148
rect 365806 3136 365812 3148
rect 365864 3136 365870 3188
rect 366358 3068 366364 3120
rect 366416 3108 366422 3120
rect 369394 3108 369400 3120
rect 366416 3080 369400 3108
rect 366416 3068 366422 3080
rect 369394 3068 369400 3080
rect 369452 3068 369458 3120
rect 171962 3000 171968 3052
rect 172020 3040 172026 3052
rect 174538 3040 174544 3052
rect 172020 3012 174544 3040
rect 172020 3000 172026 3012
rect 174538 3000 174544 3012
rect 174596 3000 174602 3052
rect 184198 3000 184204 3052
rect 184256 3040 184262 3052
rect 186130 3040 186136 3052
rect 184256 3012 186136 3040
rect 184256 3000 184262 3012
rect 186130 3000 186136 3012
rect 186188 3000 186194 3052
rect 244918 3000 244924 3052
rect 244976 3040 244982 3052
rect 249978 3040 249984 3052
rect 244976 3012 249984 3040
rect 244976 3000 244982 3012
rect 249978 3000 249984 3012
rect 250036 3000 250042 3052
rect 337470 3000 337476 3052
rect 337528 3040 337534 3052
rect 342898 3040 342904 3052
rect 337528 3012 342904 3040
rect 337528 3000 337534 3012
rect 342898 3000 342904 3012
rect 342956 3000 342962 3052
rect 125870 2932 125876 2984
rect 125928 2972 125934 2984
rect 127618 2972 127624 2984
rect 125928 2944 127624 2972
rect 125928 2932 125934 2944
rect 127618 2932 127624 2944
rect 127676 2932 127682 2984
rect 340966 2932 340972 2984
rect 341024 2972 341030 2984
rect 345658 2972 345664 2984
rect 341024 2944 345664 2972
rect 341024 2932 341030 2944
rect 345658 2932 345664 2944
rect 345716 2932 345722 2984
rect 255866 2864 255872 2916
rect 255924 2904 255930 2916
rect 260098 2904 260104 2916
rect 255924 2876 260104 2904
rect 255924 2864 255930 2876
rect 260098 2864 260104 2876
rect 260156 2864 260162 2916
rect 333974 2796 333980 2848
rect 334032 2836 334038 2848
rect 508866 2836 508872 2848
rect 334032 2808 508872 2836
rect 334032 2796 334038 2808
rect 508866 2796 508872 2808
rect 508924 2796 508930 2848
rect 415394 2728 415400 2780
rect 415452 2768 415458 2780
rect 416682 2768 416688 2780
rect 415452 2740 416688 2768
rect 415452 2728 415458 2740
rect 416682 2728 416688 2740
rect 416740 2728 416746 2780
rect 215294 2388 215300 2440
rect 215352 2428 215358 2440
rect 306742 2428 306748 2440
rect 215352 2400 306748 2428
rect 215352 2388 215358 2400
rect 306742 2388 306748 2400
rect 306800 2388 306806 2440
rect 220814 2320 220820 2372
rect 220872 2360 220878 2372
rect 324406 2360 324412 2372
rect 220872 2332 324412 2360
rect 220872 2320 220878 2332
rect 324406 2320 324412 2332
rect 324464 2320 324470 2372
rect 222194 2252 222200 2304
rect 222252 2292 222258 2304
rect 327994 2292 328000 2304
rect 222252 2264 328000 2292
rect 222252 2252 222258 2264
rect 327994 2252 328000 2264
rect 328052 2252 328058 2304
rect 249794 2184 249800 2236
rect 249852 2224 249858 2236
rect 423766 2224 423772 2236
rect 249852 2196 423772 2224
rect 249852 2184 249858 2196
rect 423766 2184 423772 2196
rect 423824 2184 423830 2236
rect 263594 2116 263600 2168
rect 263652 2156 263658 2168
rect 473446 2156 473452 2168
rect 263652 2128 473452 2156
rect 263652 2116 263658 2128
rect 473446 2116 473452 2128
rect 473504 2116 473510 2168
rect 281534 2048 281540 2100
rect 281592 2088 281598 2100
rect 537202 2088 537208 2100
rect 281592 2060 537208 2088
rect 281592 2048 281598 2060
rect 537202 2048 537208 2060
rect 537260 2048 537266 2100
rect 440234 1912 440240 1964
rect 440292 1952 440298 1964
rect 441522 1952 441528 1964
rect 440292 1924 441528 1952
rect 440292 1912 440298 1924
rect 441522 1912 441528 1924
rect 441580 1912 441586 1964
rect 273254 1300 273260 1352
rect 273312 1340 273318 1352
rect 333974 1340 333980 1352
rect 273312 1312 333980 1340
rect 273312 1300 273318 1312
rect 333974 1300 333980 1312
rect 334032 1300 334038 1352
rect 267918 144 267924 196
rect 267976 184 267982 196
rect 487246 184 487252 196
rect 267976 156 487252 184
rect 267976 144 267982 156
rect 487246 144 487252 156
rect 487304 144 487310 196
rect 271874 76 271880 128
rect 271932 116 271938 128
rect 505554 116 505560 128
rect 271932 88 505560 116
rect 271932 76 271938 88
rect 505554 76 505560 88
rect 505612 76 505618 128
rect 280154 8 280160 60
rect 280212 48 280218 60
rect 529934 48 529940 60
rect 280212 20 529940 48
rect 280212 8 280218 20
rect 529934 8 529940 20
rect 529992 8 529998 60
<< via1 >>
rect 8116 700952 8168 701004
rect 19248 700952 19300 701004
rect 72976 700952 73028 701004
rect 397460 700952 397512 701004
rect 462320 700952 462372 701004
rect 22008 700340 22060 700392
rect 89168 700340 89220 700392
rect 138020 700340 138072 700392
rect 202788 700340 202840 700392
rect 21916 700272 21968 700324
rect 218980 700272 219032 700324
rect 302148 700272 302200 700324
rect 478512 700272 478564 700324
rect 527180 700272 527232 700324
rect 543464 700272 543516 700324
rect 22100 699660 22152 699712
rect 24308 699660 24360 699712
rect 302240 698912 302292 698964
rect 413652 698912 413704 698964
rect 527272 698232 527324 698284
rect 580172 698232 580224 698284
rect 16488 697620 16540 697672
rect 138020 697620 138072 697672
rect 22192 697552 22244 697604
rect 154120 697552 154172 697604
rect 2780 606432 2832 606484
rect 15844 606432 15896 606484
rect 21916 586440 21968 586492
rect 28172 586440 28224 586492
rect 144828 586440 144880 586492
rect 149980 586440 150032 586492
rect 302148 586440 302200 586492
rect 308496 586440 308548 586492
rect 424876 586440 424928 586492
rect 429936 586440 429988 586492
rect 21824 586100 21876 586152
rect 43352 586100 43404 586152
rect 23296 586032 23348 586084
rect 48504 586032 48556 586084
rect 266268 586032 266320 586084
rect 290004 586032 290056 586084
rect 302056 586032 302108 586084
rect 313556 586032 313608 586084
rect 546316 586032 546368 586084
rect 568856 586032 568908 586084
rect 21732 585964 21784 586016
rect 53472 585964 53524 586016
rect 261576 585964 261628 586016
rect 289912 585964 289964 586016
rect 301872 585964 301924 586016
rect 318616 585964 318668 586016
rect 541256 585964 541308 586016
rect 567476 585964 567528 586016
rect 29644 585896 29696 585948
rect 104072 585896 104124 585948
rect 256516 585896 256568 585948
rect 288532 585896 288584 585948
rect 303160 585896 303212 585948
rect 323676 585896 323728 585948
rect 536196 585896 536248 585948
rect 568672 585896 568724 585948
rect 21916 585828 21968 585880
rect 33232 585828 33284 585880
rect 35164 585828 35216 585880
rect 119252 585828 119304 585880
rect 251088 585828 251140 585880
rect 289820 585828 289872 585880
rect 302148 585828 302200 585880
rect 328736 585828 328788 585880
rect 531136 585828 531188 585880
rect 569960 585828 570012 585880
rect 23112 585760 23164 585812
rect 38292 585760 38344 585812
rect 39304 585760 39356 585812
rect 124312 585760 124364 585812
rect 241336 585760 241388 585812
rect 287612 585760 287664 585812
rect 303252 585760 303304 585812
rect 333796 585760 333848 585812
rect 521016 585760 521068 585812
rect 567568 585760 567620 585812
rect 281448 585148 281500 585200
rect 288624 585148 288676 585200
rect 424324 585148 424376 585200
rect 424876 585148 424928 585200
rect 561496 585148 561548 585200
rect 568764 585148 568816 585200
rect 300676 583312 300728 583364
rect 338856 583312 338908 583364
rect 17868 583244 17920 583296
rect 93952 583244 94004 583296
rect 235908 583244 235960 583296
rect 292580 583244 292632 583296
rect 300492 583244 300544 583296
rect 343916 583244 343968 583296
rect 17776 583176 17828 583228
rect 99012 583176 99064 583228
rect 231216 583176 231268 583228
rect 288808 583176 288860 583228
rect 300768 583176 300820 583228
rect 348976 583176 349028 583228
rect 515956 583176 516008 583228
rect 570328 583176 570380 583228
rect 15108 583108 15160 583160
rect 114192 583108 114244 583160
rect 220728 583108 220780 583160
rect 291476 583108 291528 583160
rect 299296 583108 299348 583160
rect 354036 583108 354088 583160
rect 510896 583108 510948 583160
rect 570144 583108 570196 583160
rect 15016 583040 15068 583092
rect 139492 583040 139544 583092
rect 216036 583040 216088 583092
rect 291200 583040 291252 583092
rect 300584 583040 300636 583092
rect 359096 583040 359148 583092
rect 500776 583040 500828 583092
rect 568948 583040 569000 583092
rect 19156 582972 19208 583024
rect 154764 582972 154816 583024
rect 200856 582972 200908 583024
rect 293224 582972 293276 583024
rect 301964 582972 302016 583024
rect 364156 582972 364208 583024
rect 465356 582972 465408 583024
rect 567660 582972 567712 583024
rect 195796 580524 195848 580576
rect 295340 580524 295392 580576
rect 299204 580524 299256 580576
rect 374276 580524 374328 580576
rect 185676 580456 185728 580508
rect 287796 580456 287848 580508
rect 302976 580456 303028 580508
rect 379336 580456 379388 580508
rect 190368 580388 190420 580440
rect 291844 580388 291896 580440
rect 295156 580388 295208 580440
rect 394516 580388 394568 580440
rect 475476 580388 475528 580440
rect 574192 580388 574244 580440
rect 180616 580320 180668 580372
rect 295432 580320 295484 580372
rect 297824 580320 297876 580372
rect 384396 580320 384448 580372
rect 460296 580320 460348 580372
rect 572720 580320 572772 580372
rect 165436 580252 165488 580304
rect 295524 580252 295576 580304
rect 299388 580252 299440 580304
rect 399576 580252 399628 580304
rect 455236 580252 455288 580304
rect 571432 580252 571484 580304
rect 299112 577600 299164 577652
rect 408500 577600 408552 577652
rect 297916 577532 297968 577584
rect 414020 577532 414072 577584
rect 169760 577464 169812 577516
rect 292672 577464 292724 577516
rect 295248 577464 295300 577516
rect 419540 577464 419592 577516
rect 17684 574812 17736 574864
rect 35164 574812 35216 574864
rect 13728 574744 13780 574796
rect 128360 574744 128412 574796
rect 16396 572296 16448 572348
rect 29644 572296 29696 572348
rect 19064 572228 19116 572280
rect 57980 572228 58032 572280
rect 20536 572160 20588 572212
rect 67640 572160 67692 572212
rect 525800 572160 525852 572212
rect 570236 572160 570288 572212
rect 20628 572092 20680 572144
rect 73160 572092 73212 572144
rect 270500 572092 270552 572144
rect 294604 572092 294656 572144
rect 495440 572092 495492 572144
rect 571524 572092 571576 572144
rect 19248 572024 19300 572076
rect 78680 572024 78732 572076
rect 245660 572024 245712 572076
rect 290096 572024 290148 572076
rect 469220 572024 469272 572076
rect 572812 572024 572864 572076
rect 20444 571956 20496 572008
rect 88340 571956 88392 572008
rect 158720 571956 158772 572008
rect 288716 571956 288768 572008
rect 444380 571956 444432 572008
rect 575480 571956 575532 572008
rect 577688 524424 577740 524476
rect 579620 524424 579672 524476
rect 2872 514768 2924 514820
rect 4804 514768 4856 514820
rect 2780 500964 2832 501016
rect 7564 500964 7616 501016
rect 577504 484576 577556 484628
rect 580632 484576 580684 484628
rect 3332 462340 3384 462392
rect 13084 462340 13136 462392
rect 285588 461592 285640 461644
rect 292672 461592 292724 461644
rect 296536 461592 296588 461644
rect 299388 461592 299440 461644
rect 399300 461592 399352 461644
rect 24952 461116 25004 461168
rect 99012 461116 99064 461168
rect 22100 461048 22152 461100
rect 23388 461048 23440 461100
rect 16396 460980 16448 461032
rect 17592 460980 17644 461032
rect 104394 461048 104446 461100
rect 20352 460912 20404 460964
rect 109454 460980 109506 461032
rect 391940 460980 391992 461032
rect 24860 460912 24912 460964
rect 139492 460912 139544 460964
rect 17776 460844 17828 460896
rect 24952 460844 25004 460896
rect 15016 460776 15068 460828
rect 24860 460776 24912 460828
rect 17684 460708 17736 460760
rect 119252 460844 119304 460896
rect 241336 460844 241388 460896
rect 287612 460844 287664 460896
rect 295156 460844 295208 460896
rect 296720 460912 296772 460964
rect 305092 460912 305144 460964
rect 404636 460912 404688 460964
rect 296628 460844 296680 460896
rect 297824 460844 297876 460896
rect 384396 460844 384448 460896
rect 391940 460844 391992 460896
rect 394516 460844 394568 460896
rect 445116 460844 445168 460896
rect 575480 460912 575532 460964
rect 470416 460844 470468 460896
rect 572812 460844 572864 460896
rect 246396 460776 246448 460828
rect 290188 460776 290240 460828
rect 300584 460776 300636 460828
rect 359096 460776 359148 460828
rect 495716 460776 495768 460828
rect 571524 460776 571576 460828
rect 256516 460708 256568 460760
rect 286324 460708 286376 460760
rect 288532 460708 288584 460760
rect 521016 460708 521068 460760
rect 567660 460708 567712 460760
rect 526076 460640 526128 460692
rect 570236 460640 570288 460692
rect 536196 460572 536248 460624
rect 568580 460572 568632 460624
rect 285496 460232 285548 460284
rect 295524 460232 295576 460284
rect 14924 460164 14976 460216
rect 129372 460164 129424 460216
rect 190460 460164 190512 460216
rect 291844 460164 291896 460216
rect 287704 460028 287756 460080
rect 288624 460028 288676 460080
rect 300400 460028 300452 460080
rect 301780 460028 301832 460080
rect 343916 460164 343968 460216
rect 13728 459892 13780 459944
rect 14924 459892 14976 459944
rect 301872 459892 301924 459944
rect 303068 459892 303120 459944
rect 570052 459756 570104 459808
rect 570236 459756 570288 459808
rect 572812 459620 572864 459672
rect 574100 459620 574152 459672
rect 291844 459552 291896 459604
rect 293960 459552 294012 459604
rect 298928 459552 298980 459604
rect 300584 459552 300636 459604
rect 434996 459552 435048 459604
rect 438124 459552 438176 459604
rect 571524 459552 571576 459604
rect 572996 459552 573048 459604
rect 22008 459484 22060 459536
rect 28172 459484 28224 459536
rect 144828 459484 144880 459536
rect 149980 459484 150032 459536
rect 195796 459484 195848 459536
rect 295340 459484 295392 459536
rect 302056 459484 302108 459536
rect 313556 459484 313608 459536
rect 424876 459484 424928 459536
rect 429936 459484 429988 459536
rect 546316 459484 546368 459536
rect 556160 459484 556212 459536
rect 20628 459416 20680 459468
rect 73712 459416 73764 459468
rect 185676 459416 185728 459468
rect 285404 459416 285456 459468
rect 287796 459416 287848 459468
rect 301872 459416 301924 459468
rect 389456 459416 389508 459468
rect 450176 459416 450228 459468
rect 564440 459416 564492 459468
rect 19064 459348 19116 459400
rect 58532 459348 58584 459400
rect 266268 459348 266320 459400
rect 290004 459348 290056 459400
rect 299204 459348 299256 459400
rect 374276 459348 374328 459400
rect 460296 459348 460348 459400
rect 572720 459348 572772 459400
rect 20444 459280 20496 459332
rect 88892 459280 88944 459332
rect 299296 459280 299348 459332
rect 354036 459280 354088 459332
rect 465356 459280 465408 459332
rect 567752 459280 567804 459332
rect 303068 459212 303120 459264
rect 318616 459212 318668 459264
rect 531136 459212 531188 459264
rect 569960 459212 570012 459264
rect 313280 459144 313332 459196
rect 323676 459144 323728 459196
rect 308496 459076 308548 459128
rect 580264 459076 580316 459128
rect 20536 458940 20588 458992
rect 21640 458940 21692 458992
rect 34520 458940 34572 458992
rect 38292 458940 38344 458992
rect 216036 458940 216088 458992
rect 288532 458940 288584 458992
rect 291200 458940 291252 458992
rect 68652 458872 68704 458924
rect 180616 458872 180668 458924
rect 292764 458872 292816 458924
rect 295432 458872 295484 458924
rect 17868 458804 17920 458856
rect 18788 458804 18840 458856
rect 19248 458804 19300 458856
rect 20352 458804 20404 458856
rect 78772 458804 78824 458856
rect 149980 458804 150032 458856
rect 288440 458804 288492 458856
rect 556436 458804 556488 458856
rect 571432 458804 571484 458856
rect 27804 458464 27856 458516
rect 33232 458464 33284 458516
rect 110420 458192 110472 458244
rect 114192 458192 114244 458244
rect 290004 458192 290056 458244
rect 290280 458192 290332 458244
rect 23296 458124 23348 458176
rect 30932 458124 30984 458176
rect 21916 458056 21968 458108
rect 23112 458056 23164 458108
rect 27804 458056 27856 458108
rect 63592 458124 63644 458176
rect 226156 458124 226208 458176
rect 287520 458124 287572 458176
rect 298008 458124 298060 458176
rect 369216 458192 369268 458244
rect 424324 458192 424376 458244
rect 424876 458192 424928 458244
rect 500776 458192 500828 458244
rect 569960 458192 570012 458244
rect 571524 458192 571576 458244
rect 572720 458192 572772 458244
rect 575480 458192 575532 458244
rect 568948 458124 569000 458176
rect 570604 458124 570656 458176
rect 23204 457920 23256 457972
rect 21732 457852 21784 457904
rect 53472 458056 53524 458108
rect 231216 458056 231268 458108
rect 288808 458056 288860 458108
rect 291292 458056 291344 458108
rect 300676 458056 300728 458108
rect 338856 458056 338908 458108
rect 505836 458056 505888 458108
rect 565912 458056 565964 458108
rect 30932 457784 30984 457836
rect 48504 457988 48556 458040
rect 251088 457988 251140 458040
rect 289820 457988 289872 458040
rect 303252 457988 303304 458040
rect 333796 457988 333848 458040
rect 510896 457988 510948 458040
rect 570144 457988 570196 458040
rect 302148 457920 302200 457972
rect 328736 457920 328788 457972
rect 515956 457920 516008 457972
rect 570328 457920 570380 457972
rect 541256 457852 541308 457904
rect 567568 457852 567620 457904
rect 300400 457580 300452 457632
rect 303252 457580 303304 457632
rect 261576 457512 261628 457564
rect 289084 457512 289136 457564
rect 289912 457512 289964 457564
rect 21824 457444 21876 457496
rect 23020 457444 23072 457496
rect 43352 457444 43404 457496
rect 235908 457444 235960 457496
rect 291200 457444 291252 457496
rect 292580 457444 292632 457496
rect 301964 457444 302016 457496
rect 303252 457444 303304 457496
rect 364156 457444 364208 457496
rect 21732 456832 21784 456884
rect 23204 456832 23256 456884
rect 22744 456764 22796 456816
rect 23296 456764 23348 456816
rect 570328 456764 570380 456816
rect 572812 456764 572864 456816
rect 299112 456696 299164 456748
rect 409696 456696 409748 456748
rect 301872 456628 301924 456680
rect 302976 456628 303028 456680
rect 379336 456628 379388 456680
rect 305000 456016 305052 456068
rect 419816 456016 419868 456068
rect 15108 455336 15160 455388
rect 17868 455336 17920 455388
rect 19156 455336 19208 455388
rect 154764 455336 154816 455388
rect 295248 455336 295300 455388
rect 305000 455336 305052 455388
rect 440056 455336 440108 455388
rect 564900 455336 564952 455388
rect 17224 454656 17276 454708
rect 17868 454656 17920 454708
rect 110420 454656 110472 454708
rect 564900 454656 564952 454708
rect 571616 454656 571668 454708
rect 21364 444320 21416 444372
rect 24860 444320 24912 444372
rect 219440 444320 219492 444372
rect 291476 444320 291528 444372
rect 300768 444320 300820 444372
rect 347780 444320 347832 444372
rect 438124 444320 438176 444372
rect 565544 444320 565596 444372
rect 270500 444252 270552 444304
rect 297180 444252 297232 444304
rect 474740 444252 474792 444304
rect 574192 444252 574244 444304
rect 291476 443912 291528 443964
rect 292856 443912 292908 443964
rect 23480 443640 23532 443692
rect 200120 443640 200172 443692
rect 300308 443504 300360 443556
rect 300768 443504 300820 443556
rect 565544 442960 565596 443012
rect 568856 442960 568908 443012
rect 164240 442892 164292 442944
rect 284300 442892 284352 442944
rect 169760 442824 169812 442876
rect 284944 442824 284996 442876
rect 285588 442824 285640 442876
rect 13176 442212 13228 442264
rect 23480 442212 23532 442264
rect 284300 442212 284352 442264
rect 285496 442212 285548 442264
rect 296812 442212 296864 442264
rect 284944 441872 284996 441924
rect 288624 441872 288676 441924
rect 3148 410048 3200 410100
rect 6184 410048 6236 410100
rect 2780 398760 2832 398812
rect 7656 398760 7708 398812
rect 577596 364692 577648 364744
rect 580632 364692 580684 364744
rect 2964 357416 3016 357468
rect 6276 357416 6328 357468
rect 3332 345312 3384 345364
rect 8944 345312 8996 345364
rect 17408 333956 17460 334008
rect 21364 333956 21416 334008
rect 570604 333956 570656 334008
rect 574468 333956 574520 334008
rect 300492 333616 300544 333668
rect 305000 333616 305052 333668
rect 285588 333276 285640 333328
rect 292764 333276 292816 333328
rect 295248 333276 295300 333328
rect 305092 333276 305144 333328
rect 501144 333276 501196 333328
rect 570604 333276 570656 333328
rect 20444 333208 20496 333260
rect 88892 333208 88944 333260
rect 284208 333208 284260 333260
rect 296812 333208 296864 333260
rect 475752 333208 475804 333260
rect 574192 333208 574244 333260
rect 18880 332936 18932 332988
rect 20444 332936 20496 332988
rect 20352 332868 20404 332920
rect 78772 332868 78824 332920
rect 20260 332800 20312 332852
rect 109132 332800 109184 332852
rect 20168 332732 20220 332784
rect 20352 332732 20404 332784
rect 21364 332732 21416 332784
rect 124312 332732 124364 332784
rect 299112 332732 299164 332784
rect 303712 332732 303764 332784
rect 14924 332664 14976 332716
rect 15108 332664 15160 332716
rect 129372 332664 129424 332716
rect 231216 332664 231268 332716
rect 291292 332664 291344 332716
rect 296628 332664 296680 332716
rect 384028 332664 384080 332716
rect 574192 332664 574244 332716
rect 575756 332664 575808 332716
rect 15016 332596 15068 332648
rect 139492 332596 139544 332648
rect 210976 332596 211028 332648
rect 287612 332596 287664 332648
rect 305092 332596 305144 332648
rect 419816 332596 419868 332648
rect 22744 332528 22796 332580
rect 3608 332460 3660 332512
rect 23112 332460 23164 332512
rect 23664 332528 23716 332580
rect 63592 332528 63644 332580
rect 144828 332528 144880 332580
rect 149612 332528 149664 332580
rect 246396 332528 246448 332580
rect 290188 332528 290240 332580
rect 301872 332528 301924 332580
rect 306380 332528 306432 332580
rect 48412 332460 48464 332512
rect 251088 332460 251140 332512
rect 289820 332460 289872 332512
rect 303068 332460 303120 332512
rect 318616 332528 318668 332580
rect 424324 332528 424376 332580
rect 424876 332528 424928 332580
rect 429936 332528 429988 332580
rect 445116 332528 445168 332580
rect 575664 332596 575716 332648
rect 311256 332460 311308 332512
rect 333796 332460 333848 332512
rect 536196 332460 536248 332512
rect 568580 332460 568632 332512
rect 22928 332392 22980 332444
rect 43352 332392 43404 332444
rect 256516 332392 256568 332444
rect 281356 332392 281408 332444
rect 281448 332392 281500 332444
rect 287704 332392 287756 332444
rect 302148 332392 302200 332444
rect 328736 332392 328788 332444
rect 541256 332392 541308 332444
rect 567568 332392 567620 332444
rect 22836 332324 22888 332376
rect 38292 332324 38344 332376
rect 261576 332324 261628 332376
rect 282184 332324 282236 332376
rect 303160 332324 303212 332376
rect 323676 332324 323728 332376
rect 546316 332324 546368 332376
rect 568672 332324 568724 332376
rect 23020 332256 23072 332308
rect 33232 332256 33284 332308
rect 266268 332256 266320 332308
rect 290280 332256 290332 332308
rect 302056 332256 302108 332308
rect 313556 332256 313608 332308
rect 21732 332188 21784 332240
rect 23664 332188 23716 332240
rect 281356 332188 281408 332240
rect 285680 332188 285732 332240
rect 308496 332188 308548 332240
rect 580540 332188 580592 332240
rect 300400 332120 300452 332172
rect 311256 332120 311308 332172
rect 21824 331984 21876 332036
rect 22744 331984 22796 332036
rect 190368 331916 190420 331968
rect 192116 331916 192168 331968
rect 561496 331916 561548 331968
rect 568764 331916 568816 331968
rect 570236 331916 570288 331968
rect 22100 331848 22152 331900
rect 22744 331848 22796 331900
rect 53472 331848 53524 331900
rect 185676 331848 185728 331900
rect 187608 331848 187660 331900
rect 282184 331848 282236 331900
rect 289084 331848 289136 331900
rect 292580 331848 292632 331900
rect 556436 331848 556488 331900
rect 569960 331848 570012 331900
rect 299020 331304 299072 331356
rect 302148 331304 302200 331356
rect 21916 331236 21968 331288
rect 22836 331236 22888 331288
rect 16304 331100 16356 331152
rect 134432 331236 134484 331288
rect 170496 331236 170548 331288
rect 171784 331236 171836 331288
rect 172336 331236 172388 331288
rect 173808 331236 173860 331288
rect 174912 331236 174964 331288
rect 290280 331236 290332 331288
rect 292672 331236 292724 331288
rect 301964 331236 302016 331288
rect 303068 331236 303120 331288
rect 352564 331236 352616 331288
rect 354036 331236 354088 331288
rect 404636 331236 404688 331288
rect 405740 331236 405792 331288
rect 465356 331236 465408 331288
rect 467104 331236 467156 331288
rect 160100 331168 160152 331220
rect 291384 331168 291436 331220
rect 293868 331168 293920 331220
rect 296720 331168 296772 331220
rect 394516 331168 394568 331220
rect 434996 331168 435048 331220
rect 565820 331168 565872 331220
rect 172336 331100 172388 331152
rect 285772 331100 285824 331152
rect 17684 331032 17736 331084
rect 119252 331032 119304 331084
rect 220820 331032 220872 331084
rect 292856 331032 292908 331084
rect 23388 330964 23440 331016
rect 99012 330964 99064 331016
rect 19156 330896 19208 330948
rect 154672 330896 154724 330948
rect 112444 330828 112496 330880
rect 114192 330828 114244 330880
rect 292856 330692 292908 330744
rect 294144 330692 294196 330744
rect 18972 330624 19024 330676
rect 19156 330624 19208 330676
rect 187608 330556 187660 330608
rect 285496 330556 285548 330608
rect 192116 330488 192168 330540
rect 291384 330488 291436 330540
rect 293960 330488 294012 330540
rect 303620 330488 303672 330540
rect 414756 330488 414808 330540
rect 565820 330488 565872 330540
rect 568856 330488 568908 330540
rect 572904 330488 572956 330540
rect 285496 329944 285548 329996
rect 286876 329944 286928 329996
rect 17592 329740 17644 329792
rect 17776 329740 17828 329792
rect 104072 329740 104124 329792
rect 294052 329740 294104 329792
rect 295340 329740 295392 329792
rect 296536 329740 296588 329792
rect 297732 329740 297784 329792
rect 299204 329740 299256 329792
rect 300768 329740 300820 329792
rect 301780 329740 301832 329792
rect 302148 329740 302200 329792
rect 302240 329740 302292 329792
rect 373908 329740 373960 329792
rect 440240 329740 440292 329792
rect 571616 329740 571668 329792
rect 19064 329672 19116 329724
rect 58532 329672 58584 329724
rect 343916 329672 343968 329724
rect 338856 329604 338908 329656
rect 299112 329536 299164 329588
rect 302240 329536 302292 329588
rect 195980 329060 196032 329112
rect 294052 329060 294104 329112
rect 297732 329060 297784 329112
rect 297916 329060 297968 329112
rect 399576 329060 399628 329112
rect 289084 319404 289136 319456
rect 424324 319404 424376 319456
rect 3332 318792 3384 318844
rect 10324 318792 10376 318844
rect 164240 318724 164292 318776
rect 284208 318724 284260 318776
rect 303068 318724 303120 318776
rect 303712 318724 303764 318776
rect 408500 318724 408552 318776
rect 449900 318724 449952 318776
rect 567660 318724 567712 318776
rect 459560 318656 459612 318708
rect 575480 318656 575532 318708
rect 489920 318588 489972 318640
rect 575572 318588 575624 318640
rect 304264 318044 304316 318096
rect 305184 318044 305236 318096
rect 405740 318044 405792 318096
rect 469220 318044 469272 318096
rect 573364 318044 573416 318096
rect 173808 317364 173860 317416
rect 285404 317364 285456 317416
rect 573364 317364 573416 317416
rect 574100 317364 574152 317416
rect 300584 316004 300636 316056
rect 306380 316004 306432 316056
rect 571524 316004 571576 316056
rect 16396 315936 16448 315988
rect 17224 315936 17276 315988
rect 112444 315936 112496 315988
rect 179420 315936 179472 315988
rect 285588 315936 285640 315988
rect 378140 315936 378192 315988
rect 505100 315936 505152 315988
rect 566372 315936 566424 315988
rect 567108 315936 567160 315988
rect 572812 315936 572864 315988
rect 22008 315868 22060 315920
rect 82820 315868 82872 315920
rect 215208 315868 215260 315920
rect 288532 315868 288584 315920
rect 296536 315868 296588 315920
rect 298008 315868 298060 315920
rect 368480 315868 368532 315920
rect 510620 315868 510672 315920
rect 570144 315868 570196 315920
rect 571524 315868 571576 315920
rect 20628 315800 20680 315852
rect 73160 315800 73212 315852
rect 224960 315800 225012 315852
rect 287520 315800 287572 315852
rect 303252 315800 303304 315852
rect 362960 315800 363012 315852
rect 514760 315800 514812 315852
rect 572720 315800 572772 315852
rect 234620 315732 234672 315784
rect 291200 315732 291252 315784
rect 298928 315732 298980 315784
rect 358820 315732 358872 315784
rect 520280 315732 520332 315784
rect 567752 315732 567804 315784
rect 299388 315664 299440 315716
rect 352564 315664 352616 315716
rect 525800 315664 525852 315716
rect 570052 315664 570104 315716
rect 300308 315596 300360 315648
rect 347780 315596 347832 315648
rect 529940 315596 529992 315648
rect 571524 315596 571576 315648
rect 285588 315392 285640 315444
rect 290096 315392 290148 315444
rect 276020 315324 276072 315376
rect 295984 315324 296036 315376
rect 18788 315188 18840 315240
rect 19340 315188 19392 315240
rect 93860 315256 93912 315308
rect 270500 315256 270552 315308
rect 297364 315256 297416 315308
rect 297824 314644 297876 314696
rect 298928 314644 298980 314696
rect 299112 314644 299164 314696
rect 300308 314644 300360 314696
rect 567752 314644 567804 314696
rect 568764 314644 568816 314696
rect 570144 314644 570196 314696
rect 571524 314644 571576 314696
rect 305000 314576 305052 314628
rect 389180 314576 389232 314628
rect 454040 314576 454092 314628
rect 565728 314576 565780 314628
rect 467104 314508 467156 314560
rect 568856 314508 568908 314560
rect 570328 314508 570380 314560
rect 565728 314168 565780 314220
rect 568856 314168 568908 314220
rect 285496 314032 285548 314084
rect 292764 314032 292816 314084
rect 284300 313964 284352 314016
rect 296720 313964 296772 314016
rect 200120 313896 200172 313948
rect 288624 313896 288676 313948
rect 296444 313896 296496 313948
rect 305092 313964 305144 314016
rect 301872 313896 301924 313948
rect 305000 313896 305052 313948
rect 300676 313828 300728 313880
rect 303620 313828 303672 313880
rect 3332 266364 3384 266416
rect 20904 266364 20956 266416
rect 2780 240184 2832 240236
rect 4896 240184 4948 240236
rect 12348 214548 12400 214600
rect 13176 214548 13228 214600
rect 3332 213936 3384 213988
rect 13268 213936 13320 213988
rect 296444 206252 296496 206304
rect 285496 205912 285548 205964
rect 288624 205912 288676 205964
rect 303620 205912 303672 205964
rect 568028 205640 568080 205692
rect 578240 205640 578292 205692
rect 285588 204892 285640 204944
rect 291384 204892 291436 204944
rect 293868 204892 293920 204944
rect 305092 204892 305144 204944
rect 526352 204892 526404 204944
rect 570052 204892 570104 204944
rect 572904 204892 572956 204944
rect 297824 204824 297876 204876
rect 301780 204824 301832 204876
rect 298008 204756 298060 204808
rect 299388 204756 299440 204808
rect 572720 204756 572772 204808
rect 574284 204756 574336 204808
rect 17500 204688 17552 204740
rect 18972 204688 19024 204740
rect 14832 204552 14884 204604
rect 180248 204552 180300 204604
rect 16304 204484 16356 204536
rect 18788 204484 18840 204536
rect 134432 204484 134484 204536
rect 17684 204416 17736 204468
rect 119252 204416 119304 204468
rect 18972 204348 19024 204400
rect 154672 204348 154724 204400
rect 246396 204552 246448 204604
rect 290188 204552 290240 204604
rect 292856 204552 292908 204604
rect 299388 204552 299440 204604
rect 354036 204552 354088 204604
rect 531504 204552 531556 204604
rect 572812 204552 572864 204604
rect 241336 204484 241388 204536
rect 289912 204484 289964 204536
rect 301780 204484 301832 204536
rect 359096 204484 359148 204536
rect 521660 204484 521712 204536
rect 567660 204484 567712 204536
rect 568764 204484 568816 204536
rect 235908 204416 235960 204468
rect 287888 204416 287940 204468
rect 291200 204416 291252 204468
rect 300584 204416 300636 204468
rect 303896 204416 303948 204468
rect 379336 204416 379388 204468
rect 515956 204416 516008 204468
rect 572720 204416 572772 204468
rect 220728 204348 220780 204400
rect 293960 204348 294012 204400
rect 290096 204280 290148 204332
rect 20444 204212 20496 204264
rect 20628 204212 20680 204264
rect 18880 204144 18932 204196
rect 88892 204212 88944 204264
rect 144828 204212 144880 204264
rect 149612 204212 149664 204264
rect 173900 204212 173952 204264
rect 175188 204212 175240 204264
rect 251088 204212 251140 204264
rect 22008 204144 22060 204196
rect 83832 204144 83884 204196
rect 256516 204144 256568 204196
rect 285680 204144 285732 204196
rect 20352 204076 20404 204128
rect 78772 204076 78824 204128
rect 190368 204076 190420 204128
rect 192484 204076 192536 204128
rect 291200 204212 291252 204264
rect 292580 204212 292632 204264
rect 299020 204212 299072 204264
rect 299296 204212 299348 204264
rect 299388 204212 299440 204264
rect 300768 204348 300820 204400
rect 301872 204348 301924 204400
rect 305000 204348 305052 204400
rect 389456 204348 389508 204400
rect 510896 204348 510948 204400
rect 571524 204348 571576 204400
rect 302884 204280 302936 204332
rect 505836 204280 505888 204332
rect 567476 204280 567528 204332
rect 567752 204280 567804 204332
rect 291384 204144 291436 204196
rect 292672 204144 292724 204196
rect 300768 204212 300820 204264
rect 302148 204212 302200 204264
rect 343916 204212 343968 204264
rect 404636 204212 404688 204264
rect 405924 204212 405976 204264
rect 424324 204212 424376 204264
rect 424876 204212 424928 204264
rect 429936 204212 429988 204264
rect 541256 204212 541308 204264
rect 567568 204212 567620 204264
rect 333796 204144 333848 204196
rect 546316 204144 546368 204196
rect 568672 204144 568724 204196
rect 289820 204076 289872 204128
rect 294052 204076 294104 204128
rect 299296 204076 299348 204128
rect 328736 204076 328788 204128
rect 382280 204076 382332 204128
rect 384396 204076 384448 204128
rect 470416 204076 470468 204128
rect 471336 204076 471388 204128
rect 561496 204076 561548 204128
rect 570236 204076 570288 204128
rect 20444 204008 20496 204060
rect 73712 204008 73764 204060
rect 303160 204008 303212 204060
rect 323676 204008 323728 204060
rect 4804 203940 4856 203992
rect 19064 203872 19116 203924
rect 20352 203872 20404 203924
rect 23296 203940 23348 203992
rect 33232 203940 33284 203992
rect 33324 203940 33376 203992
rect 38292 203940 38344 203992
rect 301964 203940 302016 203992
rect 318616 203940 318668 203992
rect 23388 203872 23440 203924
rect 281448 203872 281500 203924
rect 287704 203872 287756 203924
rect 291292 203872 291344 203924
rect 302056 203872 302108 203924
rect 313556 203872 313608 203924
rect 286784 203736 286836 203788
rect 293224 203736 293276 203788
rect 266268 203668 266320 203720
rect 291384 203668 291436 203720
rect 261576 203600 261628 203652
rect 291200 203600 291252 203652
rect 556436 203600 556488 203652
rect 568764 203600 568816 203652
rect 20352 203532 20404 203584
rect 58532 203532 58584 203584
rect 149612 203532 149664 203584
rect 289820 203532 289872 203584
rect 551376 203532 551428 203584
rect 570052 203532 570104 203584
rect 96620 203464 96672 203516
rect 99012 203464 99064 203516
rect 566556 203396 566608 203448
rect 568856 203396 568908 203448
rect 465356 203192 465408 203244
rect 467748 203192 467800 203244
rect 170496 203056 170548 203108
rect 171140 203056 171192 203108
rect 500776 203056 500828 203108
rect 503628 203056 503680 203108
rect 103520 202852 103572 202904
rect 165436 202852 165488 202904
rect 166264 202852 166316 202904
rect 413560 202852 413612 202904
rect 414756 202852 414808 202904
rect 440056 202852 440108 202904
rect 440884 202852 440936 202904
rect 445116 202852 445168 202904
rect 446404 202852 446456 202904
rect 495716 202852 495768 202904
rect 498568 202852 498620 202904
rect 21916 202784 21968 202836
rect 23112 202784 23164 202836
rect 23388 202784 23440 202836
rect 63592 202784 63644 202836
rect 104072 202784 104124 202836
rect 296720 202784 296772 202836
rect 303620 202784 303672 202836
rect 419540 202784 419592 202836
rect 22928 202716 22980 202768
rect 53472 202716 53524 202768
rect 175280 202716 175332 202768
rect 285772 202716 285824 202768
rect 303804 202716 303856 202768
rect 408500 202716 408552 202768
rect 409696 202716 409748 202768
rect 21824 202648 21876 202700
rect 48412 202648 48464 202700
rect 195796 202648 195848 202700
rect 284944 202648 284996 202700
rect 21732 202580 21784 202632
rect 23388 202580 23440 202632
rect 226156 202580 226208 202632
rect 287520 202580 287572 202632
rect 23112 202172 23164 202224
rect 33324 202172 33376 202224
rect 455236 202172 455288 202224
rect 564348 202172 564400 202224
rect 405924 202104 405976 202156
rect 560944 202104 560996 202156
rect 185308 201424 185360 201476
rect 292764 201424 292816 201476
rect 300676 201424 300728 201476
rect 413284 201424 413336 201476
rect 413560 201424 413612 201476
rect 467748 201424 467800 201476
rect 570328 201424 570380 201476
rect 572720 201424 572772 201476
rect 573364 201424 573416 201476
rect 574376 201424 574428 201476
rect 575480 201424 575532 201476
rect 216036 201356 216088 201408
rect 288532 201356 288584 201408
rect 296444 201356 296496 201408
rect 299204 201356 299256 201408
rect 338856 201356 338908 201408
rect 471336 201356 471388 201408
rect 231216 201288 231268 201340
rect 476120 201288 476172 201340
rect 575756 201288 575808 201340
rect 291568 201220 291620 201272
rect 292672 201220 292724 201272
rect 498568 201220 498620 201272
rect 574100 201220 574152 201272
rect 503628 201152 503680 201204
rect 574468 201152 574520 201204
rect 574468 201016 574520 201068
rect 575940 201016 575992 201068
rect 299204 200812 299256 200864
rect 374276 200812 374328 200864
rect 24124 200744 24176 200796
rect 185308 200744 185360 200796
rect 210976 200744 211028 200796
rect 285680 200744 285732 200796
rect 296628 200744 296680 200796
rect 302240 200744 302292 200796
rect 382280 200744 382332 200796
rect 460296 200744 460348 200796
rect 574376 200744 574428 200796
rect 285680 200132 285732 200184
rect 286876 200132 286928 200184
rect 287612 200132 287664 200184
rect 23572 200064 23624 200116
rect 158720 200064 158772 200116
rect 15016 199996 15068 200048
rect 139400 199996 139452 200048
rect 15108 199928 15160 199980
rect 17132 199928 17184 199980
rect 128360 199928 128412 199980
rect 17776 199860 17828 199912
rect 103428 199860 103480 199912
rect 14924 199452 14976 199504
rect 23572 199452 23624 199504
rect 22008 199384 22060 199436
rect 109040 199384 109092 199436
rect 20536 199044 20588 199096
rect 22008 199044 22060 199096
rect 17592 198704 17644 198756
rect 17776 198704 17828 198756
rect 440884 198636 440936 198688
rect 571616 198636 571668 198688
rect 446404 198568 446456 198620
rect 575664 198568 575716 198620
rect 20536 197956 20588 198008
rect 166264 197956 166316 198008
rect 408500 197956 408552 198008
rect 574192 197956 574244 198008
rect 287520 189728 287572 189780
rect 424324 189728 424376 189780
rect 23664 188980 23716 189032
rect 171140 188980 171192 189032
rect 434720 188980 434772 189032
rect 565728 188980 565780 189032
rect 16396 188912 16448 188964
rect 113180 188912 113232 188964
rect 489920 188912 489972 188964
rect 575572 188912 575624 188964
rect 565728 188368 565780 188420
rect 572996 188368 573048 188420
rect 296536 188300 296588 188352
rect 300676 188300 300728 188352
rect 368480 188300 368532 188352
rect 560944 188300 560996 188352
rect 578332 188300 578384 188352
rect 2780 187688 2832 187740
rect 4804 187688 4856 187740
rect 18972 187688 19024 187740
rect 23664 187688 23716 187740
rect 575572 187688 575624 187740
rect 575756 187688 575808 187740
rect 305736 187620 305788 187672
rect 398840 187620 398892 187672
rect 297824 187552 297876 187604
rect 305092 187552 305144 187604
rect 393320 187552 393372 187604
rect 303252 187484 303304 187536
rect 362960 187484 363012 187536
rect 296536 187144 296588 187196
rect 302240 187144 302292 187196
rect 285496 187008 285548 187060
rect 294144 187008 294196 187060
rect 276020 186940 276072 186992
rect 298744 186940 298796 186992
rect 299112 186940 299164 186992
rect 303344 186940 303396 186992
rect 347780 186940 347832 186992
rect 413284 186940 413336 186992
rect 579620 186940 579672 186992
rect 297916 186396 297968 186448
rect 303712 186396 303764 186448
rect 303068 186328 303120 186380
rect 303252 186328 303304 186380
rect 192484 186260 192536 186312
rect 285128 186260 285180 186312
rect 285588 186260 285640 186312
rect 17868 185920 17920 185972
rect 23020 185852 23072 185904
rect 24124 185852 24176 185904
rect 286876 185920 286928 185972
rect 292764 185920 292816 185972
rect 173900 185852 173952 185904
rect 200120 185852 200172 185904
rect 290096 185852 290148 185904
rect 300584 185852 300636 185904
rect 305000 185852 305052 185904
rect 419540 185852 419592 185904
rect 570236 185852 570288 185904
rect 2964 149064 3016 149116
rect 6368 149064 6420 149116
rect 2780 136688 2832 136740
rect 4988 136688 5040 136740
rect 3424 110440 3476 110492
rect 9036 110440 9088 110492
rect 2780 84328 2832 84380
rect 5080 84328 5132 84380
rect 574192 79296 574244 79348
rect 574468 79296 574520 79348
rect 16396 77936 16448 77988
rect 23020 77868 23072 77920
rect 25504 77868 25556 77920
rect 114192 77868 114244 77920
rect 193220 77868 193272 77920
rect 288532 78004 288584 78056
rect 300584 78004 300636 78056
rect 240784 77868 240836 77920
rect 290096 77936 290148 77988
rect 297824 77936 297876 77988
rect 284944 77868 284996 77920
rect 294144 77868 294196 77920
rect 332600 77868 332652 77920
rect 336004 77800 336056 77852
rect 20536 77052 20588 77104
rect 23480 77052 23532 77104
rect 299204 76712 299256 76764
rect 329104 76712 329156 76764
rect 293224 76644 293276 76696
rect 418160 76644 418212 76696
rect 430580 76644 430632 76696
rect 568856 76644 568908 76696
rect 222200 76576 222252 76628
rect 300124 76576 300176 76628
rect 301504 76576 301556 76628
rect 376760 76576 376812 76628
rect 404360 76576 404412 76628
rect 571432 76576 571484 76628
rect 153016 76508 153068 76560
rect 580264 76508 580316 76560
rect 13084 76100 13136 76152
rect 28172 76100 28224 76152
rect 17684 76032 17736 76084
rect 119896 76032 119948 76084
rect 219440 76032 219492 76084
rect 297180 76032 297232 76084
rect 18972 75964 19024 76016
rect 169760 75964 169812 76016
rect 200304 75964 200356 76016
rect 291476 75964 291528 76016
rect 385040 75964 385092 76016
rect 571432 75964 571484 76016
rect 18788 75896 18840 75948
rect 134432 75896 134484 75948
rect 153108 75896 153160 75948
rect 574192 75896 574244 75948
rect 19156 75828 19208 75880
rect 88984 75828 89036 75880
rect 144828 75828 144880 75880
rect 149612 75828 149664 75880
rect 149980 75828 150032 75880
rect 188344 75828 188396 75880
rect 190368 75828 190420 75880
rect 284300 75828 284352 75880
rect 301688 75828 301740 75880
rect 301964 75828 302016 75880
rect 318616 75828 318668 75880
rect 332600 75828 332652 75880
rect 389456 75828 389508 75880
rect 423680 75828 423732 75880
rect 424876 75828 424928 75880
rect 429936 75828 429988 75880
rect 505836 75828 505888 75880
rect 567752 75828 567804 75880
rect 20444 75760 20496 75812
rect 73804 75760 73856 75812
rect 216036 75760 216088 75812
rect 217324 75760 217376 75812
rect 261576 75760 261628 75812
rect 264888 75760 264940 75812
rect 511264 75760 511316 75812
rect 571524 75760 571576 75812
rect 20352 75692 20404 75744
rect 59268 75692 59320 75744
rect 515956 75692 516008 75744
rect 574284 75692 574336 75744
rect 21824 75624 21876 75676
rect 49056 75624 49108 75676
rect 520280 75624 520332 75676
rect 521016 75624 521068 75676
rect 567660 75624 567712 75676
rect 6184 75556 6236 75608
rect 23388 75556 23440 75608
rect 526076 75556 526128 75608
rect 572904 75556 572956 75608
rect 266268 75488 266320 75540
rect 270500 75488 270552 75540
rect 529940 75488 529992 75540
rect 531136 75488 531188 75540
rect 572812 75488 572864 75540
rect 241336 75420 241388 75472
rect 248420 75420 248472 75472
rect 251088 75420 251140 75472
rect 261484 75420 261536 75472
rect 286784 75420 286836 75472
rect 308404 75420 308456 75472
rect 246396 75352 246448 75404
rect 263600 75352 263652 75404
rect 292856 75352 292908 75404
rect 235908 75284 235960 75336
rect 240048 75284 240100 75336
rect 287888 75284 287940 75336
rect 319444 75284 319496 75336
rect 333796 75284 333848 75336
rect 49056 75148 49108 75200
rect 116584 75148 116636 75200
rect 191840 75148 191892 75200
rect 200396 75148 200448 75200
rect 226156 75148 226208 75200
rect 234436 75148 234488 75200
rect 231216 75080 231268 75132
rect 235908 75080 235960 75132
rect 292672 75216 292724 75268
rect 292856 75216 292908 75268
rect 301688 75216 301740 75268
rect 307944 75216 307996 75268
rect 323676 75216 323728 75268
rect 239496 75148 239548 75200
rect 515956 75148 516008 75200
rect 271696 74808 271748 74860
rect 276112 74808 276164 74860
rect 270500 74536 270552 74588
rect 271788 74536 271840 74588
rect 414020 74536 414072 74588
rect 414756 74536 414808 74588
rect 507032 74536 507084 74588
rect 19248 74468 19300 74520
rect 94320 74468 94372 74520
rect 256608 74468 256660 74520
rect 290004 74468 290056 74520
rect 302056 74468 302108 74520
rect 313280 74468 313332 74520
rect 536104 74468 536156 74520
rect 568580 74468 568632 74520
rect 20628 74400 20680 74452
rect 68284 74400 68336 74452
rect 271788 74400 271840 74452
rect 291384 74400 291436 74452
rect 303160 74400 303212 74452
rect 307852 74400 307904 74452
rect 541256 74400 541308 74452
rect 567568 74400 567620 74452
rect 21732 74332 21784 74384
rect 64144 74332 64196 74384
rect 281448 74332 281500 74384
rect 291292 74332 291344 74384
rect 545764 74332 545816 74384
rect 568672 74332 568724 74384
rect 23204 74264 23256 74316
rect 43444 74264 43496 74316
rect 560944 74264 560996 74316
rect 570144 74264 570196 74316
rect 23112 74196 23164 74248
rect 37924 74196 37976 74248
rect 23296 74128 23348 74180
rect 33692 74128 33744 74180
rect 342352 73992 342404 74044
rect 414020 73992 414072 74044
rect 79416 73924 79468 73976
rect 322204 73924 322256 73976
rect 322296 73924 322348 73976
rect 359096 73924 359148 73976
rect 408592 73924 408644 73976
rect 568764 73924 568816 73976
rect 119896 73856 119948 73908
rect 366272 73856 366324 73908
rect 390560 73856 390612 73908
rect 570052 73856 570104 73908
rect 226432 73788 226484 73840
rect 485596 73788 485648 73840
rect 507032 73788 507084 73840
rect 534080 73788 534132 73840
rect 14832 73108 14884 73160
rect 180064 73108 180116 73160
rect 301872 73108 301924 73160
rect 322112 73108 322164 73160
rect 322296 73108 322348 73160
rect 435364 73108 435416 73160
rect 572996 73108 573048 73160
rect 17868 73040 17920 73092
rect 174544 73040 174596 73092
rect 445024 73040 445076 73092
rect 575664 73040 575716 73092
rect 14924 72972 14976 73024
rect 159364 72972 159416 73024
rect 450544 72972 450596 73024
rect 578240 72972 578292 73024
rect 23480 72904 23532 72956
rect 164240 72904 164292 72956
rect 459560 72904 459612 72956
rect 460296 72904 460348 72956
rect 574376 72904 574428 72956
rect 17500 72836 17552 72888
rect 155224 72836 155276 72888
rect 490564 72836 490616 72888
rect 575756 72836 575808 72888
rect 534080 72768 534132 72820
rect 579620 72768 579672 72820
rect 211712 72632 211764 72684
rect 288624 72632 288676 72684
rect 134432 72564 134484 72616
rect 371792 72564 371844 72616
rect 254032 72496 254084 72548
rect 529940 72496 529992 72548
rect 164240 72428 164292 72480
rect 164792 72428 164844 72480
rect 169852 72428 169904 72480
rect 459560 72428 459612 72480
rect 15016 71680 15068 71732
rect 140044 71680 140096 71732
rect 439596 71680 439648 71732
rect 571616 71680 571668 71732
rect 25596 71612 25648 71664
rect 124588 71612 124640 71664
rect 125508 71612 125560 71664
rect 469864 71612 469916 71664
rect 470416 71612 470468 71664
rect 572720 71612 572772 71664
rect 22008 71544 22060 71596
rect 109132 71544 109184 71596
rect 475384 71544 475436 71596
rect 575848 71544 575900 71596
rect 496084 71476 496136 71528
rect 574100 71476 574152 71528
rect 500776 71408 500828 71460
rect 575940 71408 575992 71460
rect 262128 71340 262180 71392
rect 289912 71340 289964 71392
rect 239404 71272 239456 71324
rect 292764 71272 292816 71324
rect 248420 71204 248472 71256
rect 261392 71204 261444 71256
rect 262128 71204 262180 71256
rect 288992 71204 289044 71256
rect 423680 71204 423732 71256
rect 114468 71136 114520 71188
rect 364432 71136 364484 71188
rect 94320 71068 94372 71120
rect 357440 71068 357492 71120
rect 33692 71000 33744 71052
rect 303712 71000 303764 71052
rect 331220 71000 331272 71052
rect 384396 71000 384448 71052
rect 109132 70388 109184 70440
rect 109684 70388 109736 70440
rect 296536 70320 296588 70372
rect 331220 70320 331272 70372
rect 405648 70320 405700 70372
rect 578332 70320 578384 70372
rect 237472 69912 237524 69964
rect 239496 69912 239548 69964
rect 264888 69844 264940 69896
rect 269120 69844 269172 69896
rect 291200 69844 291252 69896
rect 317328 69844 317380 69896
rect 343916 69844 343968 69896
rect 125508 69776 125560 69828
rect 368480 69776 368532 69828
rect 59268 69708 59320 69760
rect 313372 69708 313424 69760
rect 338120 69708 338172 69760
rect 404452 69708 404504 69760
rect 405648 69708 405700 69760
rect 410432 69708 410484 69760
rect 556436 69708 556488 69760
rect 12348 69640 12400 69692
rect 40684 69640 40736 69692
rect 252560 69640 252612 69692
rect 526076 69640 526128 69692
rect 25504 68960 25556 69012
rect 184940 68960 184992 69012
rect 300768 68960 300820 69012
rect 316592 68960 316644 69012
rect 317328 68960 317380 69012
rect 409144 68960 409196 69012
rect 574468 68960 574520 69012
rect 195152 68552 195204 68604
rect 284944 68552 284996 68604
rect 149980 68484 150032 68536
rect 272432 68484 272484 68536
rect 276112 68484 276164 68536
rect 375472 68484 375524 68536
rect 265624 68416 265676 68468
rect 520280 68416 520332 68468
rect 84108 68348 84160 68400
rect 353392 68348 353444 68400
rect 234436 68280 234488 68332
rect 244832 68280 244884 68332
rect 258080 68280 258132 68332
rect 541256 68280 541308 68332
rect 217324 67532 217376 67584
rect 240784 67532 240836 67584
rect 244832 67532 244884 67584
rect 287796 67532 287848 67584
rect 336004 67532 336056 67584
rect 393320 67532 393372 67584
rect 261484 67464 261536 67516
rect 265072 67464 265124 67516
rect 265072 67056 265124 67108
rect 294052 67056 294104 67108
rect 231952 66988 232004 67040
rect 500776 66988 500828 67040
rect 73804 66920 73856 66972
rect 349712 66920 349764 66972
rect 255872 66852 255924 66904
rect 536104 66852 536156 66904
rect 335360 66784 335412 66836
rect 336004 66784 336056 66836
rect 219532 65628 219584 65680
rect 242992 65628 243044 65680
rect 271144 65628 271196 65680
rect 480260 65628 480312 65680
rect 228272 65560 228324 65612
rect 490564 65560 490616 65612
rect 187792 65492 187844 65544
rect 194600 65492 194652 65544
rect 209780 65492 209832 65544
rect 226984 65492 227036 65544
rect 230480 65492 230532 65544
rect 496084 65492 496136 65544
rect 242992 64948 243044 65000
rect 243820 64948 243872 65000
rect 243820 64812 243872 64864
rect 293960 64812 294012 64864
rect 40684 64268 40736 64320
rect 178684 64268 178736 64320
rect 206284 64268 206336 64320
rect 465724 64268 465776 64320
rect 173072 64200 173124 64252
rect 469864 64200 469916 64252
rect 175280 64132 175332 64184
rect 475384 64132 475436 64184
rect 297916 63044 297968 63096
rect 329840 63044 329892 63096
rect 303068 62976 303120 63028
rect 324320 62976 324372 63028
rect 362960 62976 363012 63028
rect 203524 62908 203576 62960
rect 445024 62908 445076 62960
rect 154672 62840 154724 62892
rect 435364 62840 435416 62892
rect 156512 62772 156564 62824
rect 439596 62772 439648 62824
rect 299296 62024 299348 62076
rect 328460 62024 328512 62076
rect 329104 62024 329156 62076
rect 374000 62024 374052 62076
rect 300676 61616 300728 61668
rect 325884 61616 325936 61668
rect 308404 61548 308456 61600
rect 415952 61548 416004 61600
rect 116584 61480 116636 61532
rect 309232 61480 309284 61532
rect 309784 61480 309836 61532
rect 338212 61480 338264 61532
rect 52460 61412 52512 61464
rect 311072 61412 311124 61464
rect 3516 61344 3568 61396
rect 13084 61344 13136 61396
rect 43444 61344 43496 61396
rect 307760 61344 307812 61396
rect 325884 61344 325936 61396
rect 368572 61344 368624 61396
rect 412640 61344 412692 61396
rect 560944 61344 560996 61396
rect 298836 60732 298888 60784
rect 299296 60732 299348 60784
rect 297456 60324 297508 60376
rect 313280 60324 313332 60376
rect 340880 60324 340932 60376
rect 409144 60324 409196 60376
rect 298744 60256 298796 60308
rect 396080 60256 396132 60308
rect 295984 60188 296036 60240
rect 397552 60188 397604 60240
rect 109684 60120 109736 60172
rect 362960 60120 363012 60172
rect 104164 60052 104216 60104
rect 360752 60052 360804 60104
rect 98644 59984 98696 60036
rect 358912 59984 358964 60036
rect 336740 59304 336792 59356
rect 398932 59304 398984 59356
rect 140044 58760 140096 58812
rect 374000 58760 374052 58812
rect 432512 58760 432564 58812
rect 565820 58760 565872 58812
rect 88984 58692 89036 58744
rect 355232 58692 355284 58744
rect 355324 58692 355376 58744
rect 511264 58692 511316 58744
rect 68284 58624 68336 58676
rect 347872 58624 347924 58676
rect 392032 58624 392084 58676
rect 550640 58624 550692 58676
rect 329840 57876 329892 57928
rect 378140 57876 378192 57928
rect 294604 57468 294656 57520
rect 383200 57468 383252 57520
rect 129004 57400 129056 57452
rect 370320 57400 370372 57452
rect 37924 57332 37976 57384
rect 305920 57332 305972 57384
rect 64144 57264 64196 57316
rect 346400 57264 346452 57316
rect 259920 57196 259972 57248
rect 545764 57196 545816 57248
rect 299388 56516 299440 56568
rect 319444 56516 319496 56568
rect 298560 56176 298612 56228
rect 299388 56176 299440 56228
rect 294880 56108 294932 56160
rect 307852 56108 307904 56160
rect 303252 56040 303304 56092
rect 318800 56108 318852 56160
rect 347780 56108 347832 56160
rect 320640 56040 320692 56092
rect 353300 56040 353352 56092
rect 169760 55972 169812 56024
rect 178960 55972 179012 56024
rect 235908 55972 235960 56024
rect 247040 55972 247092 56024
rect 256608 55972 256660 56024
rect 267280 55972 267332 56024
rect 281448 55972 281500 56024
rect 294604 55972 294656 56024
rect 298008 55972 298060 56024
rect 344560 55972 344612 56024
rect 420184 55972 420236 56024
rect 166080 55904 166132 55956
rect 450544 55904 450596 55956
rect 167920 55836 167972 55888
rect 454040 55836 454092 55888
rect 226984 55156 227036 55208
rect 239404 55156 239456 55208
rect 278320 54816 278372 54868
rect 288440 54816 288492 54868
rect 296444 54816 296496 54868
rect 178684 54748 178736 54800
rect 174544 54680 174596 54732
rect 180800 54680 180852 54732
rect 180064 54612 180116 54664
rect 182640 54612 182692 54664
rect 282000 54748 282052 54800
rect 287612 54748 287664 54800
rect 297364 54748 297416 54800
rect 240048 54680 240100 54732
rect 248880 54680 248932 54732
rect 250720 54680 250772 54732
rect 265624 54680 265676 54732
rect 274640 54680 274692 54732
rect 289820 54680 289872 54732
rect 291200 54680 291252 54732
rect 297456 54680 297508 54732
rect 300400 54748 300452 54800
rect 309784 54748 309836 54800
rect 322204 54748 322256 54800
rect 351920 54748 351972 54800
rect 379520 54680 379572 54732
rect 197360 54612 197412 54664
rect 208400 54612 208452 54664
rect 271144 54612 271196 54664
rect 276020 54612 276072 54664
rect 394240 54612 394292 54664
rect 171600 54544 171652 54596
rect 206284 54544 206336 54596
rect 236000 54544 236052 54596
rect 355324 54544 355376 54596
rect 429200 54544 429252 54596
rect 439504 54544 439556 54596
rect 158720 54476 158772 54528
rect 203524 54476 203576 54528
rect 204260 54476 204312 54528
rect 210240 54476 210292 54528
rect 159364 54408 159416 54460
rect 162400 54408 162452 54460
rect 206560 54408 206612 54460
rect 282276 54476 282328 54528
rect 294604 54476 294656 54528
rect 414480 54476 414532 54528
rect 427360 54476 427412 54528
rect 558184 54476 558236 54528
rect 285680 54272 285732 54324
rect 289084 54272 289136 54324
rect 240784 53864 240836 53916
rect 241520 53864 241572 53916
rect 155224 53796 155276 53848
rect 160560 53796 160612 53848
rect 186320 53796 186372 53848
rect 188344 53796 188396 53848
rect 221280 53796 221332 53848
rect 285772 53796 285824 53848
rect 296720 53796 296772 53848
rect 298836 53796 298888 53848
rect 328000 53796 328052 53848
rect 329104 53796 329156 53848
rect 13268 53048 13320 53100
rect 151084 53048 151136 53100
rect 151544 53048 151596 53100
rect 577504 53048 577556 53100
rect 4988 51008 5040 51060
rect 150440 51008 150492 51060
rect 6368 49648 6420 49700
rect 150440 49648 150492 49700
rect 4896 48220 4948 48272
rect 150440 48220 150492 48272
rect 21364 48152 21416 48204
rect 150532 48152 150584 48204
rect 4804 46860 4856 46912
rect 150440 46860 150492 46912
rect 13084 45500 13136 45552
rect 150440 45500 150492 45552
rect 10324 44072 10376 44124
rect 150440 44072 150492 44124
rect 8944 42712 8996 42764
rect 150440 42712 150492 42764
rect 6276 41352 6328 41404
rect 150440 41352 150492 41404
rect 7564 39312 7616 39364
rect 151176 39312 151228 39364
rect 437388 37272 437440 37324
rect 565084 37272 565136 37324
rect 9036 36524 9088 36576
rect 151084 36524 151136 36576
rect 16488 35844 16540 35896
rect 150440 35844 150492 35896
rect 15844 34416 15896 34468
rect 150440 34416 150492 34468
rect 7656 33056 7708 33108
rect 150440 33056 150492 33108
rect 3516 31696 3568 31748
rect 150440 31696 150492 31748
rect 3424 30268 3476 30320
rect 150440 30268 150492 30320
rect 5080 28908 5132 28960
rect 150440 28908 150492 28960
rect 3608 26188 3660 26240
rect 150440 26188 150492 26240
rect 214840 23740 214892 23792
rect 299664 23740 299716 23792
rect 244096 23672 244148 23724
rect 336004 23672 336056 23724
rect 266268 23604 266320 23656
rect 480260 23604 480312 23656
rect 267372 23536 267424 23588
rect 483020 23536 483072 23588
rect 269488 23468 269540 23520
rect 489920 23468 489972 23520
rect 215484 22448 215536 22500
rect 301412 22448 301464 22500
rect 217508 22380 217560 22432
rect 309232 22380 309284 22432
rect 220544 22312 220596 22364
rect 320272 22312 320324 22364
rect 228640 22244 228692 22296
rect 349252 22244 349304 22296
rect 241796 22176 241848 22228
rect 394700 22176 394752 22228
rect 275192 22108 275244 22160
rect 512000 22108 512052 22160
rect 297364 21836 297416 21888
rect 291844 21768 291896 21820
rect 250904 21700 250956 21752
rect 276020 21700 276072 21752
rect 278688 21700 278740 21752
rect 297456 21700 297508 21752
rect 226616 21632 226668 21684
rect 246304 21632 246356 21684
rect 254032 21632 254084 21684
rect 383476 21768 383528 21820
rect 388444 21768 388496 21820
rect 307576 21700 307628 21752
rect 315304 21700 315356 21752
rect 322756 21700 322808 21752
rect 350632 21700 350684 21752
rect 358176 21700 358228 21752
rect 385500 21700 385552 21752
rect 394608 21700 394660 21752
rect 398656 21700 398708 21752
rect 437572 21700 437624 21752
rect 230664 21564 230716 21616
rect 262864 21564 262916 21616
rect 298468 21564 298520 21616
rect 323584 21632 323636 21684
rect 342996 21632 343048 21684
rect 369308 21632 369360 21684
rect 371148 21632 371200 21684
rect 386512 21632 386564 21684
rect 426808 21632 426860 21684
rect 338948 21564 339000 21616
rect 342904 21564 342956 21616
rect 354128 21564 354180 21616
rect 388536 21564 388588 21616
rect 440240 21564 440292 21616
rect 164332 21496 164384 21548
rect 176016 21496 176068 21548
rect 193220 21496 193272 21548
rect 210332 21496 210384 21548
rect 211436 21496 211488 21548
rect 249984 21496 250036 21548
rect 263048 21496 263100 21548
rect 278136 21496 278188 21548
rect 279424 21496 279476 21548
rect 199292 21428 199344 21480
rect 228364 21428 228416 21480
rect 242164 21428 242216 21480
rect 301504 21428 301556 21480
rect 304264 21428 304316 21480
rect 312636 21428 312688 21480
rect 127624 21360 127676 21412
rect 164884 21360 164936 21412
rect 206284 21360 206336 21412
rect 303528 21360 303580 21412
rect 302884 21292 302936 21344
rect 311624 21360 311676 21412
rect 311164 21292 311216 21344
rect 316684 21292 316736 21344
rect 320824 21496 320876 21548
rect 333980 21496 334032 21548
rect 340972 21496 341024 21548
rect 343640 21496 343692 21548
rect 356152 21496 356204 21548
rect 371332 21496 371384 21548
rect 377496 21496 377548 21548
rect 381452 21496 381504 21548
rect 387064 21496 387116 21548
rect 392584 21496 392636 21548
rect 456892 21496 456944 21548
rect 345020 21428 345072 21480
rect 390560 21428 390612 21480
rect 465080 21428 465132 21480
rect 334900 21360 334952 21412
rect 325700 21292 325752 21344
rect 351092 21360 351144 21412
rect 368296 21360 368348 21412
rect 378784 21360 378836 21412
rect 394516 21360 394568 21412
rect 478880 21360 478932 21412
rect 312544 21224 312596 21276
rect 319720 21224 319772 21276
rect 309784 21156 309836 21208
rect 318708 21156 318760 21208
rect 322756 21156 322808 21208
rect 325792 21156 325844 21208
rect 300952 21088 301004 21140
rect 306564 21088 306616 21140
rect 375380 21020 375432 21072
rect 382924 21020 382976 21072
rect 306564 20952 306616 21004
rect 308588 20952 308640 21004
rect 347780 20952 347832 21004
rect 357164 20952 357216 21004
rect 363236 20952 363288 21004
rect 366364 20952 366416 21004
rect 174544 20884 174596 20936
rect 178040 20884 178092 20936
rect 184112 20816 184164 20868
rect 185584 20816 185636 20868
rect 234712 20816 234764 20868
rect 240784 20816 240836 20868
rect 380440 20816 380492 20868
rect 384396 20816 384448 20868
rect 178040 20748 178092 20800
rect 180064 20748 180116 20800
rect 182088 20748 182140 20800
rect 184204 20748 184256 20800
rect 317052 20748 317104 20800
rect 323768 20748 323820 20800
rect 366272 20748 366324 20800
rect 367744 20748 367796 20800
rect 171784 20680 171836 20732
rect 177028 20680 177080 20732
rect 177304 20680 177356 20732
rect 179052 20680 179104 20732
rect 181076 20680 181128 20732
rect 182180 20680 182232 20732
rect 183100 20680 183152 20732
rect 184296 20680 184348 20732
rect 210424 20680 210476 20732
rect 211804 20680 211856 20732
rect 298744 20680 298796 20732
rect 304540 20680 304592 20732
rect 307116 20680 307168 20732
rect 309600 20680 309652 20732
rect 311256 20680 311308 20732
rect 314660 20680 314712 20732
rect 318064 20680 318116 20732
rect 320732 20680 320784 20732
rect 356704 20680 356756 20732
rect 359188 20680 359240 20732
rect 359464 20680 359516 20732
rect 360200 20680 360252 20732
rect 362224 20680 362276 20732
rect 363604 20680 363656 20732
rect 365260 20680 365312 20732
rect 366456 20680 366508 20732
rect 378416 20680 378468 20732
rect 380164 20680 380216 20732
rect 384488 20680 384540 20732
rect 392584 20680 392636 20732
rect 249984 20340 250036 20392
rect 288440 20340 288492 20392
rect 301596 20340 301648 20392
rect 331864 20340 331916 20392
rect 237380 20272 237432 20324
rect 322756 20272 322808 20324
rect 201500 20204 201552 20256
rect 315672 20204 315724 20256
rect 334624 20204 334676 20256
rect 350080 20204 350132 20256
rect 394608 20204 394660 20256
rect 447140 20204 447192 20256
rect 176660 20136 176712 20188
rect 306564 20136 306616 20188
rect 330484 20136 330536 20188
rect 347044 20136 347096 20188
rect 378784 20136 378836 20188
rect 386420 20136 386472 20188
rect 396632 20136 396684 20188
rect 485780 20136 485832 20188
rect 169760 20068 169812 20120
rect 300952 20068 301004 20120
rect 319444 20068 319496 20120
rect 339960 20068 340012 20120
rect 371148 20068 371200 20120
rect 390744 20068 390796 20120
rect 397644 20068 397696 20120
rect 490012 20068 490064 20120
rect 138020 20000 138072 20052
rect 278688 20000 278740 20052
rect 291200 20000 291252 20052
rect 333980 20000 334032 20052
rect 367284 20000 367336 20052
rect 382280 20000 382332 20052
rect 382924 20000 382976 20052
rect 411260 20000 411312 20052
rect 411812 20000 411864 20052
rect 539600 20000 539652 20052
rect 165620 19932 165672 19984
rect 166540 19932 166592 19984
rect 169852 19932 169904 19984
rect 170588 19932 170640 19984
rect 173900 19932 173952 19984
rect 174636 19932 174688 19984
rect 189080 19932 189132 19984
rect 189908 19932 189960 19984
rect 195980 19932 196032 19984
rect 196900 19932 196952 19984
rect 208400 19932 208452 19984
rect 209044 19932 209096 19984
rect 245752 19932 245804 19984
rect 246580 19932 246632 19984
rect 271880 19932 271932 19984
rect 272892 19932 272944 19984
rect 278136 19932 278188 19984
rect 469220 19932 469272 19984
rect 287060 19864 287112 19916
rect 287980 19864 288032 19916
rect 332600 19864 332652 19916
rect 333612 19864 333664 19916
rect 336740 19864 336792 19916
rect 337660 19864 337712 19916
rect 401600 19864 401652 19916
rect 402428 19864 402480 19916
rect 408592 19864 408644 19916
rect 409420 19864 409472 19916
rect 412732 19864 412784 19916
rect 413468 19864 413520 19916
rect 389548 19524 389600 19576
rect 393964 19524 394016 19576
rect 185216 18912 185268 18964
rect 310612 18912 310664 18964
rect 420920 18912 420972 18964
rect 421564 18912 421616 18964
rect 135260 18844 135312 18896
rect 296444 18844 296496 18896
rect 298100 18844 298152 18896
rect 323584 18844 323636 18896
rect 257988 18776 258040 18828
rect 451280 18776 451332 18828
rect 259000 18708 259052 18760
rect 455420 18708 455472 18760
rect 202328 18640 202380 18692
rect 256700 18640 256752 18692
rect 260012 18640 260064 18692
rect 458180 18640 458232 18692
rect 203340 18572 203392 18624
rect 259460 18572 259512 18624
rect 261024 18572 261076 18624
rect 462320 18572 462372 18624
rect 230480 17552 230532 17604
rect 317052 17552 317104 17604
rect 142160 17484 142212 17536
rect 254032 17484 254084 17536
rect 276020 17484 276072 17536
rect 426440 17484 426492 17536
rect 426808 17484 426860 17536
rect 449900 17484 449952 17536
rect 131120 17416 131172 17468
rect 295432 17416 295484 17468
rect 416872 17416 416924 17468
rect 556160 17416 556212 17468
rect 251916 17348 251968 17400
rect 430580 17348 430632 17400
rect 198280 17280 198332 17332
rect 242900 17280 242952 17332
rect 252928 17280 252980 17332
rect 433340 17280 433392 17332
rect 440240 17280 440292 17332
rect 456800 17280 456852 17332
rect 456892 17280 456944 17332
rect 471980 17280 472032 17332
rect 201316 17212 201368 17264
rect 252560 17212 252612 17264
rect 253940 17212 253992 17264
rect 437480 17212 437532 17264
rect 437572 17212 437624 17264
rect 492680 17212 492732 17264
rect 204260 16668 204312 16720
rect 204996 16668 205048 16720
rect 145472 16192 145524 16244
rect 247684 16192 247736 16244
rect 273904 16192 273956 16244
rect 305000 16192 305052 16244
rect 307024 16192 307076 16244
rect 329932 16192 329984 16244
rect 401692 16192 401744 16244
rect 503720 16192 503772 16244
rect 198740 16124 198792 16176
rect 311256 16124 311308 16176
rect 402980 16124 403032 16176
rect 511264 16124 511316 16176
rect 244280 16056 244332 16108
rect 406016 16056 406068 16108
rect 228364 15988 228416 16040
rect 196072 15920 196124 15972
rect 234620 15920 234672 15972
rect 200120 15852 200172 15904
rect 244924 15852 244976 15904
rect 245844 15988 245896 16040
rect 409144 16056 409196 16108
rect 408684 15988 408736 16040
rect 528560 15988 528612 16040
rect 245752 15920 245804 15972
rect 412640 15920 412692 15972
rect 412824 15920 412876 15972
rect 542728 15920 542780 15972
rect 245936 15852 245988 15904
rect 247040 15852 247092 15904
rect 415400 15852 415452 15904
rect 260104 14764 260156 14816
rect 330392 14764 330444 14816
rect 380164 14764 380216 14816
rect 422576 14764 422628 14816
rect 213368 14696 213420 14748
rect 309784 14696 309836 14748
rect 384396 14696 384448 14748
rect 429200 14696 429252 14748
rect 236000 14628 236052 14680
rect 347044 14628 347096 14680
rect 388444 14628 388496 14680
rect 440332 14628 440384 14680
rect 190460 14560 190512 14612
rect 218060 14560 218112 14612
rect 237472 14560 237524 14612
rect 370504 14560 370556 14612
rect 376760 14560 376812 14612
rect 418528 14560 418580 14612
rect 419540 14560 419592 14612
rect 567568 14560 567620 14612
rect 194600 14492 194652 14544
rect 231860 14492 231912 14544
rect 238852 14492 238904 14544
rect 377404 14492 377456 14544
rect 421012 14492 421064 14544
rect 571340 14492 571392 14544
rect 195980 14424 196032 14476
rect 238944 14424 238996 14476
rect 381544 14424 381596 14476
rect 420920 14424 420972 14476
rect 575112 14424 575164 14476
rect 239312 14356 239364 14408
rect 262864 13404 262916 13456
rect 356336 13404 356388 13456
rect 219992 13336 220044 13388
rect 318064 13336 318116 13388
rect 378692 13336 378744 13388
rect 425704 13336 425756 13388
rect 229100 13268 229152 13320
rect 337384 13268 337436 13320
rect 381728 13268 381780 13320
rect 515496 13268 515548 13320
rect 230848 13200 230900 13252
rect 359372 13200 359424 13252
rect 375472 13200 375524 13252
rect 231952 13132 232004 13184
rect 363420 13132 363472 13184
rect 369860 13132 369912 13184
rect 381636 13132 381688 13184
rect 193312 13064 193364 13116
rect 228272 13064 228324 13116
rect 233240 13064 233292 13116
rect 365812 13064 365864 13116
rect 366456 13064 366508 13116
rect 376024 13064 376076 13116
rect 412732 13200 412784 13252
rect 546500 13200 546552 13252
rect 386696 13132 386748 13184
rect 413284 13132 413336 13184
rect 414020 13132 414072 13184
rect 550272 13132 550324 13184
rect 415492 13064 415544 13116
rect 415584 13064 415636 13116
rect 553768 13064 553820 13116
rect 276664 12044 276716 12096
rect 336832 12044 336884 12096
rect 210332 11976 210384 12028
rect 225144 11976 225196 12028
rect 227536 11976 227588 12028
rect 315304 11976 315356 12028
rect 387064 11976 387116 12028
rect 431960 11976 432012 12028
rect 151820 11908 151872 11960
rect 242164 11908 242216 11960
rect 246304 11908 246356 11960
rect 340972 11908 341024 11960
rect 405832 11908 405884 11960
rect 494796 11908 494848 11960
rect 223580 11840 223632 11892
rect 331220 11840 331272 11892
rect 405924 11840 405976 11892
rect 521660 11840 521712 11892
rect 189172 11772 189224 11824
rect 209780 11772 209832 11824
rect 223672 11772 223724 11824
rect 334624 11772 334676 11824
rect 337476 11772 337528 11824
rect 352196 11772 352248 11824
rect 372712 11772 372764 11824
rect 404452 11772 404504 11824
rect 407212 11772 407264 11824
rect 525432 11772 525484 11824
rect 157800 11704 157852 11756
rect 173992 11704 174044 11756
rect 189080 11704 189132 11756
rect 214472 11704 214524 11756
rect 225052 11704 225104 11756
rect 338672 11704 338724 11756
rect 338764 11704 338816 11756
rect 351920 11704 351972 11756
rect 363512 11704 363564 11756
rect 372896 11704 372948 11756
rect 374000 11704 374052 11756
rect 407120 11704 407172 11756
rect 408592 11704 408644 11756
rect 532056 11704 532108 11756
rect 393320 10956 393372 11008
rect 399484 10956 399536 11008
rect 280712 10616 280764 10668
rect 336740 10616 336792 10668
rect 262496 10548 262548 10600
rect 332692 10548 332744 10600
rect 382372 10548 382424 10600
rect 436744 10548 436796 10600
rect 191840 10480 191892 10532
rect 221096 10480 221148 10532
rect 241704 10480 241756 10532
rect 325884 10480 325936 10532
rect 398840 10480 398892 10532
rect 497096 10480 497148 10532
rect 218152 10412 218204 10464
rect 305644 10412 305696 10464
rect 330576 10412 330628 10464
rect 345112 10412 345164 10464
rect 345664 10412 345716 10464
rect 354680 10412 354732 10464
rect 367744 10412 367796 10464
rect 379520 10412 379572 10464
rect 400220 10412 400272 10464
rect 500592 10412 500644 10464
rect 143540 10344 143592 10396
rect 169944 10344 169996 10396
rect 186320 10344 186372 10396
rect 203432 10344 203484 10396
rect 219532 10344 219584 10396
rect 316040 10344 316092 10396
rect 316684 10344 316736 10396
rect 335360 10344 335412 10396
rect 337568 10344 337620 10396
rect 348332 10344 348384 10396
rect 377496 10344 377548 10396
rect 397736 10344 397788 10396
rect 401600 10344 401652 10396
rect 507216 10344 507268 10396
rect 141424 10276 141476 10328
rect 168380 10276 168432 10328
rect 187700 10276 187752 10328
rect 207112 10276 207164 10328
rect 209872 10276 209924 10328
rect 317512 10276 317564 10328
rect 336096 10276 336148 10328
rect 347872 10276 347924 10328
rect 371516 10276 371568 10328
rect 400864 10276 400916 10328
rect 409880 10276 409932 10328
rect 536104 10276 536156 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 248788 9324 248840 9376
rect 328460 9324 328512 9376
rect 211620 9256 211672 9308
rect 292580 9256 292632 9308
rect 195612 9188 195664 9240
rect 313280 9188 313332 9240
rect 174268 9120 174320 9172
rect 297364 9120 297416 9172
rect 329656 9120 329708 9172
rect 343732 9120 343784 9172
rect 394792 9120 394844 9172
rect 482836 9120 482888 9172
rect 181444 9052 181496 9104
rect 307116 9052 307168 9104
rect 307760 9052 307812 9104
rect 332600 9052 332652 9104
rect 404360 9052 404412 9104
rect 514760 9052 514812 9104
rect 136456 8984 136508 9036
rect 167000 8984 167052 9036
rect 291292 8984 291344 9036
rect 555424 8984 555476 9036
rect 129372 8916 129424 8968
rect 165712 8916 165764 8968
rect 284392 8916 284444 8968
rect 291844 8916 291896 8968
rect 292672 8916 292724 8968
rect 576308 8916 576360 8968
rect 300492 8168 300544 8220
rect 302332 8168 302384 8220
rect 207020 7896 207072 7948
rect 274824 7896 274876 7948
rect 277492 7896 277544 7948
rect 299572 7896 299624 7948
rect 305552 7896 305604 7948
rect 320824 7896 320876 7948
rect 252468 7828 252520 7880
rect 324320 7828 324372 7880
rect 206192 7760 206244 7812
rect 311164 7760 311216 7812
rect 323584 7760 323636 7812
rect 341064 7760 341116 7812
rect 392584 7760 392636 7812
rect 443828 7760 443880 7812
rect 234896 7692 234948 7744
rect 348516 7692 348568 7744
rect 417056 7692 417108 7744
rect 560852 7692 560904 7744
rect 154212 7624 154264 7676
rect 172520 7624 172572 7676
rect 185032 7624 185084 7676
rect 196808 7624 196860 7676
rect 208492 7624 208544 7676
rect 278320 7624 278372 7676
rect 284484 7624 284536 7676
rect 547880 7624 547932 7676
rect 132960 7556 133012 7608
rect 165620 7556 165672 7608
rect 185124 7556 185176 7608
rect 200304 7556 200356 7608
rect 208400 7556 208452 7608
rect 281908 7556 281960 7608
rect 285680 7556 285732 7608
rect 551468 7556 551520 7608
rect 3424 6808 3476 6860
rect 151084 6808 151136 6860
rect 270040 6536 270092 6588
rect 279424 6536 279476 6588
rect 245200 6468 245252 6520
rect 327080 6468 327132 6520
rect 216864 6400 216916 6452
rect 312544 6400 312596 6452
rect 188528 6332 188580 6384
rect 302884 6332 302936 6384
rect 422300 6332 422352 6384
rect 468760 6332 468812 6384
rect 277400 6264 277452 6316
rect 523040 6264 523092 6316
rect 150624 6196 150676 6248
rect 171140 6196 171192 6248
rect 205640 6196 205692 6248
rect 271236 6196 271288 6248
rect 278780 6196 278832 6248
rect 526628 6196 526680 6248
rect 160100 6128 160152 6180
rect 206284 6128 206336 6180
rect 212540 6128 212592 6180
rect 280068 6128 280120 6180
rect 284300 6128 284352 6180
rect 544384 6128 544436 6180
rect 211804 5108 211856 5160
rect 285404 5108 285456 5160
rect 223948 5040 224000 5092
rect 321652 5040 321704 5092
rect 192024 4972 192076 5024
rect 304264 4972 304316 5024
rect 240784 4904 240836 4956
rect 370596 4904 370648 4956
rect 418160 4904 418212 4956
rect 564440 4904 564492 4956
rect 161296 4836 161348 4888
rect 173900 4836 173952 4888
rect 204352 4836 204404 4888
rect 264152 4836 264204 4888
rect 269120 4836 269172 4888
rect 487160 4836 487212 4888
rect 147680 4768 147732 4820
rect 169852 4768 169904 4820
rect 185584 4768 185636 4820
rect 193220 4768 193272 4820
rect 204260 4768 204312 4820
rect 267740 4768 267792 4820
rect 270500 4768 270552 4820
rect 498200 4768 498252 4820
rect 333888 3952 333940 4004
rect 337476 3952 337528 4004
rect 168380 3884 168432 3936
rect 171784 3884 171836 3936
rect 319720 3884 319772 3936
rect 337568 3884 337620 3936
rect 301964 3816 302016 3868
rect 329656 3816 329708 3868
rect 266544 3748 266596 3800
rect 307760 3748 307812 3800
rect 316224 3748 316276 3800
rect 336096 3748 336148 3800
rect 234712 3680 234764 3732
rect 252468 3680 252520 3732
rect 259552 3680 259604 3732
rect 301596 3680 301648 3732
rect 312636 3680 312688 3732
rect 330484 3680 330536 3732
rect 336004 3680 336056 3732
rect 402520 3680 402572 3732
rect 413284 3680 413336 3732
rect 454500 3680 454552 3732
rect 175464 3612 175516 3664
rect 177304 3612 177356 3664
rect 252376 3612 252428 3664
rect 307024 3612 307076 3664
rect 309048 3612 309100 3664
rect 330576 3612 330628 3664
rect 337384 3612 337436 3664
rect 352840 3612 352892 3664
rect 370504 3612 370556 3664
rect 381176 3612 381228 3664
rect 381544 3612 381596 3664
rect 388260 3612 388312 3664
rect 390560 3612 390612 3664
rect 151820 3544 151872 3596
rect 153016 3544 153068 3596
rect 167184 3544 167236 3596
rect 273904 3544 273956 3596
rect 294880 3544 294932 3596
rect 323584 3544 323636 3596
rect 330392 3544 330444 3596
rect 338764 3544 338816 3596
rect 348516 3544 348568 3596
rect 374092 3544 374144 3596
rect 381636 3544 381688 3596
rect 390284 3544 390336 3596
rect 140044 3476 140096 3528
rect 141424 3476 141476 3528
rect 149520 3476 149572 3528
rect 277492 3476 277544 3528
rect 287796 3476 287848 3528
rect 319444 3476 319496 3528
rect 323308 3476 323360 3528
rect 334716 3476 334768 3528
rect 340972 3476 341024 3528
rect 342168 3476 342220 3528
rect 347044 3476 347096 3528
rect 377680 3476 377732 3528
rect 382280 3476 382332 3528
rect 383568 3476 383620 3528
rect 384304 3476 384356 3528
rect 391848 3476 391900 3528
rect 393964 3612 394016 3664
rect 461584 3612 461636 3664
rect 487160 3612 487212 3664
rect 494704 3612 494756 3664
rect 494796 3612 494848 3664
rect 518348 3612 518400 3664
rect 399484 3544 399536 3596
rect 475752 3544 475804 3596
rect 480260 3544 480312 3596
rect 554964 3544 555016 3596
rect 555424 3544 555476 3596
rect 569132 3544 569184 3596
rect 468668 3476 468720 3528
rect 468760 3476 468812 3528
rect 578608 3476 578660 3528
rect 128176 3408 128228 3460
rect 269212 3408 269264 3460
rect 273628 3408 273680 3460
rect 316684 3408 316736 3460
rect 329104 3408 329156 3460
rect 562048 3408 562100 3460
rect 565084 3408 565136 3460
rect 579804 3408 579856 3460
rect 176660 3340 176712 3392
rect 177856 3340 177908 3392
rect 201500 3340 201552 3392
rect 202696 3340 202748 3392
rect 234620 3340 234672 3392
rect 235816 3340 235868 3392
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 355232 3340 355284 3392
rect 356704 3340 356756 3392
rect 358728 3340 358780 3392
rect 359464 3340 359516 3392
rect 365812 3340 365864 3392
rect 367008 3340 367060 3392
rect 377404 3340 377456 3392
rect 384764 3340 384816 3392
rect 390284 3340 390336 3392
rect 394240 3340 394292 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 489920 3340 489972 3392
rect 490748 3340 490800 3392
rect 184296 3272 184348 3324
rect 189724 3272 189776 3324
rect 363604 3136 363656 3188
rect 365812 3136 365864 3188
rect 366364 3068 366416 3120
rect 369400 3068 369452 3120
rect 171968 3000 172020 3052
rect 174544 3000 174596 3052
rect 184204 3000 184256 3052
rect 186136 3000 186188 3052
rect 244924 3000 244976 3052
rect 249984 3000 250036 3052
rect 337476 3000 337528 3052
rect 342904 3000 342956 3052
rect 125876 2932 125928 2984
rect 127624 2932 127676 2984
rect 340972 2932 341024 2984
rect 345664 2932 345716 2984
rect 255872 2864 255924 2916
rect 260104 2864 260156 2916
rect 333980 2796 334032 2848
rect 508872 2796 508924 2848
rect 415400 2728 415452 2780
rect 416688 2728 416740 2780
rect 215300 2388 215352 2440
rect 306748 2388 306800 2440
rect 220820 2320 220872 2372
rect 324412 2320 324464 2372
rect 222200 2252 222252 2304
rect 328000 2252 328052 2304
rect 249800 2184 249852 2236
rect 423772 2184 423824 2236
rect 263600 2116 263652 2168
rect 473452 2116 473504 2168
rect 281540 2048 281592 2100
rect 537208 2048 537260 2100
rect 440240 1912 440292 1964
rect 441528 1912 441580 1964
rect 273260 1300 273312 1352
rect 333980 1300 334032 1352
rect 267924 144 267976 196
rect 487252 144 487304 196
rect 271880 76 271932 128
rect 505560 76 505612 128
rect 280160 8 280212 60
rect 529940 8 529992 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 701010 8156 703520
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 19248 701004 19300 701010
rect 19248 700946 19300 700952
rect 19260 699825 19288 700946
rect 22008 700392 22060 700398
rect 22008 700334 22060 700340
rect 21916 700324 21968 700330
rect 21916 700266 21968 700272
rect 19246 699816 19302 699825
rect 19246 699751 19302 699760
rect 16488 697672 16540 697678
rect 16488 697614 16540 697620
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 606490 2820 658135
rect 2780 606484 2832 606490
rect 2780 606426 2832 606432
rect 2792 606121 2820 606426
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 2792 501809 2820 553823
rect 2870 514856 2926 514865
rect 2870 514791 2872 514800
rect 2924 514791 2926 514800
rect 2872 514762 2924 514768
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 501022 2820 501735
rect 2780 501016 2832 501022
rect 2780 500958 2832 500964
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 398818 2820 449511
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 410106 3188 410479
rect 3148 410100 3200 410106
rect 3148 410042 3200 410048
rect 2780 398812 2832 398818
rect 2780 398754 2832 398760
rect 2792 397497 2820 398754
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 2962 358456 3018 358465
rect 2962 358391 3018 358400
rect 2976 357474 3004 358391
rect 2964 357468 3016 357474
rect 2964 357410 3016 357416
rect 3330 345400 3386 345409
rect 3330 345335 3332 345344
rect 3384 345335 3386 345344
rect 3332 345306 3384 345312
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3344 266422 3372 267135
rect 3332 266416 3384 266422
rect 3332 266358 3384 266364
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3436 204105 3464 566879
rect 3528 332489 3556 671191
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3620 332518 3648 619103
rect 15844 606484 15896 606490
rect 15844 606426 15896 606432
rect 15108 583160 15160 583166
rect 15108 583102 15160 583108
rect 15016 583092 15068 583098
rect 15016 583034 15068 583040
rect 13728 574796 13780 574802
rect 13728 574738 13780 574744
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3608 332512 3660 332518
rect 3514 332480 3570 332489
rect 3608 332454 3660 332460
rect 3514 332415 3570 332424
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3422 204096 3478 204105
rect 3422 204031 3478 204040
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 2792 187746 2820 188799
rect 2780 187740 2832 187746
rect 2780 187682 2832 187688
rect 2962 149832 3018 149841
rect 2962 149767 3018 149776
rect 2976 149122 3004 149767
rect 2964 149116 3016 149122
rect 2964 149058 3016 149064
rect 2778 136776 2834 136785
rect 2778 136711 2780 136720
rect 2832 136711 2834 136720
rect 2780 136682 2832 136688
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3436 110498 3464 110599
rect 3424 110492 3476 110498
rect 3424 110434 3476 110440
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2792 84386 2820 84623
rect 2780 84380 2832 84386
rect 2780 84322 2832 84328
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 30326 3464 71567
rect 3528 61402 3556 293111
rect 4816 203998 4844 514762
rect 7564 501016 7616 501022
rect 7564 500958 7616 500964
rect 6184 410100 6236 410106
rect 6184 410042 6236 410048
rect 4896 240236 4948 240242
rect 4896 240178 4948 240184
rect 4804 203992 4856 203998
rect 4804 203934 4856 203940
rect 4804 187740 4856 187746
rect 4804 187682 4856 187688
rect 3516 61396 3568 61402
rect 3516 61338 3568 61344
rect 4816 46918 4844 187682
rect 4908 48278 4936 240178
rect 4988 136740 5040 136746
rect 4988 136682 5040 136688
rect 5000 51066 5028 136682
rect 5080 84380 5132 84386
rect 5080 84322 5132 84328
rect 4988 51060 5040 51066
rect 4988 51002 5040 51008
rect 4896 48272 4948 48278
rect 4896 48214 4948 48220
rect 4804 46912 4856 46918
rect 4804 46854 4856 46860
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3528 31754 3556 45455
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 3516 31748 3568 31754
rect 3516 31690 3568 31696
rect 3424 30320 3476 30326
rect 3424 30262 3476 30268
rect 3620 26246 3648 32399
rect 5092 28966 5120 84322
rect 6196 75614 6224 410042
rect 6276 357468 6328 357474
rect 6276 357410 6328 357416
rect 6184 75608 6236 75614
rect 6184 75550 6236 75556
rect 6288 41410 6316 357410
rect 6368 149116 6420 149122
rect 6368 149058 6420 149064
rect 6380 49706 6408 149058
rect 6368 49700 6420 49706
rect 6368 49642 6420 49648
rect 6276 41404 6328 41410
rect 6276 41346 6328 41352
rect 7576 39370 7604 500958
rect 13084 462392 13136 462398
rect 13084 462334 13136 462340
rect 7656 398812 7708 398818
rect 7656 398754 7708 398760
rect 7564 39364 7616 39370
rect 7564 39306 7616 39312
rect 7668 33114 7696 398754
rect 8944 345364 8996 345370
rect 8944 345306 8996 345312
rect 8956 42770 8984 345306
rect 10324 318844 10376 318850
rect 10324 318786 10376 318792
rect 9036 110492 9088 110498
rect 9036 110434 9088 110440
rect 8944 42764 8996 42770
rect 8944 42706 8996 42712
rect 9048 36582 9076 110434
rect 10336 44130 10364 318786
rect 12348 214600 12400 214606
rect 12348 214542 12400 214548
rect 12360 69698 12388 214542
rect 13096 76158 13124 462334
rect 13740 459950 13768 574738
rect 15028 460834 15056 583034
rect 15016 460828 15068 460834
rect 15016 460770 15068 460776
rect 14924 460216 14976 460222
rect 14924 460158 14976 460164
rect 14936 459950 14964 460158
rect 13728 459944 13780 459950
rect 13728 459886 13780 459892
rect 14924 459944 14976 459950
rect 14924 459886 14976 459892
rect 13176 442264 13228 442270
rect 13176 442206 13228 442212
rect 13188 214606 13216 442206
rect 14936 332722 14964 459886
rect 14924 332716 14976 332722
rect 14924 332658 14976 332664
rect 15028 332654 15056 460770
rect 15120 455394 15148 583102
rect 15108 455388 15160 455394
rect 15108 455330 15160 455336
rect 15108 332716 15160 332722
rect 15108 332658 15160 332664
rect 15016 332648 15068 332654
rect 15016 332590 15068 332596
rect 13176 214600 13228 214606
rect 13176 214542 13228 214548
rect 13268 213988 13320 213994
rect 13268 213930 13320 213936
rect 13084 76152 13136 76158
rect 13084 76094 13136 76100
rect 12348 69692 12400 69698
rect 12348 69634 12400 69640
rect 13084 61396 13136 61402
rect 13084 61338 13136 61344
rect 13096 45558 13124 61338
rect 13280 53106 13308 213930
rect 14832 204604 14884 204610
rect 14832 204546 14884 204552
rect 14844 73166 14872 204546
rect 15028 200054 15056 332590
rect 15016 200048 15068 200054
rect 15016 199990 15068 199996
rect 14924 199504 14976 199510
rect 14924 199446 14976 199452
rect 14832 73160 14884 73166
rect 14832 73102 14884 73108
rect 14936 73030 14964 199446
rect 14924 73024 14976 73030
rect 14924 72966 14976 72972
rect 15028 71738 15056 199990
rect 15120 199986 15148 332658
rect 15108 199980 15160 199986
rect 15108 199922 15160 199928
rect 15016 71732 15068 71738
rect 15016 71674 15068 71680
rect 13268 53100 13320 53106
rect 13268 53042 13320 53048
rect 13084 45552 13136 45558
rect 13084 45494 13136 45500
rect 10324 44124 10376 44130
rect 10324 44066 10376 44072
rect 9036 36576 9088 36582
rect 9036 36518 9088 36524
rect 15856 34474 15884 606426
rect 16396 572348 16448 572354
rect 16396 572290 16448 572296
rect 16408 461038 16436 572290
rect 16396 461032 16448 461038
rect 16396 460974 16448 460980
rect 16394 460184 16450 460193
rect 16394 460119 16450 460128
rect 16408 335354 16436 460119
rect 16316 335326 16436 335354
rect 16316 331158 16344 335326
rect 16304 331152 16356 331158
rect 16304 331094 16356 331100
rect 16316 204542 16344 331094
rect 16396 315988 16448 315994
rect 16396 315930 16448 315936
rect 16304 204536 16356 204542
rect 16304 204478 16356 204484
rect 16408 188970 16436 315930
rect 16396 188964 16448 188970
rect 16396 188906 16448 188912
rect 16408 77994 16436 188906
rect 16396 77988 16448 77994
rect 16396 77930 16448 77936
rect 16500 35902 16528 697614
rect 21928 586498 21956 700266
rect 21916 586492 21968 586498
rect 21916 586434 21968 586440
rect 21824 586152 21876 586158
rect 21824 586094 21876 586100
rect 21732 586016 21784 586022
rect 21732 585958 21784 585964
rect 17868 583296 17920 583302
rect 17868 583238 17920 583244
rect 17776 583228 17828 583234
rect 17776 583170 17828 583176
rect 17684 574864 17736 574870
rect 17684 574806 17736 574812
rect 17592 461032 17644 461038
rect 17592 460974 17644 460980
rect 17224 454708 17276 454714
rect 17224 454650 17276 454656
rect 17236 315994 17264 454650
rect 17408 334008 17460 334014
rect 17408 333950 17460 333956
rect 17224 315988 17276 315994
rect 17224 315930 17276 315936
rect 17132 199980 17184 199986
rect 17132 199922 17184 199928
rect 17144 199209 17172 199922
rect 17130 199200 17186 199209
rect 17130 199135 17186 199144
rect 17420 186017 17448 333950
rect 17604 329798 17632 460974
rect 17696 460766 17724 574806
rect 17788 460902 17816 583170
rect 17776 460896 17828 460902
rect 17776 460838 17828 460844
rect 17684 460760 17736 460766
rect 17684 460702 17736 460708
rect 17696 331090 17724 460702
rect 17880 458862 17908 583238
rect 19156 583024 19208 583030
rect 19156 582966 19208 582972
rect 19064 572280 19116 572286
rect 19064 572222 19116 572228
rect 19076 459406 19104 572222
rect 19064 459400 19116 459406
rect 19064 459342 19116 459348
rect 17868 458856 17920 458862
rect 18788 458856 18840 458862
rect 17868 458798 17920 458804
rect 18786 458824 18788 458833
rect 18840 458824 18842 458833
rect 18786 458759 18842 458768
rect 17868 455388 17920 455394
rect 17868 455330 17920 455336
rect 17880 454714 17908 455330
rect 17868 454708 17920 454714
rect 17868 454650 17920 454656
rect 17684 331084 17736 331090
rect 17684 331026 17736 331032
rect 17592 329792 17644 329798
rect 17592 329734 17644 329740
rect 17500 204740 17552 204746
rect 17500 204682 17552 204688
rect 17406 186008 17462 186017
rect 17406 185943 17462 185952
rect 17512 72894 17540 204682
rect 17696 204474 17724 331026
rect 17776 329792 17828 329798
rect 17776 329734 17828 329740
rect 17684 204468 17736 204474
rect 17684 204410 17736 204416
rect 17592 198756 17644 198762
rect 17592 198698 17644 198704
rect 17604 74497 17632 198698
rect 17696 76090 17724 204410
rect 17788 199918 17816 329734
rect 18800 315246 18828 458759
rect 18880 332988 18932 332994
rect 18880 332930 18932 332936
rect 18788 315240 18840 315246
rect 18788 315182 18840 315188
rect 18788 204536 18840 204542
rect 18788 204478 18840 204484
rect 17776 199912 17828 199918
rect 17776 199854 17828 199860
rect 17788 198762 17816 199854
rect 17776 198756 17828 198762
rect 17776 198698 17828 198704
rect 17868 185972 17920 185978
rect 17868 185914 17920 185920
rect 17684 76084 17736 76090
rect 17684 76026 17736 76032
rect 17590 74488 17646 74497
rect 17590 74423 17646 74432
rect 17880 73098 17908 185914
rect 18800 75954 18828 204478
rect 18892 204202 18920 332930
rect 18972 330676 19024 330682
rect 18972 330618 19024 330624
rect 18984 204746 19012 330618
rect 19076 329730 19104 459342
rect 19168 455394 19196 582966
rect 20536 572212 20588 572218
rect 20536 572154 20588 572160
rect 19248 572076 19300 572082
rect 19248 572018 19300 572024
rect 19260 458862 19288 572018
rect 20444 572008 20496 572014
rect 20350 571976 20406 571985
rect 20444 571950 20496 571956
rect 20350 571911 20406 571920
rect 20364 460970 20392 571911
rect 20352 460964 20404 460970
rect 20272 460912 20352 460934
rect 20272 460906 20404 460912
rect 19248 458856 19300 458862
rect 19248 458798 19300 458804
rect 19156 455388 19208 455394
rect 19156 455330 19208 455336
rect 19168 330954 19196 455330
rect 20272 332858 20300 460906
rect 20456 459338 20484 571950
rect 20444 459332 20496 459338
rect 20444 459274 20496 459280
rect 20352 458856 20404 458862
rect 20352 458798 20404 458804
rect 20364 332926 20392 458798
rect 20456 333266 20484 459274
rect 20548 458998 20576 572154
rect 20628 572144 20680 572150
rect 20628 572086 20680 572092
rect 20640 459474 20668 572086
rect 20628 459468 20680 459474
rect 20628 459410 20680 459416
rect 20536 458992 20588 458998
rect 20536 458934 20588 458940
rect 20444 333260 20496 333266
rect 20444 333202 20496 333208
rect 20456 332994 20484 333202
rect 20444 332988 20496 332994
rect 20444 332930 20496 332936
rect 20352 332920 20404 332926
rect 20352 332862 20404 332868
rect 20260 332852 20312 332858
rect 20260 332794 20312 332800
rect 20168 332784 20220 332790
rect 20168 332726 20220 332732
rect 19156 330948 19208 330954
rect 19156 330890 19208 330896
rect 19168 330682 19196 330890
rect 19156 330676 19208 330682
rect 19156 330618 19208 330624
rect 19064 329724 19116 329730
rect 19064 329666 19116 329672
rect 18972 204740 19024 204746
rect 18972 204682 19024 204688
rect 18984 204406 19012 204682
rect 18972 204400 19024 204406
rect 18972 204342 19024 204348
rect 18880 204196 18932 204202
rect 18880 204138 18932 204144
rect 18892 200114 18920 204138
rect 19076 203930 19104 329666
rect 19340 315240 19392 315246
rect 19340 315182 19392 315188
rect 19352 204762 19380 315182
rect 20180 229094 20208 332726
rect 20272 325694 20300 332794
rect 20364 332790 20392 332862
rect 20352 332784 20404 332790
rect 20352 332726 20404 332732
rect 20272 325666 20576 325694
rect 20180 229066 20392 229094
rect 19260 204734 19380 204762
rect 19260 203946 19288 204734
rect 20364 204241 20392 229066
rect 20444 204264 20496 204270
rect 20350 204232 20406 204241
rect 20444 204206 20496 204212
rect 20350 204167 20406 204176
rect 20364 204134 20392 204167
rect 20352 204128 20404 204134
rect 20352 204070 20404 204076
rect 20456 204066 20484 204206
rect 20444 204060 20496 204066
rect 20444 204002 20496 204008
rect 19338 203960 19394 203969
rect 19064 203924 19116 203930
rect 19064 203866 19116 203872
rect 19260 203918 19338 203946
rect 18892 200086 19196 200114
rect 18972 187740 19024 187746
rect 18972 187682 19024 187688
rect 18984 76022 19012 187682
rect 18972 76016 19024 76022
rect 18972 75958 19024 75964
rect 18788 75948 18840 75954
rect 18788 75890 18840 75896
rect 19168 75886 19196 200086
rect 19156 75880 19208 75886
rect 19156 75822 19208 75828
rect 19260 74526 19288 203918
rect 19338 203895 19394 203904
rect 20352 203924 20404 203930
rect 20352 203866 20404 203872
rect 20364 203590 20392 203866
rect 20352 203584 20404 203590
rect 20352 203526 20404 203532
rect 20364 75750 20392 203526
rect 20456 75818 20484 204002
rect 20548 199102 20576 325666
rect 20640 315858 20668 459410
rect 21640 458992 21692 458998
rect 21640 458934 21692 458940
rect 21364 444372 21416 444378
rect 21364 444314 21416 444320
rect 21376 334014 21404 444314
rect 21364 334008 21416 334014
rect 21364 333950 21416 333956
rect 21376 332790 21404 333950
rect 21364 332784 21416 332790
rect 21364 332726 21416 332732
rect 21652 331809 21680 458934
rect 21744 457910 21772 585958
rect 21732 457904 21784 457910
rect 21732 457846 21784 457852
rect 21744 457042 21772 457846
rect 21836 457502 21864 586094
rect 21916 585880 21968 585886
rect 21916 585822 21968 585828
rect 21928 458114 21956 585822
rect 22020 459542 22048 700334
rect 24320 699718 24348 703520
rect 72988 701010 73016 703520
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 89180 700398 89208 703520
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 137848 700210 137876 703520
rect 138020 700392 138072 700398
rect 138020 700334 138072 700340
rect 138032 700210 138060 700334
rect 137848 700182 138060 700210
rect 22100 699712 22152 699718
rect 22100 699654 22152 699660
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 22112 461106 22140 699654
rect 138032 697678 138060 700182
rect 138020 697672 138072 697678
rect 138020 697614 138072 697620
rect 154132 697610 154160 703520
rect 202800 700398 202828 703520
rect 202788 700392 202840 700398
rect 202788 700334 202840 700340
rect 218992 700330 219020 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 397472 700369 397500 700946
rect 397458 700360 397514 700369
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 302148 700324 302200 700330
rect 397458 700295 397514 700304
rect 302148 700266 302200 700272
rect 22192 697604 22244 697610
rect 22192 697546 22244 697552
rect 154120 697604 154172 697610
rect 154120 697546 154172 697552
rect 22204 596174 22232 697546
rect 22204 596146 23060 596174
rect 23032 588690 23060 596146
rect 23032 588662 23460 588690
rect 28184 587302 28520 587330
rect 33244 587302 33580 587330
rect 38304 587302 38640 587330
rect 43364 587302 43700 587330
rect 48516 587302 48760 587330
rect 53484 587302 53820 587330
rect 57992 587302 58880 587330
rect 63604 587302 63940 587330
rect 67652 587302 69000 587330
rect 73172 587302 74060 587330
rect 78692 587302 79120 587330
rect 83844 587302 84180 587330
rect 88352 587302 89240 587330
rect 93964 587302 94300 587330
rect 99024 587302 99360 587330
rect 104084 587302 104420 587330
rect 109052 587302 109480 587330
rect 114204 587302 114540 587330
rect 119264 587302 119600 587330
rect 124324 587302 124660 587330
rect 128372 587302 129720 587330
rect 134444 587302 134780 587330
rect 139504 587302 139840 587330
rect 144840 587302 144900 587330
rect 28184 586498 28212 587302
rect 28172 586492 28224 586498
rect 28172 586434 28224 586440
rect 23296 586084 23348 586090
rect 23296 586026 23348 586032
rect 23202 585848 23258 585857
rect 23112 585812 23164 585818
rect 23202 585783 23258 585792
rect 23112 585754 23164 585760
rect 22100 461100 22152 461106
rect 22100 461042 22152 461048
rect 23124 460934 23152 585754
rect 22940 460906 23152 460934
rect 22008 459536 22060 459542
rect 22008 459478 22060 459484
rect 22940 458969 22968 460906
rect 22926 458960 22982 458969
rect 22926 458895 22982 458904
rect 21916 458108 21968 458114
rect 21916 458050 21968 458056
rect 21824 457496 21876 457502
rect 21824 457438 21876 457444
rect 21744 457014 21864 457042
rect 21732 456884 21784 456890
rect 21732 456826 21784 456832
rect 21744 332246 21772 456826
rect 21836 451274 21864 457014
rect 22744 456816 22796 456822
rect 22744 456758 22796 456764
rect 21836 451246 22048 451274
rect 21732 332240 21784 332246
rect 21732 332182 21784 332188
rect 21638 331800 21694 331809
rect 21638 331735 21694 331744
rect 20628 315852 20680 315858
rect 20628 315794 20680 315800
rect 20640 204270 20668 315794
rect 20904 266416 20956 266422
rect 20904 266358 20956 266364
rect 20916 258074 20944 266358
rect 20916 258046 21404 258074
rect 20628 204264 20680 204270
rect 20628 204206 20680 204212
rect 20626 202872 20682 202881
rect 20626 202807 20682 202816
rect 20536 199096 20588 199102
rect 20536 199038 20588 199044
rect 20536 198008 20588 198014
rect 20536 197950 20588 197956
rect 20548 77110 20576 197950
rect 20536 77104 20588 77110
rect 20536 77046 20588 77052
rect 20444 75812 20496 75818
rect 20444 75754 20496 75760
rect 20352 75744 20404 75750
rect 20352 75686 20404 75692
rect 19248 74520 19300 74526
rect 19248 74462 19300 74468
rect 20640 74458 20668 202807
rect 20628 74452 20680 74458
rect 20628 74394 20680 74400
rect 17868 73092 17920 73098
rect 17868 73034 17920 73040
rect 17500 72888 17552 72894
rect 17500 72830 17552 72836
rect 21376 48210 21404 258046
rect 21744 202638 21772 332182
rect 21824 332036 21876 332042
rect 21824 331978 21876 331984
rect 21836 202706 21864 331978
rect 22020 331922 22048 451246
rect 22756 332586 22784 456758
rect 22940 345014 22968 458895
rect 23112 458108 23164 458114
rect 23112 458050 23164 458056
rect 23020 457496 23072 457502
rect 23020 457438 23072 457444
rect 22848 344986 22968 345014
rect 22744 332580 22796 332586
rect 22744 332522 22796 332528
rect 22756 332042 22784 332522
rect 22848 332382 22876 344986
rect 23032 335354 23060 457438
rect 22940 335326 23060 335354
rect 22940 332450 22968 335326
rect 23124 333418 23152 458050
rect 23216 457978 23244 585783
rect 23308 458182 23336 586026
rect 29644 585948 29696 585954
rect 29644 585890 29696 585896
rect 29656 572354 29684 585890
rect 33244 585886 33272 587302
rect 33232 585880 33284 585886
rect 33232 585822 33284 585828
rect 35164 585880 35216 585886
rect 35164 585822 35216 585828
rect 35176 574870 35204 585822
rect 38304 585818 38332 587302
rect 43364 586158 43392 587302
rect 43352 586152 43404 586158
rect 43352 586094 43404 586100
rect 48516 586090 48544 587302
rect 48504 586084 48556 586090
rect 48504 586026 48556 586032
rect 53484 586022 53512 587302
rect 53472 586016 53524 586022
rect 53472 585958 53524 585964
rect 38292 585812 38344 585818
rect 38292 585754 38344 585760
rect 39304 585812 39356 585818
rect 39304 585754 39356 585760
rect 35164 574864 35216 574870
rect 35164 574806 35216 574812
rect 29644 572348 29696 572354
rect 29644 572290 29696 572296
rect 39316 570625 39344 585754
rect 57992 572286 58020 587302
rect 63604 585857 63632 587302
rect 63590 585848 63646 585857
rect 63590 585783 63646 585792
rect 57980 572280 58032 572286
rect 57980 572222 58032 572228
rect 67652 572218 67680 587302
rect 67640 572212 67692 572218
rect 67640 572154 67692 572160
rect 73172 572150 73200 587302
rect 73160 572144 73212 572150
rect 73160 572086 73212 572092
rect 78692 572082 78720 587302
rect 83844 585721 83872 587302
rect 83830 585712 83886 585721
rect 83830 585647 83886 585656
rect 78680 572076 78732 572082
rect 78680 572018 78732 572024
rect 88352 572014 88380 587302
rect 93964 583302 93992 587302
rect 93952 583296 94004 583302
rect 93952 583238 94004 583244
rect 99024 583234 99052 587302
rect 104084 585954 104112 587302
rect 104072 585948 104124 585954
rect 104072 585890 104124 585896
rect 99012 583228 99064 583234
rect 99012 583170 99064 583176
rect 88340 572008 88392 572014
rect 109052 571985 109080 587302
rect 114204 583166 114232 587302
rect 119264 585886 119292 587302
rect 119252 585880 119304 585886
rect 119252 585822 119304 585828
rect 124324 585818 124352 587302
rect 124312 585812 124364 585818
rect 124312 585754 124364 585760
rect 114192 583160 114244 583166
rect 114192 583102 114244 583108
rect 128372 574802 128400 587302
rect 134444 583001 134472 587302
rect 139504 583098 139532 587302
rect 144840 586498 144868 587302
rect 149946 587058 149974 587316
rect 154776 587302 155020 587330
rect 158732 587302 160080 587330
rect 165140 587302 165476 587330
rect 149946 587030 150020 587058
rect 149992 586498 150020 587030
rect 144828 586492 144880 586498
rect 144828 586434 144880 586440
rect 149980 586492 150032 586498
rect 149980 586434 150032 586440
rect 149992 585857 150020 586434
rect 149978 585848 150034 585857
rect 149978 585783 150034 585792
rect 139492 583092 139544 583098
rect 139492 583034 139544 583040
rect 154776 583030 154804 587302
rect 154764 583024 154816 583030
rect 134430 582992 134486 583001
rect 154764 582966 154816 582972
rect 134430 582927 134486 582936
rect 128360 574796 128412 574802
rect 128360 574738 128412 574744
rect 158732 572014 158760 587302
rect 165448 580310 165476 587302
rect 169772 587302 170200 587330
rect 175200 587302 175260 587330
rect 180320 587302 180656 587330
rect 185380 587302 185716 587330
rect 165436 580304 165488 580310
rect 165436 580246 165488 580252
rect 169772 577522 169800 587302
rect 175200 580281 175228 587302
rect 180628 580378 180656 587302
rect 185688 580514 185716 587302
rect 190380 587302 190440 587330
rect 195500 587302 195836 587330
rect 200560 587302 200896 587330
rect 185676 580508 185728 580514
rect 185676 580450 185728 580456
rect 190380 580446 190408 587302
rect 195808 580582 195836 587302
rect 200868 583030 200896 587302
rect 204272 587302 205620 587330
rect 210680 587302 211016 587330
rect 215740 587302 216076 587330
rect 200856 583024 200908 583030
rect 200856 582966 200908 582972
rect 195796 580576 195848 580582
rect 195796 580518 195848 580524
rect 190368 580440 190420 580446
rect 190368 580382 190420 580388
rect 180616 580372 180668 580378
rect 180616 580314 180668 580320
rect 175186 580272 175242 580281
rect 175186 580207 175242 580216
rect 169760 577516 169812 577522
rect 169760 577458 169812 577464
rect 158720 572008 158772 572014
rect 88340 571950 88392 571956
rect 109038 571976 109094 571985
rect 204272 571985 204300 587302
rect 210988 583001 211016 587302
rect 216048 583098 216076 587302
rect 220740 587302 220800 587330
rect 225860 587302 226196 587330
rect 230920 587302 231256 587330
rect 220740 583166 220768 587302
rect 226168 585721 226196 587302
rect 226154 585712 226210 585721
rect 226154 585647 226210 585656
rect 231228 583234 231256 587302
rect 235920 587302 235980 587330
rect 241040 587302 241376 587330
rect 235920 583302 235948 587302
rect 241348 585818 241376 587302
rect 245672 587302 246100 587330
rect 251100 587302 251160 587330
rect 256220 587302 256556 587330
rect 261280 587302 261616 587330
rect 241336 585812 241388 585818
rect 241336 585754 241388 585760
rect 235908 583296 235960 583302
rect 235908 583238 235960 583244
rect 231216 583228 231268 583234
rect 231216 583170 231268 583176
rect 220728 583160 220780 583166
rect 220728 583102 220780 583108
rect 216036 583092 216088 583098
rect 216036 583034 216088 583040
rect 210974 582992 211030 583001
rect 210974 582927 211030 582936
rect 245672 572082 245700 587302
rect 251100 585886 251128 587302
rect 256528 585954 256556 587302
rect 261588 586022 261616 587302
rect 266280 587302 266340 587330
rect 270512 587302 271400 587330
rect 276032 587302 276460 587330
rect 281460 587302 281520 587330
rect 286428 587302 286580 587330
rect 266280 586090 266308 587302
rect 266268 586084 266320 586090
rect 266268 586026 266320 586032
rect 261576 586016 261628 586022
rect 261576 585958 261628 585964
rect 256516 585948 256568 585954
rect 256516 585890 256568 585896
rect 251088 585880 251140 585886
rect 251088 585822 251140 585828
rect 270512 572150 270540 587302
rect 270500 572144 270552 572150
rect 276032 572121 276060 587302
rect 281460 585206 281488 587302
rect 281448 585200 281500 585206
rect 286428 585177 286456 587302
rect 302160 586498 302188 700266
rect 413664 698970 413692 703520
rect 462332 701010 462360 703520
rect 462320 701004 462372 701010
rect 462320 700946 462372 700952
rect 478524 700330 478552 703520
rect 527192 702434 527220 703520
rect 527192 702406 527312 702434
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 302240 698964 302292 698970
rect 302240 698906 302292 698912
rect 413652 698964 413704 698970
rect 413652 698906 413704 698912
rect 302252 596174 302280 698906
rect 527192 697513 527220 700266
rect 527284 699825 527312 702406
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 527270 699816 527326 699825
rect 527270 699751 527326 699760
rect 527284 698290 527312 699751
rect 527272 698284 527324 698290
rect 527272 698226 527324 698232
rect 580172 698284 580224 698290
rect 580172 698226 580224 698232
rect 527178 697504 527234 697513
rect 527178 697439 527234 697448
rect 580184 697241 580212 698226
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 302252 596146 303016 596174
rect 302988 588690 303016 596146
rect 302988 588662 303462 588690
rect 308508 586498 308536 587316
rect 302148 586492 302200 586498
rect 302148 586434 302200 586440
rect 308496 586492 308548 586498
rect 308496 586434 308548 586440
rect 313568 586090 313596 587316
rect 290004 586084 290056 586090
rect 290004 586026 290056 586032
rect 302056 586084 302108 586090
rect 302056 586026 302108 586032
rect 313556 586084 313608 586090
rect 313556 586026 313608 586032
rect 289912 586016 289964 586022
rect 289912 585958 289964 585964
rect 288532 585948 288584 585954
rect 288532 585890 288584 585896
rect 287612 585812 287664 585818
rect 287612 585754 287664 585760
rect 287518 585712 287574 585721
rect 287518 585647 287574 585656
rect 281448 585142 281500 585148
rect 286414 585168 286470 585177
rect 286414 585103 286470 585112
rect 270500 572086 270552 572092
rect 276018 572112 276074 572121
rect 245660 572076 245712 572082
rect 276018 572047 276074 572056
rect 245660 572018 245712 572024
rect 158720 571950 158772 571956
rect 204258 571976 204314 571985
rect 109038 571911 109094 571920
rect 204258 571911 204314 571920
rect 39302 570616 39358 570625
rect 39302 570551 39358 570560
rect 286230 461952 286286 461961
rect 286230 461887 286286 461896
rect 285588 461644 285640 461650
rect 285588 461586 285640 461592
rect 23400 461230 23460 461258
rect 28184 461230 28520 461258
rect 33244 461230 33580 461258
rect 38304 461230 38640 461258
rect 43364 461230 43700 461258
rect 48516 461230 48760 461258
rect 53484 461230 53820 461258
rect 58544 461230 58880 461258
rect 63604 461230 63940 461258
rect 68664 461230 69000 461258
rect 73724 461230 74060 461258
rect 78784 461230 79120 461258
rect 83844 461230 84180 461258
rect 88904 461230 89240 461258
rect 93964 461230 94300 461258
rect 99024 461230 99360 461258
rect 23400 461106 23428 461230
rect 24952 461168 25004 461174
rect 24952 461110 25004 461116
rect 23388 461100 23440 461106
rect 23388 461042 23440 461048
rect 24860 460964 24912 460970
rect 24860 460906 24912 460912
rect 24872 460834 24900 460906
rect 24964 460902 24992 461110
rect 24952 460896 25004 460902
rect 24952 460838 25004 460844
rect 24860 460828 24912 460834
rect 24860 460770 24912 460776
rect 24858 460320 24914 460329
rect 24858 460255 24914 460264
rect 23296 458176 23348 458182
rect 23296 458118 23348 458124
rect 23204 457972 23256 457978
rect 23204 457914 23256 457920
rect 23216 456890 23244 457914
rect 23204 456884 23256 456890
rect 23204 456826 23256 456832
rect 23308 456822 23336 458118
rect 23296 456816 23348 456822
rect 23296 456758 23348 456764
rect 24872 444378 24900 460255
rect 24860 444372 24912 444378
rect 24860 444314 24912 444320
rect 24964 444281 24992 460838
rect 28184 459542 28212 461230
rect 28172 459536 28224 459542
rect 28172 459478 28224 459484
rect 33244 458522 33272 461230
rect 38304 458998 38332 461230
rect 34520 458992 34572 458998
rect 34518 458960 34520 458969
rect 38292 458992 38344 458998
rect 34572 458960 34574 458969
rect 38292 458934 38344 458940
rect 34518 458895 34574 458904
rect 27804 458516 27856 458522
rect 27804 458458 27856 458464
rect 33232 458516 33284 458522
rect 33232 458458 33284 458464
rect 27816 458114 27844 458458
rect 30932 458176 30984 458182
rect 30932 458118 30984 458124
rect 27804 458108 27856 458114
rect 27804 458050 27856 458056
rect 30944 457842 30972 458118
rect 30932 457836 30984 457842
rect 30932 457778 30984 457784
rect 43364 457502 43392 461230
rect 48516 458046 48544 461230
rect 53484 458114 53512 461230
rect 58544 459406 58572 461230
rect 58532 459400 58584 459406
rect 58532 459342 58584 459348
rect 63604 458182 63632 461230
rect 68664 458930 68692 461230
rect 73724 459474 73752 461230
rect 73712 459468 73764 459474
rect 73712 459410 73764 459416
rect 68652 458924 68704 458930
rect 68652 458866 68704 458872
rect 78784 458862 78812 461230
rect 78772 458856 78824 458862
rect 78772 458798 78824 458804
rect 63592 458176 63644 458182
rect 83844 458153 83872 461230
rect 88904 459338 88932 461230
rect 88892 459332 88944 459338
rect 88892 459274 88944 459280
rect 93964 458833 93992 461230
rect 99024 461174 99052 461230
rect 99012 461168 99064 461174
rect 99012 461110 99064 461116
rect 104406 461106 104434 461244
rect 104394 461100 104446 461106
rect 104394 461042 104446 461048
rect 109466 461038 109494 461244
rect 114204 461230 114540 461258
rect 119264 461230 119600 461258
rect 124324 461230 124660 461258
rect 129384 461230 129720 461258
rect 134444 461230 134780 461258
rect 139504 461230 139840 461258
rect 144840 461230 144900 461258
rect 109454 461032 109506 461038
rect 109454 460974 109506 460980
rect 93950 458824 94006 458833
rect 93950 458759 94006 458768
rect 114204 458250 114232 461230
rect 119264 460902 119292 461230
rect 119252 460896 119304 460902
rect 119252 460838 119304 460844
rect 124324 460329 124352 461230
rect 124310 460320 124366 460329
rect 124310 460255 124366 460264
rect 129384 460222 129412 461230
rect 129372 460216 129424 460222
rect 134444 460193 134472 461230
rect 139504 460970 139532 461230
rect 139492 460964 139544 460970
rect 139492 460906 139544 460912
rect 129372 460158 129424 460164
rect 134430 460184 134486 460193
rect 134430 460119 134486 460128
rect 144840 459542 144868 461230
rect 149946 461122 149974 461244
rect 154776 461230 155020 461258
rect 160020 461230 160080 461258
rect 164252 461230 165140 461258
rect 169772 461230 170200 461258
rect 175200 461230 175260 461258
rect 180320 461230 180656 461258
rect 185380 461230 185716 461258
rect 149946 461094 150020 461122
rect 149992 459542 150020 461094
rect 144828 459536 144880 459542
rect 144828 459478 144880 459484
rect 149980 459536 150032 459542
rect 149980 459478 150032 459484
rect 149992 458862 150020 459478
rect 149980 458856 150032 458862
rect 149980 458798 150032 458804
rect 110420 458244 110472 458250
rect 110420 458186 110472 458192
rect 114192 458244 114244 458250
rect 114192 458186 114244 458192
rect 63592 458118 63644 458124
rect 83830 458144 83886 458153
rect 53472 458108 53524 458114
rect 83830 458079 83886 458088
rect 53472 458050 53524 458056
rect 48504 458040 48556 458046
rect 48504 457982 48556 457988
rect 43352 457496 43404 457502
rect 43352 457438 43404 457444
rect 110432 454714 110460 458186
rect 154776 455394 154804 461230
rect 160020 460873 160048 461230
rect 160006 460864 160062 460873
rect 160006 460799 160062 460808
rect 154764 455388 154816 455394
rect 154764 455330 154816 455336
rect 110420 454708 110472 454714
rect 110420 454650 110472 454656
rect 24950 444272 25006 444281
rect 24950 444207 25006 444216
rect 23480 443692 23532 443698
rect 23480 443634 23532 443640
rect 23492 442270 23520 443634
rect 164252 442950 164280 461230
rect 164240 442944 164292 442950
rect 164240 442886 164292 442892
rect 169772 442882 169800 461230
rect 175200 460193 175228 461230
rect 175186 460184 175242 460193
rect 175186 460119 175242 460128
rect 180628 458930 180656 461230
rect 185688 459474 185716 461230
rect 190426 460934 190454 461244
rect 195500 461230 195836 461258
rect 190426 460906 190500 460934
rect 190472 460222 190500 460906
rect 190460 460216 190512 460222
rect 190460 460158 190512 460164
rect 195808 459542 195836 461230
rect 200132 461230 200560 461258
rect 204272 461230 205620 461258
rect 210680 461230 211108 461258
rect 215740 461230 216076 461258
rect 195796 459536 195848 459542
rect 195796 459478 195848 459484
rect 185676 459468 185728 459474
rect 185676 459410 185728 459416
rect 180616 458924 180668 458930
rect 180616 458866 180668 458872
rect 200132 443698 200160 461230
rect 204272 443737 204300 461230
rect 211080 459490 211108 461230
rect 211080 459462 211200 459490
rect 211172 458153 211200 459462
rect 216048 458998 216076 461230
rect 219452 461230 220800 461258
rect 225860 461230 226196 461258
rect 230920 461230 231256 461258
rect 216036 458992 216088 458998
rect 216036 458934 216088 458940
rect 211158 458144 211214 458153
rect 211158 458079 211214 458088
rect 219452 444378 219480 461230
rect 226168 458182 226196 461230
rect 226156 458176 226208 458182
rect 226156 458118 226208 458124
rect 231228 458114 231256 461230
rect 235920 461230 235980 461258
rect 241040 461230 241376 461258
rect 246100 461230 246436 461258
rect 231216 458108 231268 458114
rect 231216 458050 231268 458056
rect 235920 457502 235948 461230
rect 241348 460902 241376 461230
rect 241336 460896 241388 460902
rect 241336 460838 241388 460844
rect 246408 460834 246436 461230
rect 251100 461230 251160 461258
rect 256220 461230 256556 461258
rect 261280 461230 261616 461258
rect 246396 460828 246448 460834
rect 246396 460770 246448 460776
rect 251100 458046 251128 461230
rect 256528 460766 256556 461230
rect 256516 460760 256568 460766
rect 256516 460702 256568 460708
rect 251088 458040 251140 458046
rect 251088 457982 251140 457988
rect 261588 457570 261616 461230
rect 266280 461230 266340 461258
rect 270512 461230 271400 461258
rect 276460 461230 276796 461258
rect 266280 459406 266308 461230
rect 266268 459400 266320 459406
rect 266268 459342 266320 459348
rect 261576 457564 261628 457570
rect 261576 457506 261628 457512
rect 235908 457496 235960 457502
rect 235908 457438 235960 457444
rect 219440 444372 219492 444378
rect 219440 444314 219492 444320
rect 270512 444310 270540 461230
rect 276768 459105 276796 461230
rect 281460 461230 281520 461258
rect 281460 459513 281488 461230
rect 285496 460284 285548 460290
rect 285496 460226 285548 460232
rect 285310 460184 285366 460193
rect 285310 460119 285366 460128
rect 281446 459504 281502 459513
rect 281446 459439 281502 459448
rect 276754 459096 276810 459105
rect 276754 459031 276810 459040
rect 285324 451274 285352 460119
rect 285404 459468 285456 459474
rect 285404 459410 285456 459416
rect 285416 458289 285444 459410
rect 285402 458280 285458 458289
rect 285402 458215 285458 458224
rect 285324 451246 285444 451274
rect 270500 444304 270552 444310
rect 270500 444246 270552 444252
rect 285416 443873 285444 451246
rect 285402 443864 285458 443873
rect 285402 443799 285458 443808
rect 204258 443728 204314 443737
rect 200120 443692 200172 443698
rect 204258 443663 204314 443672
rect 200120 443634 200172 443640
rect 284300 442944 284352 442950
rect 284300 442886 284352 442892
rect 169760 442876 169812 442882
rect 169760 442818 169812 442824
rect 284312 442270 284340 442886
rect 284944 442876 284996 442882
rect 284944 442818 284996 442824
rect 23480 442264 23532 442270
rect 23480 442206 23532 442212
rect 284300 442264 284352 442270
rect 284300 442206 284352 442212
rect 284956 441930 284984 442818
rect 285508 442270 285536 460226
rect 285600 442882 285628 461586
rect 286244 456929 286272 461887
rect 286580 461230 286916 461258
rect 286324 460760 286376 460766
rect 286322 460728 286324 460737
rect 286376 460728 286378 460737
rect 286322 460663 286378 460672
rect 286888 458969 286916 461230
rect 286874 458960 286930 458969
rect 286874 458895 286930 458904
rect 287532 458182 287560 585647
rect 287624 460902 287652 585754
rect 287796 580508 287848 580514
rect 287796 580450 287848 580456
rect 287612 460896 287664 460902
rect 287612 460838 287664 460844
rect 287624 459649 287652 460838
rect 287704 460080 287756 460086
rect 287704 460022 287756 460028
rect 287610 459640 287666 459649
rect 287610 459575 287666 459584
rect 287716 459513 287744 460022
rect 287702 459504 287758 459513
rect 287808 459474 287836 580450
rect 288544 460766 288572 585890
rect 289820 585880 289872 585886
rect 289820 585822 289872 585828
rect 288624 585200 288676 585206
rect 288624 585142 288676 585148
rect 288532 460760 288584 460766
rect 288532 460702 288584 460708
rect 288636 460086 288664 585142
rect 288808 583228 288860 583234
rect 288808 583170 288860 583176
rect 288716 572008 288768 572014
rect 288716 571950 288768 571956
rect 288728 460329 288756 571950
rect 288714 460320 288770 460329
rect 288714 460255 288770 460264
rect 288624 460080 288676 460086
rect 288624 460022 288676 460028
rect 288728 459785 288756 460255
rect 288714 459776 288770 459785
rect 288714 459711 288770 459720
rect 287702 459439 287758 459448
rect 287796 459468 287848 459474
rect 287520 458176 287572 458182
rect 287520 458118 287572 458124
rect 286230 456920 286286 456929
rect 286230 456855 286286 456864
rect 285588 442876 285640 442882
rect 285588 442818 285640 442824
rect 285496 442264 285548 442270
rect 285496 442206 285548 442212
rect 284944 441924 284996 441930
rect 284944 441866 284996 441872
rect 285770 333840 285826 333849
rect 285770 333775 285826 333784
rect 286966 333840 287022 333849
rect 286966 333775 287022 333784
rect 23032 333390 23152 333418
rect 22928 332444 22980 332450
rect 22928 332386 22980 332392
rect 22836 332376 22888 332382
rect 22836 332318 22888 332324
rect 22744 332036 22796 332042
rect 22744 331978 22796 331984
rect 22020 331906 22140 331922
rect 22020 331900 22152 331906
rect 22020 331894 22100 331900
rect 22100 331842 22152 331848
rect 22744 331900 22796 331906
rect 22744 331842 22796 331848
rect 22650 331800 22706 331809
rect 22650 331735 22706 331744
rect 21916 331288 21968 331294
rect 21916 331230 21968 331236
rect 21928 202842 21956 331230
rect 22664 325694 22692 331735
rect 22756 330834 22784 331842
rect 22848 331294 22876 332318
rect 22836 331288 22888 331294
rect 22836 331230 22888 331236
rect 22940 330970 22968 332386
rect 23032 332314 23060 333390
rect 285588 333328 285640 333334
rect 23124 333254 23460 333282
rect 28184 333254 28520 333282
rect 33244 333254 33580 333282
rect 38304 333254 38640 333282
rect 43364 333254 43700 333282
rect 48424 333254 48760 333282
rect 53484 333254 53820 333282
rect 58544 333254 58880 333282
rect 63604 333254 63940 333282
rect 68664 333254 69000 333282
rect 73172 333254 74060 333282
rect 78784 333254 79120 333282
rect 82832 333254 84180 333282
rect 88904 333266 89240 333282
rect 88892 333260 89240 333266
rect 23124 332518 23152 333254
rect 23664 332580 23716 332586
rect 23664 332522 23716 332528
rect 23112 332512 23164 332518
rect 23112 332454 23164 332460
rect 23020 332308 23072 332314
rect 23020 332250 23072 332256
rect 23032 331106 23060 332250
rect 23676 332246 23704 332522
rect 28184 332489 28212 333254
rect 28170 332480 28226 332489
rect 28170 332415 28226 332424
rect 33244 332314 33272 333254
rect 38304 332382 38332 333254
rect 43364 332450 43392 333254
rect 48424 332518 48452 333254
rect 48412 332512 48464 332518
rect 48412 332454 48464 332460
rect 43352 332444 43404 332450
rect 43352 332386 43404 332392
rect 38292 332376 38344 332382
rect 38292 332318 38344 332324
rect 33232 332308 33284 332314
rect 33232 332250 33284 332256
rect 23664 332240 23716 332246
rect 23664 332182 23716 332188
rect 53484 331906 53512 333254
rect 53472 331900 53524 331906
rect 53472 331842 53524 331848
rect 23032 331078 23336 331106
rect 22940 330942 23060 330970
rect 22756 330806 22968 330834
rect 22664 325666 22784 325694
rect 22008 315920 22060 315926
rect 22006 315888 22008 315897
rect 22060 315888 22062 315897
rect 22006 315823 22062 315832
rect 22006 204232 22062 204241
rect 22006 204167 22008 204176
rect 22060 204167 22062 204176
rect 22190 204232 22246 204241
rect 22190 204167 22246 204176
rect 22008 204138 22060 204144
rect 22204 203969 22232 204167
rect 22190 203960 22246 203969
rect 22190 203895 22246 203904
rect 22756 202881 22784 325666
rect 22742 202872 22798 202881
rect 21916 202836 21968 202842
rect 22742 202807 22798 202816
rect 21916 202778 21968 202784
rect 22940 202774 22968 330806
rect 23032 325694 23060 330942
rect 23032 325666 23244 325694
rect 23216 209774 23244 325666
rect 23032 209746 23244 209774
rect 23032 203969 23060 209746
rect 23308 203998 23336 331078
rect 23388 331016 23440 331022
rect 23386 330984 23388 330993
rect 23440 330984 23442 330993
rect 23386 330919 23442 330928
rect 58544 329730 58572 333254
rect 63604 332586 63632 333254
rect 63592 332580 63644 332586
rect 63592 332522 63644 332528
rect 68664 331809 68692 333254
rect 68650 331800 68706 331809
rect 68650 331735 68706 331744
rect 58532 329724 58584 329730
rect 58532 329666 58584 329672
rect 73172 315858 73200 333254
rect 78784 332926 78812 333254
rect 78772 332920 78824 332926
rect 78772 332862 78824 332868
rect 82832 315926 82860 333254
rect 88944 333254 89240 333260
rect 93872 333254 94300 333282
rect 99024 333254 99360 333282
rect 104084 333254 104420 333282
rect 109144 333254 109480 333282
rect 114204 333254 114540 333282
rect 119264 333254 119600 333282
rect 124324 333254 124660 333282
rect 129384 333254 129720 333282
rect 134444 333254 134780 333282
rect 139504 333254 139840 333282
rect 144840 333254 144900 333282
rect 149624 333254 149960 333282
rect 154684 333254 155020 333282
rect 160020 333254 160080 333282
rect 164252 333254 165140 333282
rect 170200 333254 170536 333282
rect 88892 333202 88944 333208
rect 82820 315920 82872 315926
rect 82820 315862 82872 315868
rect 73160 315852 73212 315858
rect 73160 315794 73212 315800
rect 93872 315314 93900 333254
rect 99024 331022 99052 333254
rect 99012 331016 99064 331022
rect 99012 330958 99064 330964
rect 104084 329798 104112 333254
rect 109144 332858 109172 333254
rect 109132 332852 109184 332858
rect 109132 332794 109184 332800
rect 114204 330886 114232 333254
rect 119264 331090 119292 333254
rect 124324 332790 124352 333254
rect 124312 332784 124364 332790
rect 124312 332726 124364 332732
rect 129384 332722 129412 333254
rect 129372 332716 129424 332722
rect 129372 332658 129424 332664
rect 134444 331294 134472 333254
rect 139504 332654 139532 333254
rect 139492 332648 139544 332654
rect 139492 332590 139544 332596
rect 144840 332586 144868 333254
rect 149624 332586 149652 333254
rect 144828 332580 144880 332586
rect 144828 332522 144880 332528
rect 149612 332580 149664 332586
rect 149612 332522 149664 332528
rect 149624 331809 149652 332522
rect 149610 331800 149666 331809
rect 149610 331735 149666 331744
rect 134432 331288 134484 331294
rect 134432 331230 134484 331236
rect 119252 331084 119304 331090
rect 119252 331026 119304 331032
rect 154684 330954 154712 333254
rect 160020 332466 160048 333254
rect 160020 332438 160140 332466
rect 160112 331226 160140 332438
rect 160100 331220 160152 331226
rect 160100 331162 160152 331168
rect 154672 330948 154724 330954
rect 154672 330890 154724 330896
rect 112444 330880 112496 330886
rect 112444 330822 112496 330828
rect 114192 330880 114244 330886
rect 114192 330822 114244 330828
rect 104072 329792 104124 329798
rect 104072 329734 104124 329740
rect 112456 315994 112484 330822
rect 160112 330449 160140 331162
rect 160098 330440 160154 330449
rect 160098 330375 160154 330384
rect 164252 318782 164280 333254
rect 170508 331294 170536 333254
rect 174924 333254 175260 333282
rect 179432 333254 180320 333282
rect 185380 333254 185716 333282
rect 174924 331294 174952 333254
rect 170496 331288 170548 331294
rect 170496 331230 170548 331236
rect 171784 331288 171836 331294
rect 171784 331230 171836 331236
rect 172336 331288 172388 331294
rect 172336 331230 172388 331236
rect 173808 331288 173860 331294
rect 173808 331230 173860 331236
rect 174912 331288 174964 331294
rect 174912 331230 174964 331236
rect 164240 318776 164292 318782
rect 164240 318718 164292 318724
rect 112444 315988 112496 315994
rect 112444 315930 112496 315936
rect 171796 315353 171824 331230
rect 172348 331158 172376 331230
rect 172336 331152 172388 331158
rect 172336 331094 172388 331100
rect 173820 317422 173848 331230
rect 173808 317416 173860 317422
rect 173808 317358 173860 317364
rect 179432 315994 179460 333254
rect 185688 331906 185716 333254
rect 190380 333254 190440 333282
rect 195500 333254 195928 333282
rect 190380 331974 190408 333254
rect 190368 331968 190420 331974
rect 190368 331910 190420 331916
rect 192116 331968 192168 331974
rect 192116 331910 192168 331916
rect 185676 331900 185728 331906
rect 185676 331842 185728 331848
rect 187608 331900 187660 331906
rect 187608 331842 187660 331848
rect 187620 330614 187648 331842
rect 187608 330608 187660 330614
rect 187608 330550 187660 330556
rect 192128 330546 192156 331910
rect 195900 331242 195928 333254
rect 200132 333254 200560 333282
rect 204272 333254 205620 333282
rect 210680 333254 211016 333282
rect 195900 331214 196020 331242
rect 192116 330540 192168 330546
rect 192116 330482 192168 330488
rect 195992 329118 196020 331214
rect 195980 329112 196032 329118
rect 195980 329054 196032 329060
rect 179420 315988 179472 315994
rect 179420 315930 179472 315936
rect 171782 315344 171838 315353
rect 93860 315308 93912 315314
rect 171782 315279 171838 315288
rect 93860 315250 93912 315256
rect 200132 313954 200160 333254
rect 204272 315353 204300 333254
rect 210988 332654 211016 333254
rect 215312 333254 215740 333282
rect 220740 333254 220800 333282
rect 224972 333254 225860 333282
rect 230920 333254 231256 333282
rect 210976 332648 211028 332654
rect 210976 332590 211028 332596
rect 215312 331242 215340 333254
rect 215220 331214 215340 331242
rect 220740 331242 220768 333254
rect 220740 331214 220860 331242
rect 215220 315926 215248 331214
rect 220832 331090 220860 331214
rect 220820 331084 220872 331090
rect 220820 331026 220872 331032
rect 215208 315920 215260 315926
rect 215208 315862 215260 315868
rect 224972 315858 225000 333254
rect 231228 332722 231256 333254
rect 234632 333254 235980 333282
rect 241040 333254 241376 333282
rect 246100 333254 246436 333282
rect 231216 332716 231268 332722
rect 231216 332658 231268 332664
rect 224960 315852 225012 315858
rect 224960 315794 225012 315800
rect 234632 315790 234660 333254
rect 241348 332489 241376 333254
rect 246408 332586 246436 333254
rect 251100 333254 251160 333282
rect 256220 333254 256556 333282
rect 261280 333254 261616 333282
rect 246396 332580 246448 332586
rect 246396 332522 246448 332528
rect 251100 332518 251128 333254
rect 251088 332512 251140 332518
rect 241334 332480 241390 332489
rect 251088 332454 251140 332460
rect 256528 332450 256556 333254
rect 241334 332415 241390 332424
rect 256516 332444 256568 332450
rect 256516 332386 256568 332392
rect 261588 332382 261616 333254
rect 266280 333254 266340 333282
rect 270512 333254 271400 333282
rect 276032 333254 276460 333282
rect 281460 333254 281520 333282
rect 285588 333270 285640 333276
rect 284208 333260 284260 333266
rect 261576 332376 261628 332382
rect 261576 332318 261628 332324
rect 266280 332314 266308 333254
rect 266268 332308 266320 332314
rect 266268 332250 266320 332256
rect 234620 315784 234672 315790
rect 234620 315726 234672 315732
rect 204258 315344 204314 315353
rect 270512 315314 270540 333254
rect 276032 315382 276060 333254
rect 281460 332450 281488 333254
rect 284208 333202 284260 333208
rect 281356 332444 281408 332450
rect 281356 332386 281408 332392
rect 281448 332444 281500 332450
rect 281448 332386 281500 332392
rect 281368 332246 281396 332386
rect 282184 332376 282236 332382
rect 282184 332318 282236 332324
rect 281356 332240 281408 332246
rect 281356 332182 281408 332188
rect 282196 331906 282224 332318
rect 282184 331900 282236 331906
rect 282184 331842 282236 331848
rect 284220 318782 284248 333202
rect 285496 330608 285548 330614
rect 285496 330550 285548 330556
rect 285508 330002 285536 330550
rect 285496 329996 285548 330002
rect 285496 329938 285548 329944
rect 284208 318776 284260 318782
rect 284260 318724 284340 318730
rect 284208 318718 284340 318724
rect 284220 318702 284340 318718
rect 284220 318653 284248 318702
rect 276020 315376 276072 315382
rect 276020 315318 276072 315324
rect 204258 315279 204314 315288
rect 270500 315308 270552 315314
rect 270500 315250 270552 315256
rect 284312 314022 284340 318702
rect 285404 317416 285456 317422
rect 285404 317358 285456 317364
rect 285416 316713 285444 317358
rect 285402 316704 285458 316713
rect 285402 316639 285458 316648
rect 285508 314090 285536 329938
rect 285600 315994 285628 333270
rect 285680 332240 285732 332246
rect 285678 332208 285680 332217
rect 285732 332208 285734 332217
rect 285678 332143 285734 332152
rect 285784 331158 285812 333775
rect 286874 333704 286930 333713
rect 286874 333639 286930 333648
rect 286580 333254 286732 333282
rect 286704 331265 286732 333254
rect 286690 331256 286746 331265
rect 286690 331191 286746 331200
rect 285772 331152 285824 331158
rect 285772 331094 285824 331100
rect 286888 330002 286916 333639
rect 286876 329996 286928 330002
rect 286876 329938 286928 329944
rect 285588 315988 285640 315994
rect 285588 315930 285640 315936
rect 285600 315450 285628 315930
rect 286980 315489 287008 333775
rect 287532 315858 287560 458118
rect 287610 458008 287666 458017
rect 287610 457943 287666 457952
rect 287624 332654 287652 457943
rect 287612 332648 287664 332654
rect 287612 332590 287664 332596
rect 287520 315852 287572 315858
rect 287520 315794 287572 315800
rect 286966 315480 287022 315489
rect 285588 315444 285640 315450
rect 286966 315415 287022 315424
rect 285588 315386 285640 315392
rect 285496 314084 285548 314090
rect 285496 314026 285548 314032
rect 284300 314016 284352 314022
rect 284300 313958 284352 313964
rect 200120 313948 200172 313954
rect 200120 313890 200172 313896
rect 285496 205964 285548 205970
rect 285496 205906 285548 205912
rect 23846 205864 23902 205873
rect 23846 205799 23902 205808
rect 23754 205728 23810 205737
rect 23584 205686 23754 205714
rect 23400 205278 23460 205306
rect 23296 203992 23348 203998
rect 23018 203960 23074 203969
rect 23018 203895 23074 203904
rect 23202 203960 23258 203969
rect 23296 203934 23348 203940
rect 23202 203895 23258 203904
rect 23112 202836 23164 202842
rect 23112 202778 23164 202784
rect 22928 202768 22980 202774
rect 22926 202736 22928 202745
rect 22980 202736 22982 202745
rect 21824 202700 21876 202706
rect 22926 202671 22982 202680
rect 21824 202642 21876 202648
rect 21732 202632 21784 202638
rect 21732 202574 21784 202580
rect 21744 74390 21772 202574
rect 21836 75682 21864 202642
rect 23124 202230 23152 202778
rect 23112 202224 23164 202230
rect 23112 202166 23164 202172
rect 22008 199436 22060 199442
rect 22008 199378 22060 199384
rect 22020 199102 22048 199378
rect 22008 199096 22060 199102
rect 22008 199038 22060 199044
rect 21824 75676 21876 75682
rect 21824 75618 21876 75624
rect 21732 74384 21784 74390
rect 21732 74326 21784 74332
rect 22020 71602 22048 199038
rect 23020 185904 23072 185910
rect 23020 185846 23072 185852
rect 23032 77926 23060 185846
rect 23020 77920 23072 77926
rect 23020 77862 23072 77868
rect 23124 74254 23152 202166
rect 23216 74322 23244 203895
rect 23204 74316 23256 74322
rect 23204 74258 23256 74264
rect 23112 74248 23164 74254
rect 23112 74190 23164 74196
rect 23308 74186 23336 203934
rect 23400 203930 23428 205278
rect 23388 203924 23440 203930
rect 23388 203866 23440 203872
rect 23388 202836 23440 202842
rect 23388 202778 23440 202784
rect 23400 202638 23428 202778
rect 23388 202632 23440 202638
rect 23388 202574 23440 202580
rect 23584 200122 23612 205686
rect 23754 205663 23810 205672
rect 23572 200116 23624 200122
rect 23860 200114 23888 205799
rect 284942 205728 284998 205737
rect 284942 205663 284998 205672
rect 28184 205278 28520 205306
rect 33244 205278 33580 205306
rect 38304 205278 38640 205306
rect 43364 205278 43700 205306
rect 48424 205278 48760 205306
rect 53484 205278 53820 205306
rect 58544 205278 58880 205306
rect 63604 205278 63940 205306
rect 68664 205278 69000 205306
rect 73724 205278 74060 205306
rect 78784 205278 79120 205306
rect 83844 205278 84180 205306
rect 88904 205278 89240 205306
rect 94056 205278 94300 205306
rect 99024 205278 99360 205306
rect 104084 205278 104420 205306
rect 109052 205278 109480 205306
rect 113192 205278 114540 205306
rect 119264 205278 119600 205306
rect 124232 205278 124660 205306
rect 128372 205278 129720 205306
rect 134444 205278 134780 205306
rect 139412 205278 139840 205306
rect 144840 205278 144900 205306
rect 149624 205278 149960 205306
rect 154684 205278 155020 205306
rect 158732 205278 160080 205306
rect 165140 205278 165476 205306
rect 170200 205278 170536 205306
rect 28184 204105 28212 205278
rect 28170 204096 28226 204105
rect 28170 204031 28226 204040
rect 33244 203998 33272 205278
rect 38304 203998 38332 205278
rect 33232 203992 33284 203998
rect 33232 203934 33284 203940
rect 33324 203992 33376 203998
rect 33324 203934 33376 203940
rect 38292 203992 38344 203998
rect 43364 203969 43392 205278
rect 38292 203934 38344 203940
rect 43350 203960 43406 203969
rect 33336 202230 33364 203934
rect 43350 203895 43406 203904
rect 48424 202706 48452 205278
rect 53484 202774 53512 205278
rect 58544 203590 58572 205278
rect 58532 203584 58584 203590
rect 58532 203526 58584 203532
rect 63604 202842 63632 205278
rect 68664 202881 68692 205278
rect 73724 204066 73752 205278
rect 78784 204134 78812 205278
rect 83844 204202 83872 205278
rect 88904 204270 88932 205278
rect 88892 204264 88944 204270
rect 94056 204241 94084 205278
rect 88892 204206 88944 204212
rect 94042 204232 94098 204241
rect 83832 204196 83884 204202
rect 94042 204167 94098 204176
rect 83832 204138 83884 204144
rect 78772 204128 78824 204134
rect 78772 204070 78824 204076
rect 73712 204060 73764 204066
rect 73712 204002 73764 204008
rect 99024 203522 99052 205278
rect 96620 203516 96672 203522
rect 96620 203458 96672 203464
rect 99012 203516 99064 203522
rect 99012 203458 99064 203464
rect 68650 202872 68706 202881
rect 63592 202836 63644 202842
rect 68650 202807 68706 202816
rect 63592 202778 63644 202784
rect 53472 202768 53524 202774
rect 53472 202710 53524 202716
rect 48412 202700 48464 202706
rect 48412 202642 48464 202648
rect 33324 202224 33376 202230
rect 24858 202192 24914 202201
rect 96632 202201 96660 203458
rect 103520 202904 103572 202910
rect 103440 202852 103520 202874
rect 103440 202846 103572 202852
rect 33324 202166 33376 202172
rect 96618 202192 96674 202201
rect 24858 202127 24914 202136
rect 96618 202127 96674 202136
rect 24124 200796 24176 200802
rect 24124 200738 24176 200744
rect 23572 200058 23624 200064
rect 23676 200086 23888 200114
rect 23584 199510 23612 200058
rect 23572 199504 23624 199510
rect 23572 199446 23624 199452
rect 23676 189038 23704 200086
rect 23664 189032 23716 189038
rect 23664 188974 23716 188980
rect 23676 187746 23704 188974
rect 23664 187740 23716 187746
rect 23664 187682 23716 187688
rect 24136 185910 24164 200738
rect 24872 186425 24900 202127
rect 103440 199918 103468 202846
rect 104084 202842 104112 205278
rect 104072 202836 104124 202842
rect 104072 202778 104124 202784
rect 103428 199912 103480 199918
rect 103428 199854 103480 199860
rect 109052 199442 109080 205278
rect 109040 199436 109092 199442
rect 109040 199378 109092 199384
rect 113192 188970 113220 205278
rect 119264 204474 119292 205278
rect 119252 204468 119304 204474
rect 119252 204410 119304 204416
rect 113180 188964 113232 188970
rect 113180 188906 113232 188912
rect 24858 186416 24914 186425
rect 24858 186351 24914 186360
rect 124232 186017 124260 205278
rect 128372 199986 128400 205278
rect 134444 204542 134472 205278
rect 134432 204536 134484 204542
rect 134432 204478 134484 204484
rect 139412 200054 139440 205278
rect 144840 204270 144868 205278
rect 149624 204270 149652 205278
rect 154684 204406 154712 205278
rect 154672 204400 154724 204406
rect 154672 204342 154724 204348
rect 144828 204264 144880 204270
rect 144828 204206 144880 204212
rect 149612 204264 149664 204270
rect 149612 204206 149664 204212
rect 149624 203590 149652 204206
rect 149612 203584 149664 203590
rect 149612 203526 149664 203532
rect 158732 200122 158760 205278
rect 165448 202910 165476 205278
rect 170508 203114 170536 205278
rect 175200 205278 175260 205306
rect 180260 205278 180320 205306
rect 185320 205278 185380 205306
rect 190380 205278 190440 205306
rect 195500 205278 195836 205306
rect 175200 204270 175228 205278
rect 180260 204610 180288 205278
rect 180248 204604 180300 204610
rect 180248 204546 180300 204552
rect 173900 204264 173952 204270
rect 173900 204206 173952 204212
rect 175188 204264 175240 204270
rect 175188 204206 175240 204212
rect 170496 203108 170548 203114
rect 170496 203050 170548 203056
rect 171140 203108 171192 203114
rect 171140 203050 171192 203056
rect 165436 202904 165488 202910
rect 165436 202846 165488 202852
rect 166264 202904 166316 202910
rect 166264 202846 166316 202852
rect 158720 200116 158772 200122
rect 158720 200058 158772 200064
rect 139400 200048 139452 200054
rect 139400 199990 139452 199996
rect 128360 199980 128412 199986
rect 128360 199922 128412 199928
rect 166276 198014 166304 202846
rect 166264 198008 166316 198014
rect 166264 197950 166316 197956
rect 171152 189038 171180 203050
rect 171140 189032 171192 189038
rect 171140 188974 171192 188980
rect 124218 186008 124274 186017
rect 124218 185943 124274 185952
rect 173912 185910 173940 204206
rect 175200 202858 175228 204206
rect 175200 202830 175320 202858
rect 175292 202774 175320 202830
rect 175280 202768 175332 202774
rect 175280 202710 175332 202716
rect 185320 201482 185348 205278
rect 190380 204134 190408 205278
rect 190368 204128 190420 204134
rect 190368 204070 190420 204076
rect 192484 204128 192536 204134
rect 192484 204070 192536 204076
rect 185308 201476 185360 201482
rect 185308 201418 185360 201424
rect 185320 200802 185348 201418
rect 185308 200796 185360 200802
rect 185308 200738 185360 200744
rect 192496 186318 192524 204070
rect 195808 202706 195836 205278
rect 200132 205278 200560 205306
rect 204272 205278 205620 205306
rect 210680 205278 211016 205306
rect 215740 205278 216076 205306
rect 195796 202700 195848 202706
rect 195796 202642 195848 202648
rect 192484 186312 192536 186318
rect 192484 186254 192536 186260
rect 200132 185910 200160 205278
rect 204272 188329 204300 205278
rect 210988 200802 211016 205278
rect 216048 201414 216076 205278
rect 220740 205278 220800 205306
rect 225860 205278 226196 205306
rect 230920 205278 231256 205306
rect 220740 204406 220768 205278
rect 220728 204400 220780 204406
rect 220728 204342 220780 204348
rect 226168 202638 226196 205278
rect 226156 202632 226208 202638
rect 226156 202574 226208 202580
rect 216036 201408 216088 201414
rect 216036 201350 216088 201356
rect 231228 201346 231256 205278
rect 235920 205278 235980 205306
rect 241040 205278 241376 205306
rect 246100 205278 246436 205306
rect 235920 204474 235948 205278
rect 241348 204542 241376 205278
rect 246408 204610 246436 205278
rect 251100 205278 251160 205306
rect 256220 205278 256556 205306
rect 261280 205278 261616 205306
rect 246396 204604 246448 204610
rect 246396 204546 246448 204552
rect 241336 204536 241388 204542
rect 241336 204478 241388 204484
rect 235908 204468 235960 204474
rect 235908 204410 235960 204416
rect 251100 204270 251128 205278
rect 251088 204264 251140 204270
rect 251088 204206 251140 204212
rect 256528 204202 256556 205278
rect 256516 204196 256568 204202
rect 256516 204138 256568 204144
rect 261588 203658 261616 205278
rect 266280 205278 266340 205306
rect 271400 205278 271736 205306
rect 266280 203726 266308 205278
rect 266268 203720 266320 203726
rect 266268 203662 266320 203668
rect 261576 203652 261628 203658
rect 261576 203594 261628 203600
rect 271708 203561 271736 205278
rect 276032 205278 276460 205306
rect 281460 205278 281520 205306
rect 271694 203552 271750 203561
rect 271694 203487 271750 203496
rect 231216 201340 231268 201346
rect 231216 201282 231268 201288
rect 210976 200796 211028 200802
rect 210976 200738 211028 200744
rect 204258 188320 204314 188329
rect 204258 188255 204314 188264
rect 276032 186998 276060 205278
rect 281460 203930 281488 205278
rect 281448 203924 281500 203930
rect 281448 203866 281500 203872
rect 284956 202706 284984 205663
rect 284944 202700 284996 202706
rect 284944 202642 284996 202648
rect 276020 186992 276072 186998
rect 276020 186934 276072 186940
rect 284956 186017 284984 202642
rect 285508 187066 285536 205906
rect 285770 205864 285826 205873
rect 285770 205799 285826 205808
rect 285588 204944 285640 204950
rect 285588 204886 285640 204892
rect 285496 187060 285548 187066
rect 285496 187002 285548 187008
rect 285600 186318 285628 204886
rect 285680 204196 285732 204202
rect 285680 204138 285732 204144
rect 285692 203697 285720 204138
rect 285678 203688 285734 203697
rect 285678 203623 285734 203632
rect 285784 202774 285812 205799
rect 286580 205278 286824 205306
rect 286796 203794 286824 205278
rect 286966 204912 287022 204921
rect 286966 204847 287022 204856
rect 286784 203788 286836 203794
rect 286784 203730 286836 203736
rect 285772 202768 285824 202774
rect 285772 202710 285824 202716
rect 285680 200796 285732 200802
rect 285680 200738 285732 200744
rect 285692 200190 285720 200738
rect 285680 200184 285732 200190
rect 285680 200126 285732 200132
rect 286876 200184 286928 200190
rect 286876 200126 286928 200132
rect 285128 186312 285180 186318
rect 285128 186254 285180 186260
rect 285588 186312 285640 186318
rect 285588 186254 285640 186260
rect 284942 186008 284998 186017
rect 284942 185943 284998 185952
rect 24124 185904 24176 185910
rect 24124 185846 24176 185852
rect 173900 185904 173952 185910
rect 173900 185846 173952 185852
rect 200120 185904 200172 185910
rect 285140 185881 285168 186254
rect 286888 185978 286916 200126
rect 286980 186153 287008 204847
rect 287532 202638 287560 315794
rect 287520 202632 287572 202638
rect 287520 202574 287572 202580
rect 287532 190454 287560 202574
rect 287624 200190 287652 332590
rect 287716 332450 287744 459439
rect 287796 459410 287848 459416
rect 288532 458992 288584 458998
rect 288532 458934 288584 458940
rect 288440 458856 288492 458862
rect 288440 458798 288492 458804
rect 287704 332444 287756 332450
rect 287704 332386 287756 332392
rect 287716 203930 287744 332386
rect 287888 204468 287940 204474
rect 287888 204410 287940 204416
rect 287704 203924 287756 203930
rect 287704 203866 287756 203872
rect 287612 200184 287664 200190
rect 287612 200126 287664 200132
rect 287532 190426 287836 190454
rect 287520 189780 287572 189786
rect 287520 189722 287572 189728
rect 286966 186144 287022 186153
rect 286966 186079 287022 186088
rect 286876 185972 286928 185978
rect 286876 185914 286928 185920
rect 200120 185846 200172 185852
rect 285126 185872 285182 185881
rect 285126 185807 285182 185816
rect 25504 77920 25556 77926
rect 114192 77920 114244 77926
rect 25504 77862 25556 77868
rect 25594 77888 25650 77897
rect 23400 77302 23460 77330
rect 23400 75614 23428 77302
rect 23480 77104 23532 77110
rect 23480 77046 23532 77052
rect 23388 75608 23440 75614
rect 23388 75550 23440 75556
rect 23296 74180 23348 74186
rect 23296 74122 23348 74128
rect 23492 72962 23520 77046
rect 23480 72956 23532 72962
rect 23480 72898 23532 72904
rect 22008 71596 22060 71602
rect 22008 71538 22060 71544
rect 25516 69018 25544 77862
rect 193220 77920 193272 77926
rect 114244 77868 114540 77874
rect 114192 77862 114540 77868
rect 240784 77920 240836 77926
rect 193220 77862 193272 77868
rect 194598 77888 194654 77897
rect 114204 77846 114540 77862
rect 25594 77823 25650 77832
rect 25608 71670 25636 77823
rect 28184 77302 28520 77330
rect 33580 77302 33732 77330
rect 28184 76158 28212 77302
rect 28172 76152 28224 76158
rect 28172 76094 28224 76100
rect 33704 74186 33732 77302
rect 37936 77302 38640 77330
rect 43456 77302 43700 77330
rect 48760 77302 49096 77330
rect 37936 74254 37964 77302
rect 43456 74322 43484 77302
rect 49068 75682 49096 77302
rect 53806 77081 53834 77316
rect 58880 77302 59308 77330
rect 63940 77302 64184 77330
rect 52458 77072 52514 77081
rect 52458 77007 52514 77016
rect 53792 77072 53848 77081
rect 53792 77007 53848 77016
rect 52472 75993 52500 77007
rect 52458 75984 52514 75993
rect 52458 75919 52514 75928
rect 49056 75676 49108 75682
rect 49056 75618 49108 75624
rect 49068 75206 49096 75618
rect 49056 75200 49108 75206
rect 49056 75142 49108 75148
rect 43444 74316 43496 74322
rect 43444 74258 43496 74264
rect 37924 74248 37976 74254
rect 37924 74190 37976 74196
rect 33692 74180 33744 74186
rect 33692 74122 33744 74128
rect 25596 71664 25648 71670
rect 25596 71606 25648 71612
rect 33704 71058 33732 74122
rect 33692 71052 33744 71058
rect 33692 70994 33744 71000
rect 25504 69012 25556 69018
rect 25504 68954 25556 68960
rect 37936 57390 37964 74190
rect 40684 69692 40736 69698
rect 40684 69634 40736 69640
rect 40696 64326 40724 69634
rect 40684 64320 40736 64326
rect 40684 64262 40736 64268
rect 43456 61402 43484 74258
rect 52472 61470 52500 75919
rect 59280 75750 59308 77302
rect 59268 75744 59320 75750
rect 59268 75686 59320 75692
rect 59280 69766 59308 75686
rect 64156 74390 64184 77302
rect 68664 77302 69000 77330
rect 73816 77302 74060 77330
rect 79120 77302 79456 77330
rect 68664 74534 68692 77302
rect 73816 75818 73844 77302
rect 73804 75812 73856 75818
rect 73804 75754 73856 75760
rect 68296 74506 68692 74534
rect 68296 74458 68324 74506
rect 68284 74452 68336 74458
rect 68284 74394 68336 74400
rect 64144 74384 64196 74390
rect 64144 74326 64196 74332
rect 59268 69760 59320 69766
rect 59268 69702 59320 69708
rect 52460 61464 52512 61470
rect 52460 61406 52512 61412
rect 43444 61396 43496 61402
rect 43444 61338 43496 61344
rect 37924 57384 37976 57390
rect 37924 57326 37976 57332
rect 64156 57322 64184 74326
rect 68296 58682 68324 74394
rect 73816 66978 73844 75754
rect 79428 75585 79456 77302
rect 84120 77302 84180 77330
rect 88996 77302 89240 77330
rect 84120 75721 84148 77302
rect 88996 75886 89024 77302
rect 94286 77058 94314 77316
rect 98656 77302 99360 77330
rect 104176 77302 104420 77330
rect 109144 77302 109480 77330
rect 94286 77030 94360 77058
rect 88984 75880 89036 75886
rect 88984 75822 89036 75828
rect 84106 75712 84162 75721
rect 84106 75647 84162 75656
rect 79414 75576 79470 75585
rect 79414 75511 79470 75520
rect 79428 73982 79456 75511
rect 79416 73976 79468 73982
rect 79416 73918 79468 73924
rect 84120 68406 84148 75647
rect 84108 68400 84160 68406
rect 84108 68342 84160 68348
rect 73804 66972 73856 66978
rect 73804 66914 73856 66920
rect 88996 58750 89024 75822
rect 94332 74526 94360 77030
rect 98656 75857 98684 77302
rect 98642 75848 98698 75857
rect 98642 75783 98698 75792
rect 94320 74520 94372 74526
rect 94320 74462 94372 74468
rect 94332 71126 94360 74462
rect 94320 71120 94372 71126
rect 94320 71062 94372 71068
rect 98656 60042 98684 75783
rect 104176 74497 104204 77302
rect 104162 74488 104218 74497
rect 104162 74423 104218 74432
rect 104176 60110 104204 74423
rect 109144 71602 109172 77302
rect 109132 71596 109184 71602
rect 109132 71538 109184 71544
rect 109144 70446 109172 71538
rect 114480 71194 114508 77846
rect 119600 77302 119936 77330
rect 119908 76090 119936 77302
rect 124600 77302 124660 77330
rect 129384 77302 129720 77330
rect 134444 77302 134780 77330
rect 139840 77302 140084 77330
rect 119896 76084 119948 76090
rect 119896 76026 119948 76032
rect 116584 75200 116636 75206
rect 116584 75142 116636 75148
rect 114468 71188 114520 71194
rect 114468 71130 114520 71136
rect 109132 70440 109184 70446
rect 109132 70382 109184 70388
rect 109684 70440 109736 70446
rect 109684 70382 109736 70388
rect 109696 60178 109724 70382
rect 116596 61538 116624 75142
rect 119908 73914 119936 76026
rect 119896 73908 119948 73914
rect 119896 73850 119948 73856
rect 124600 71670 124628 77302
rect 129384 74534 129412 77302
rect 134444 75954 134472 77302
rect 134432 75948 134484 75954
rect 134432 75890 134484 75896
rect 129016 74506 129412 74534
rect 129016 71777 129044 74506
rect 134444 72622 134472 75890
rect 134432 72616 134484 72622
rect 134432 72558 134484 72564
rect 129002 71768 129058 71777
rect 140056 71738 140084 77302
rect 144840 77302 144900 77330
rect 149624 77302 149960 77330
rect 155020 77302 155264 77330
rect 144840 75886 144868 77302
rect 149624 75886 149652 77302
rect 153016 76560 153068 76566
rect 151726 76528 151782 76537
rect 153016 76502 153068 76508
rect 151726 76463 151782 76472
rect 144828 75880 144880 75886
rect 144828 75822 144880 75828
rect 149612 75880 149664 75886
rect 149612 75822 149664 75828
rect 149980 75880 150032 75886
rect 149980 75822 150032 75828
rect 129002 71703 129058 71712
rect 140044 71732 140096 71738
rect 124588 71664 124640 71670
rect 124588 71606 124640 71612
rect 125508 71664 125560 71670
rect 125508 71606 125560 71612
rect 125520 69834 125548 71606
rect 125508 69828 125560 69834
rect 125508 69770 125560 69776
rect 116584 61532 116636 61538
rect 116584 61474 116636 61480
rect 109684 60172 109736 60178
rect 109684 60114 109736 60120
rect 104164 60104 104216 60110
rect 104164 60046 104216 60052
rect 98644 60036 98696 60042
rect 98644 59978 98696 59984
rect 88984 58744 89036 58750
rect 88984 58686 89036 58692
rect 68284 58676 68336 58682
rect 68284 58618 68336 58624
rect 129016 57458 129044 71703
rect 140044 71674 140096 71680
rect 140056 58818 140084 71674
rect 149992 68542 150020 75822
rect 149980 68536 150032 68542
rect 149980 68478 150032 68484
rect 140044 58812 140096 58818
rect 140044 58754 140096 58760
rect 129004 57452 129056 57458
rect 129004 57394 129056 57400
rect 64144 57316 64196 57322
rect 64144 57258 64196 57264
rect 151634 53136 151690 53145
rect 151084 53100 151136 53106
rect 151084 53042 151136 53048
rect 151544 53100 151596 53106
rect 151634 53071 151690 53080
rect 151544 53042 151596 53048
rect 150440 51060 150492 51066
rect 150440 51002 150492 51008
rect 150452 50561 150480 51002
rect 150438 50552 150494 50561
rect 150438 50487 150494 50496
rect 150440 49700 150492 49706
rect 150440 49642 150492 49648
rect 150452 49609 150480 49642
rect 150438 49600 150494 49609
rect 150438 49535 150494 49544
rect 150440 48272 150492 48278
rect 150438 48240 150440 48249
rect 150492 48240 150494 48249
rect 21364 48204 21416 48210
rect 150438 48175 150494 48184
rect 150532 48204 150584 48210
rect 21364 48146 21416 48152
rect 150532 48146 150584 48152
rect 150544 47705 150572 48146
rect 150530 47696 150586 47705
rect 150530 47631 150586 47640
rect 150440 46912 150492 46918
rect 150440 46854 150492 46860
rect 150452 46753 150480 46854
rect 150438 46744 150494 46753
rect 150438 46679 150494 46688
rect 150440 45552 150492 45558
rect 151096 45529 151124 53042
rect 150440 45494 150492 45500
rect 151082 45520 151138 45529
rect 150452 44849 150480 45494
rect 151082 45455 151138 45464
rect 150438 44840 150494 44849
rect 150438 44775 150494 44784
rect 150440 44124 150492 44130
rect 150440 44066 150492 44072
rect 150452 43897 150480 44066
rect 150438 43888 150494 43897
rect 150438 43823 150494 43832
rect 150440 42764 150492 42770
rect 150440 42706 150492 42712
rect 150452 42537 150480 42706
rect 150438 42528 150494 42537
rect 150438 42463 150494 42472
rect 150440 41404 150492 41410
rect 150440 41346 150492 41352
rect 150452 41313 150480 41346
rect 150438 41304 150494 41313
rect 150438 41239 150494 41248
rect 151556 39953 151584 53042
rect 151542 39944 151598 39953
rect 151542 39879 151598 39888
rect 151176 39364 151228 39370
rect 151176 39306 151228 39312
rect 151084 36576 151136 36582
rect 151084 36518 151136 36524
rect 16488 35896 16540 35902
rect 150440 35896 150492 35902
rect 16488 35838 16540 35844
rect 150438 35864 150440 35873
rect 150492 35864 150494 35873
rect 150438 35799 150494 35808
rect 15844 34468 15896 34474
rect 15844 34410 15896 34416
rect 150440 34468 150492 34474
rect 150440 34410 150492 34416
rect 150452 34377 150480 34410
rect 150438 34368 150494 34377
rect 150438 34303 150494 34312
rect 7656 33108 7708 33114
rect 7656 33050 7708 33056
rect 150440 33108 150492 33114
rect 150440 33050 150492 33056
rect 150452 32473 150480 33050
rect 150438 32464 150494 32473
rect 150438 32399 150494 32408
rect 150440 31748 150492 31754
rect 150440 31690 150492 31696
rect 150452 31521 150480 31690
rect 150438 31512 150494 31521
rect 150438 31447 150494 31456
rect 150440 30320 150492 30326
rect 150440 30262 150492 30268
rect 150452 30161 150480 30262
rect 150438 30152 150494 30161
rect 150438 30087 150494 30096
rect 5080 28960 5132 28966
rect 150440 28960 150492 28966
rect 5080 28902 5132 28908
rect 150438 28928 150440 28937
rect 150492 28928 150494 28937
rect 150438 28863 150494 28872
rect 151096 28529 151124 36518
rect 151188 33153 151216 39306
rect 151648 37233 151676 53071
rect 151740 38185 151768 76463
rect 153028 40429 153056 76502
rect 153108 75948 153160 75954
rect 153108 75890 153160 75896
rect 153014 40420 153070 40429
rect 153014 40355 153070 40364
rect 153120 38729 153148 75890
rect 155236 72894 155264 77302
rect 159744 77302 160080 77330
rect 164804 77302 165140 77330
rect 169772 77302 170200 77330
rect 174924 77302 175260 77330
rect 180076 77302 180320 77330
rect 184952 77302 185380 77330
rect 190380 77302 190440 77330
rect 159744 74534 159772 77302
rect 159376 74506 159772 74534
rect 159376 73030 159404 74506
rect 159364 73024 159416 73030
rect 159364 72966 159416 72972
rect 155224 72888 155276 72894
rect 155224 72830 155276 72836
rect 154672 62892 154724 62898
rect 154672 62834 154724 62840
rect 154684 52714 154712 62834
rect 155236 53854 155264 72830
rect 156512 62824 156564 62830
rect 156512 62766 156564 62772
rect 155224 53848 155276 53854
rect 155224 53790 155276 53796
rect 156524 52714 156552 62766
rect 158720 54528 158772 54534
rect 158720 54470 158772 54476
rect 154684 52686 155066 52714
rect 156524 52686 156906 52714
rect 158732 52700 158760 54470
rect 159376 54466 159404 72966
rect 164240 72956 164292 72962
rect 164240 72898 164292 72904
rect 164252 72486 164280 72898
rect 164804 72486 164832 77302
rect 169772 76022 169800 77302
rect 169760 76016 169812 76022
rect 169760 75958 169812 75964
rect 164240 72480 164292 72486
rect 164240 72422 164292 72428
rect 164792 72480 164844 72486
rect 164792 72422 164844 72428
rect 159364 54460 159416 54466
rect 159364 54402 159416 54408
rect 162400 54460 162452 54466
rect 162400 54402 162452 54408
rect 160560 53848 160612 53854
rect 160560 53790 160612 53796
rect 160572 52700 160600 53790
rect 162412 52700 162440 54402
rect 164252 52700 164280 72422
rect 169772 56030 169800 75958
rect 174924 74534 174952 77302
rect 174556 74506 174952 74534
rect 174556 73098 174584 74506
rect 180076 73166 180104 77302
rect 180064 73160 180116 73166
rect 180064 73102 180116 73108
rect 174544 73092 174596 73098
rect 174544 73034 174596 73040
rect 169852 72480 169904 72486
rect 169852 72422 169904 72428
rect 169760 56024 169812 56030
rect 169760 55966 169812 55972
rect 166080 55956 166132 55962
rect 166080 55898 166132 55904
rect 166092 52700 166120 55898
rect 167920 55888 167972 55894
rect 167920 55830 167972 55836
rect 167932 52700 167960 55830
rect 169864 52714 169892 72422
rect 173072 64252 173124 64258
rect 173072 64194 173124 64200
rect 171600 54596 171652 54602
rect 171600 54538 171652 54544
rect 169786 52686 169892 52714
rect 171612 52700 171640 54538
rect 173084 52714 173112 64194
rect 174556 54738 174584 73034
rect 178684 64320 178736 64326
rect 178684 64262 178736 64268
rect 175280 64184 175332 64190
rect 175280 64126 175332 64132
rect 174544 54732 174596 54738
rect 174544 54674 174596 54680
rect 173084 52686 173466 52714
rect 175292 52700 175320 64126
rect 178696 54806 178724 64262
rect 178960 56024 179012 56030
rect 178960 55966 179012 55972
rect 178684 54800 178736 54806
rect 178684 54742 178736 54748
rect 178972 52700 179000 55966
rect 180076 54670 180104 73102
rect 184952 69018 184980 77302
rect 190380 75886 190408 77302
rect 188344 75880 188396 75886
rect 188344 75822 188396 75828
rect 190368 75880 190420 75886
rect 190368 75822 190420 75828
rect 184940 69012 184992 69018
rect 184940 68954 184992 68960
rect 184952 55214 184980 68954
rect 187792 65544 187844 65550
rect 187792 65486 187844 65492
rect 184860 55186 184980 55214
rect 180800 54732 180852 54738
rect 180800 54674 180852 54680
rect 180064 54664 180116 54670
rect 180064 54606 180116 54612
rect 180812 52700 180840 54674
rect 182640 54664 182692 54670
rect 182640 54606 182692 54612
rect 182652 52700 182680 54606
rect 184860 52714 184888 55186
rect 186320 53848 186372 53854
rect 186320 53790 186372 53796
rect 184506 52686 184888 52714
rect 186332 52700 186360 53790
rect 187804 52714 187832 65486
rect 188356 53854 188384 75822
rect 191840 75200 191892 75206
rect 191840 75142 191892 75148
rect 188344 53848 188396 53854
rect 188344 53790 188396 53796
rect 187804 52686 188186 52714
rect 191852 52700 191880 75142
rect 193232 74534 193260 77862
rect 195794 77888 195850 77897
rect 195500 77846 195794 77874
rect 194598 77823 194654 77832
rect 240784 77862 240836 77868
rect 284944 77920 284996 77926
rect 284944 77862 284996 77868
rect 195794 77823 195850 77832
rect 193232 74506 193352 74534
rect 193324 52714 193352 74506
rect 194612 65550 194640 77823
rect 200408 77302 200560 77330
rect 204272 77302 205620 77330
rect 209792 77302 210680 77330
rect 215740 77302 216076 77330
rect 200304 76016 200356 76022
rect 200304 75958 200356 75964
rect 200316 74534 200344 75958
rect 200408 75206 200436 77302
rect 200396 75200 200448 75206
rect 200396 75142 200448 75148
rect 200316 74506 200712 74534
rect 195152 68604 195204 68610
rect 195152 68546 195204 68552
rect 194600 65544 194652 65550
rect 194600 65486 194652 65492
rect 195164 52714 195192 68546
rect 198830 68232 198886 68241
rect 198830 68167 198886 68176
rect 197360 54664 197412 54670
rect 197360 54606 197412 54612
rect 193324 52686 193706 52714
rect 195164 52686 195546 52714
rect 197372 52700 197400 54606
rect 198844 52714 198872 68167
rect 200684 52714 200712 74506
rect 203524 62960 203576 62966
rect 203524 62902 203576 62908
rect 203536 54534 203564 62902
rect 204272 54534 204300 77302
rect 204350 73808 204406 73817
rect 204350 73743 204406 73752
rect 203524 54528 203576 54534
rect 202878 54496 202934 54505
rect 203524 54470 203576 54476
rect 204260 54528 204312 54534
rect 204260 54470 204312 54476
rect 202878 54431 202934 54440
rect 198844 52686 199226 52714
rect 200684 52686 201066 52714
rect 202892 52700 202920 54431
rect 204364 52714 204392 73743
rect 209792 65550 209820 77302
rect 216048 75818 216076 77302
rect 219544 77302 220800 77330
rect 225860 77302 226196 77330
rect 230920 77302 231256 77330
rect 219440 76084 219492 76090
rect 219440 76026 219492 76032
rect 216036 75812 216088 75818
rect 216036 75754 216088 75760
rect 217324 75812 217376 75818
rect 217324 75754 217376 75760
rect 211712 72684 211764 72690
rect 211712 72626 211764 72632
rect 209780 65544 209832 65550
rect 209780 65486 209832 65492
rect 206284 64320 206336 64326
rect 206284 64262 206336 64268
rect 206296 54602 206324 64262
rect 208400 54664 208452 54670
rect 208400 54606 208452 54612
rect 206284 54596 206336 54602
rect 206284 54538 206336 54544
rect 206560 54460 206612 54466
rect 206560 54402 206612 54408
rect 204364 52686 204746 52714
rect 206572 52700 206600 54402
rect 208412 52700 208440 54606
rect 210240 54528 210292 54534
rect 210240 54470 210292 54476
rect 210252 52700 210280 54470
rect 211724 52714 211752 72626
rect 217336 67590 217364 75754
rect 217324 67584 217376 67590
rect 217324 67526 217376 67532
rect 217230 59936 217286 59945
rect 217230 59871 217286 59880
rect 215758 57488 215814 57497
rect 215758 57423 215814 57432
rect 213918 57352 213974 57361
rect 213918 57287 213974 57296
rect 211724 52686 212106 52714
rect 213932 52700 213960 57287
rect 215772 52700 215800 57423
rect 217244 52714 217272 59871
rect 217244 52686 217626 52714
rect 219452 52700 219480 76026
rect 219544 65686 219572 77302
rect 224958 76664 225014 76673
rect 222200 76628 222252 76634
rect 224958 76599 225014 76608
rect 222200 76570 222252 76576
rect 222212 74534 222240 76570
rect 222212 74506 222792 74534
rect 219532 65680 219584 65686
rect 219532 65622 219584 65628
rect 221280 53848 221332 53854
rect 221280 53790 221332 53796
rect 221292 52700 221320 53790
rect 222764 52714 222792 74506
rect 222764 52686 223146 52714
rect 224972 52700 225000 76599
rect 226168 75206 226196 77302
rect 226156 75200 226208 75206
rect 226156 75142 226208 75148
rect 231228 75138 231256 77302
rect 235920 77302 235980 77330
rect 235920 75342 235948 77302
rect 235908 75336 235960 75342
rect 235908 75278 235960 75284
rect 240048 75336 240100 75342
rect 240048 75278 240100 75284
rect 234436 75200 234488 75206
rect 233238 75168 233294 75177
rect 231216 75132 231268 75138
rect 234436 75142 234488 75148
rect 239496 75200 239548 75206
rect 239496 75142 239548 75148
rect 233238 75103 233294 75112
rect 231216 75074 231268 75080
rect 233252 74534 233280 75103
rect 233252 74506 233832 74534
rect 226432 73840 226484 73846
rect 226432 73782 226484 73788
rect 226444 52714 226472 73782
rect 231952 67040 232004 67046
rect 231952 66982 232004 66988
rect 228272 65612 228324 65618
rect 228272 65554 228324 65560
rect 226984 65544 227036 65550
rect 226984 65486 227036 65492
rect 226996 55214 227024 65486
rect 226984 55208 227036 55214
rect 226984 55150 227036 55156
rect 228284 52714 228312 65554
rect 230480 65544 230532 65550
rect 230480 65486 230532 65492
rect 226444 52686 226826 52714
rect 228284 52686 228666 52714
rect 230492 52700 230520 65486
rect 231964 52714 231992 66982
rect 233804 52714 233832 74506
rect 234448 68338 234476 75142
rect 235908 75132 235960 75138
rect 235908 75074 235960 75080
rect 234436 68332 234488 68338
rect 234436 68274 234488 68280
rect 235920 56030 235948 75074
rect 239404 71324 239456 71330
rect 239404 71266 239456 71272
rect 237472 69964 237524 69970
rect 237472 69906 237524 69912
rect 235908 56024 235960 56030
rect 235908 55966 235960 55972
rect 236000 54596 236052 54602
rect 236000 54538 236052 54544
rect 231964 52686 232346 52714
rect 233804 52686 234186 52714
rect 236012 52700 236040 54538
rect 237484 52714 237512 69906
rect 239416 55214 239444 71266
rect 239508 69970 239536 75142
rect 239496 69964 239548 69970
rect 239496 69906 239548 69912
rect 239404 55208 239456 55214
rect 239404 55150 239456 55156
rect 239416 52714 239444 55150
rect 240060 54738 240088 75278
rect 240796 67590 240824 77862
rect 284298 77752 284354 77761
rect 284298 77687 284354 77696
rect 241040 77302 241376 77330
rect 246100 77302 246436 77330
rect 241348 75478 241376 77302
rect 241336 75472 241388 75478
rect 241336 75414 241388 75420
rect 246408 75410 246436 77302
rect 251100 77302 251160 77330
rect 256220 77302 256648 77330
rect 261280 77302 261616 77330
rect 251100 75478 251128 77302
rect 248420 75472 248472 75478
rect 248420 75414 248472 75420
rect 251088 75472 251140 75478
rect 251088 75414 251140 75420
rect 246396 75404 246448 75410
rect 246396 75346 246448 75352
rect 248432 71262 248460 75414
rect 256620 74526 256648 77302
rect 261588 75818 261616 77302
rect 266280 77302 266340 77330
rect 271400 77302 271736 77330
rect 261576 75812 261628 75818
rect 261576 75754 261628 75760
rect 264888 75812 264940 75818
rect 264888 75754 264940 75760
rect 261484 75472 261536 75478
rect 261484 75414 261536 75420
rect 256608 74520 256660 74526
rect 256608 74462 256660 74468
rect 254032 72548 254084 72554
rect 254032 72490 254084 72496
rect 248420 71256 248472 71262
rect 248420 71198 248472 71204
rect 252560 69692 252612 69698
rect 252560 69634 252612 69640
rect 244832 68332 244884 68338
rect 244832 68274 244884 68280
rect 244844 67590 244872 68274
rect 240784 67584 240836 67590
rect 240784 67526 240836 67532
rect 244832 67584 244884 67590
rect 244832 67526 244884 67532
rect 240048 54732 240100 54738
rect 240048 54674 240100 54680
rect 240796 53922 240824 67526
rect 242992 65680 243044 65686
rect 242992 65622 243044 65628
rect 243004 65006 243032 65622
rect 242992 65000 243044 65006
rect 242992 64942 243044 64948
rect 243820 65000 243872 65006
rect 243820 64942 243872 64948
rect 240784 53916 240836 53922
rect 240784 53858 240836 53864
rect 241520 53916 241572 53922
rect 241520 53858 241572 53864
rect 237484 52686 237866 52714
rect 239416 52686 239706 52714
rect 241532 52700 241560 53858
rect 243004 52714 243032 64942
rect 243832 64870 243860 64942
rect 243820 64864 243872 64870
rect 243820 64806 243872 64812
rect 244844 52714 244872 67526
rect 247040 56024 247092 56030
rect 247040 55966 247092 55972
rect 243004 52686 243386 52714
rect 244844 52686 245226 52714
rect 247052 52700 247080 55966
rect 248880 54732 248932 54738
rect 248880 54674 248932 54680
rect 250720 54732 250772 54738
rect 250720 54674 250772 54680
rect 248892 52700 248920 54674
rect 250732 52700 250760 54674
rect 252572 52700 252600 69634
rect 254044 52714 254072 72490
rect 255872 66904 255924 66910
rect 255872 66846 255924 66852
rect 255884 52714 255912 66846
rect 256620 56030 256648 74462
rect 261392 71256 261444 71262
rect 261392 71198 261444 71204
rect 258080 68332 258132 68338
rect 258080 68274 258132 68280
rect 256608 56024 256660 56030
rect 256608 55966 256660 55972
rect 254044 52686 254426 52714
rect 255884 52686 256266 52714
rect 258092 52700 258120 68274
rect 259920 57248 259972 57254
rect 259920 57190 259972 57196
rect 259932 52700 259960 57190
rect 261404 52714 261432 71198
rect 261496 67522 261524 75414
rect 263600 75404 263652 75410
rect 263600 75346 263652 75352
rect 262128 71392 262180 71398
rect 262128 71334 262180 71340
rect 262140 71262 262168 71334
rect 262128 71256 262180 71262
rect 262128 71198 262180 71204
rect 261484 67516 261536 67522
rect 261484 67458 261536 67464
rect 261404 52686 261786 52714
rect 263612 52700 263640 75346
rect 264900 69902 264928 75754
rect 266280 75546 266308 77302
rect 266268 75540 266320 75546
rect 266268 75482 266320 75488
rect 270500 75540 270552 75546
rect 270500 75482 270552 75488
rect 270512 74594 270540 75482
rect 271708 74866 271736 77302
rect 276032 77302 276460 77330
rect 281460 77302 281520 77330
rect 271696 74860 271748 74866
rect 271696 74802 271748 74808
rect 270500 74588 270552 74594
rect 270500 74530 270552 74536
rect 271788 74588 271840 74594
rect 271788 74530 271840 74536
rect 264888 69896 264940 69902
rect 264888 69838 264940 69844
rect 269120 69896 269172 69902
rect 269120 69838 269172 69844
rect 265624 68468 265676 68474
rect 265624 68410 265676 68416
rect 265072 67516 265124 67522
rect 265072 67458 265124 67464
rect 265084 67114 265112 67458
rect 265072 67108 265124 67114
rect 265072 67050 265124 67056
rect 265084 52714 265112 67050
rect 265636 54738 265664 68410
rect 267280 56024 267332 56030
rect 267280 55966 267332 55972
rect 265624 54732 265676 54738
rect 265624 54674 265676 54680
rect 265084 52686 265466 52714
rect 267292 52700 267320 55966
rect 269132 52700 269160 69838
rect 270512 64874 270540 74530
rect 271800 74458 271828 74530
rect 271788 74452 271840 74458
rect 271788 74394 271840 74400
rect 272432 68536 272484 68542
rect 272432 68478 272484 68484
rect 271144 65680 271196 65686
rect 271144 65622 271196 65628
rect 270512 64846 270632 64874
rect 270604 52714 270632 64846
rect 271156 54670 271184 65622
rect 271144 54664 271196 54670
rect 271144 54606 271196 54612
rect 272444 52714 272472 68478
rect 274640 54732 274692 54738
rect 274640 54674 274692 54680
rect 270604 52686 270986 52714
rect 272444 52686 272826 52714
rect 274652 52700 274680 54674
rect 276032 54670 276060 77302
rect 276112 74860 276164 74866
rect 276112 74802 276164 74808
rect 276124 68542 276152 74802
rect 281460 74390 281488 77302
rect 282182 76800 282238 76809
rect 282182 76735 282238 76744
rect 281448 74384 281500 74390
rect 281448 74326 281500 74332
rect 276112 68536 276164 68542
rect 276112 68478 276164 68484
rect 281460 56030 281488 74326
rect 281448 56024 281500 56030
rect 281448 55966 281500 55972
rect 278320 54868 278372 54874
rect 278320 54810 278372 54816
rect 276020 54664 276072 54670
rect 276020 54606 276072 54612
rect 276478 54632 276534 54641
rect 276478 54567 276534 54576
rect 276492 52700 276520 54567
rect 278332 52700 278360 54810
rect 282000 54800 282052 54806
rect 280158 54768 280214 54777
rect 282000 54742 282052 54748
rect 280158 54703 280214 54712
rect 280172 52700 280200 54703
rect 282012 52700 282040 54742
rect 282196 54505 282224 76735
rect 284312 75886 284340 77687
rect 284300 75880 284352 75886
rect 284300 75822 284352 75828
rect 282274 73944 282330 73953
rect 282274 73879 282330 73888
rect 282288 54534 282316 73879
rect 284956 68610 284984 77862
rect 286580 77302 286824 77330
rect 286796 75478 286824 77302
rect 286784 75472 286836 75478
rect 286784 75414 286836 75420
rect 284944 68604 284996 68610
rect 284944 68546 284996 68552
rect 282276 54528 282328 54534
rect 282182 54496 282238 54505
rect 282276 54470 282328 54476
rect 283838 54496 283894 54505
rect 282182 54431 282238 54440
rect 283838 54431 283894 54440
rect 283852 52700 283880 54431
rect 285680 54324 285732 54330
rect 285680 54266 285732 54272
rect 285692 52700 285720 54266
rect 285770 53952 285826 53961
rect 285770 53887 285826 53896
rect 285784 53854 285812 53887
rect 285772 53848 285824 53854
rect 285772 53790 285824 53796
rect 287532 52700 287560 189722
rect 287808 67590 287836 190426
rect 287900 75342 287928 204410
rect 287888 75336 287940 75342
rect 287888 75278 287940 75284
rect 287796 67584 287848 67590
rect 287796 67526 287848 67532
rect 287610 54904 287666 54913
rect 288452 54874 288480 458798
rect 288544 315926 288572 458934
rect 288820 458114 288848 583170
rect 288808 458108 288860 458114
rect 288808 458050 288860 458056
rect 289832 458046 289860 585822
rect 289820 458040 289872 458046
rect 289820 457982 289872 457988
rect 289084 457564 289136 457570
rect 289084 457506 289136 457512
rect 288624 441924 288676 441930
rect 288624 441866 288676 441872
rect 288636 334257 288664 441866
rect 288622 334248 288678 334257
rect 288622 334183 288678 334192
rect 289096 331906 289124 457506
rect 289832 451274 289860 457982
rect 289924 457570 289952 585958
rect 290016 459406 290044 586026
rect 301872 586016 301924 586022
rect 301872 585958 301924 585964
rect 300676 583364 300728 583370
rect 300676 583306 300728 583312
rect 292580 583296 292632 583302
rect 292580 583238 292632 583244
rect 300492 583296 300544 583302
rect 300492 583238 300544 583244
rect 291476 583160 291528 583166
rect 291476 583102 291528 583108
rect 291200 583092 291252 583098
rect 291200 583034 291252 583040
rect 290096 572076 290148 572082
rect 290096 572018 290148 572024
rect 290108 480254 290136 572018
rect 290108 480226 290228 480254
rect 290200 460834 290228 480226
rect 290188 460828 290240 460834
rect 290188 460770 290240 460776
rect 290004 459400 290056 459406
rect 290004 459342 290056 459348
rect 290016 458250 290044 459342
rect 290004 458244 290056 458250
rect 290004 458186 290056 458192
rect 289912 457564 289964 457570
rect 289912 457506 289964 457512
rect 289832 451246 290044 451274
rect 290016 335354 290044 451246
rect 290094 433936 290150 433945
rect 290094 433871 290150 433880
rect 289832 335326 290044 335354
rect 289832 332518 289860 335326
rect 290108 334121 290136 433871
rect 290094 334112 290150 334121
rect 290094 334047 290150 334056
rect 290200 332586 290228 460770
rect 291212 458998 291240 583034
rect 291382 459776 291438 459785
rect 291382 459711 291438 459720
rect 291200 458992 291252 458998
rect 291200 458934 291252 458940
rect 290280 458244 290332 458250
rect 290280 458186 290332 458192
rect 290188 332580 290240 332586
rect 290188 332522 290240 332528
rect 289820 332512 289872 332518
rect 289820 332454 289872 332460
rect 289910 332480 289966 332489
rect 289084 331900 289136 331906
rect 289084 331842 289136 331848
rect 289084 319456 289136 319462
rect 289084 319398 289136 319404
rect 288532 315920 288584 315926
rect 288532 315862 288584 315868
rect 288544 201414 288572 315862
rect 288624 313948 288676 313954
rect 288624 313890 288676 313896
rect 288636 205970 288664 313890
rect 288624 205964 288676 205970
rect 288624 205906 288676 205912
rect 288532 201408 288584 201414
rect 288532 201350 288584 201356
rect 288544 78062 288572 201350
rect 288622 177984 288678 177993
rect 288622 177919 288678 177928
rect 288532 78056 288584 78062
rect 288532 77998 288584 78004
rect 288636 72690 288664 177919
rect 288624 72684 288676 72690
rect 288624 72626 288676 72632
rect 288992 71256 289044 71262
rect 288992 71198 289044 71204
rect 287610 54839 287666 54848
rect 288440 54868 288492 54874
rect 287624 54806 287652 54839
rect 288440 54810 288492 54816
rect 287612 54800 287664 54806
rect 287612 54742 287664 54748
rect 289004 52714 289032 71198
rect 289096 54330 289124 319398
rect 289832 204134 289860 332454
rect 289910 332415 289966 332424
rect 289924 204542 289952 332415
rect 290096 315444 290148 315450
rect 290096 315386 290148 315392
rect 289912 204536 289964 204542
rect 289912 204478 289964 204484
rect 289820 204128 289872 204134
rect 289820 204070 289872 204076
rect 289820 203584 289872 203590
rect 289820 203526 289872 203532
rect 289832 54738 289860 203526
rect 289924 71398 289952 204478
rect 290108 204338 290136 315386
rect 290200 204610 290228 332522
rect 290292 332314 290320 458186
rect 291292 458108 291344 458114
rect 291292 458050 291344 458056
rect 291200 457496 291252 457502
rect 291200 457438 291252 457444
rect 290280 332308 290332 332314
rect 290280 332250 290332 332256
rect 290292 331294 290320 332250
rect 290280 331288 290332 331294
rect 290280 331230 290332 331236
rect 291212 315790 291240 457438
rect 291304 332722 291332 458050
rect 291292 332716 291344 332722
rect 291292 332658 291344 332664
rect 291304 331106 291332 332658
rect 291396 331226 291424 459711
rect 291488 444378 291516 583102
rect 291844 580440 291896 580446
rect 291844 580382 291896 580388
rect 291856 460222 291884 580382
rect 291844 460216 291896 460222
rect 291844 460158 291896 460164
rect 291856 459610 291884 460158
rect 291844 459604 291896 459610
rect 291844 459546 291896 459552
rect 292592 457502 292620 583238
rect 299296 583160 299348 583166
rect 299296 583102 299348 583108
rect 293224 583024 293276 583030
rect 293224 582966 293276 582972
rect 298006 582992 298062 583001
rect 292672 577516 292724 577522
rect 292672 577458 292724 577464
rect 292684 461650 292712 577458
rect 292672 461644 292724 461650
rect 292672 461586 292724 461592
rect 292764 458924 292816 458930
rect 292764 458866 292816 458872
rect 292580 457496 292632 457502
rect 292580 457438 292632 457444
rect 291476 444372 291528 444378
rect 291476 444314 291528 444320
rect 291488 443970 291516 444314
rect 291476 443964 291528 443970
rect 291476 443906 291528 443912
rect 292776 333334 292804 458866
rect 292856 443964 292908 443970
rect 292856 443906 292908 443912
rect 292764 333328 292816 333334
rect 292764 333270 292816 333276
rect 292580 331900 292632 331906
rect 292580 331842 292632 331848
rect 291384 331220 291436 331226
rect 291384 331162 291436 331168
rect 291304 331078 291516 331106
rect 291384 330540 291436 330546
rect 291384 330482 291436 330488
rect 291200 315784 291252 315790
rect 291200 315726 291252 315732
rect 290188 204604 290240 204610
rect 290188 204546 290240 204552
rect 291212 204474 291240 315726
rect 291396 204950 291424 330482
rect 291488 325694 291516 331078
rect 291488 325666 291608 325694
rect 291474 305688 291530 305697
rect 291474 305623 291530 305632
rect 291488 206009 291516 305623
rect 291474 206000 291530 206009
rect 291474 205935 291530 205944
rect 291384 204944 291436 204950
rect 291384 204886 291436 204892
rect 291200 204468 291252 204474
rect 291200 204410 291252 204416
rect 290096 204332 290148 204338
rect 290096 204274 290148 204280
rect 291200 204264 291252 204270
rect 291200 204206 291252 204212
rect 290002 203688 290058 203697
rect 291212 203658 291240 204206
rect 291384 204196 291436 204202
rect 291384 204138 291436 204144
rect 291292 203924 291344 203930
rect 291292 203866 291344 203872
rect 290002 203623 290058 203632
rect 291200 203652 291252 203658
rect 290016 74526 290044 203623
rect 291200 203594 291252 203600
rect 290096 185904 290148 185910
rect 290096 185846 290148 185852
rect 290108 77994 290136 185846
rect 290096 77988 290148 77994
rect 290096 77930 290148 77936
rect 290004 74520 290056 74526
rect 290004 74462 290056 74468
rect 289912 71392 289964 71398
rect 289912 71334 289964 71340
rect 291212 69902 291240 203594
rect 291304 74390 291332 203866
rect 291396 203726 291424 204138
rect 291384 203720 291436 203726
rect 291384 203662 291436 203668
rect 291396 74458 291424 203662
rect 291580 201278 291608 325666
rect 292592 204270 292620 331842
rect 292672 331288 292724 331294
rect 292672 331230 292724 331236
rect 292580 204264 292632 204270
rect 292580 204206 292632 204212
rect 292684 204202 292712 331230
rect 292868 331090 292896 443906
rect 293236 331945 293264 582966
rect 298006 582927 298062 582936
rect 295340 580576 295392 580582
rect 295340 580518 295392 580524
rect 295156 580440 295208 580446
rect 295156 580382 295208 580388
rect 294604 572144 294656 572150
rect 294604 572086 294656 572092
rect 293960 459604 294012 459610
rect 293960 459546 294012 459552
rect 293222 331936 293278 331945
rect 293222 331871 293278 331880
rect 293868 331220 293920 331226
rect 293868 331162 293920 331168
rect 292856 331084 292908 331090
rect 292856 331026 292908 331032
rect 292868 330750 292896 331026
rect 292856 330744 292908 330750
rect 292856 330686 292908 330692
rect 292764 314084 292816 314090
rect 292764 314026 292816 314032
rect 292672 204196 292724 204202
rect 292672 204138 292724 204144
rect 292776 201482 292804 314026
rect 293880 204950 293908 331162
rect 293972 330546 294000 459546
rect 294144 330744 294196 330750
rect 294144 330686 294196 330692
rect 293960 330540 294012 330546
rect 293960 330482 294012 330488
rect 294052 329792 294104 329798
rect 294052 329734 294104 329740
rect 294064 329118 294092 329734
rect 294052 329112 294104 329118
rect 294052 329054 294104 329060
rect 294064 205737 294092 329054
rect 294050 205728 294106 205737
rect 294050 205663 294106 205672
rect 293868 204944 293920 204950
rect 293868 204886 293920 204892
rect 294156 204762 294184 330686
rect 293972 204734 294184 204762
rect 292856 204604 292908 204610
rect 292856 204546 292908 204552
rect 292764 201476 292816 201482
rect 292764 201418 292816 201424
rect 291568 201272 291620 201278
rect 291568 201214 291620 201220
rect 292672 201272 292724 201278
rect 292672 201214 292724 201220
rect 291474 185872 291530 185881
rect 291474 185807 291530 185816
rect 291488 77761 291516 185807
rect 291474 77752 291530 77761
rect 291474 77687 291530 77696
rect 291474 76392 291530 76401
rect 291474 76327 291530 76336
rect 291488 76022 291516 76327
rect 291476 76016 291528 76022
rect 291476 75958 291528 75964
rect 292684 75274 292712 201214
rect 292764 185972 292816 185978
rect 292764 185914 292816 185920
rect 292672 75268 292724 75274
rect 292672 75210 292724 75216
rect 291384 74452 291436 74458
rect 291384 74394 291436 74400
rect 291292 74384 291344 74390
rect 291292 74326 291344 74332
rect 292776 71330 292804 185914
rect 292868 75410 292896 204546
rect 293972 204406 294000 204734
rect 293960 204400 294012 204406
rect 293960 204342 294012 204348
rect 293224 203788 293276 203794
rect 293224 203730 293276 203736
rect 293236 76702 293264 203730
rect 293224 76696 293276 76702
rect 293224 76638 293276 76644
rect 292856 75404 292908 75410
rect 292856 75346 292908 75352
rect 292856 75268 292908 75274
rect 292856 75210 292908 75216
rect 292764 71324 292816 71330
rect 292764 71266 292816 71272
rect 291200 69896 291252 69902
rect 291200 69838 291252 69844
rect 289820 54732 289872 54738
rect 289820 54674 289872 54680
rect 291200 54732 291252 54738
rect 291200 54674 291252 54680
rect 289084 54324 289136 54330
rect 289084 54266 289136 54272
rect 289004 52686 289386 52714
rect 291212 52700 291240 54674
rect 292868 52714 292896 75210
rect 293972 64870 294000 204342
rect 294052 204128 294104 204134
rect 294052 204070 294104 204076
rect 294064 67114 294092 204070
rect 294144 187060 294196 187066
rect 294144 187002 294196 187008
rect 294156 77926 294184 187002
rect 294144 77920 294196 77926
rect 294144 77862 294196 77868
rect 294052 67108 294104 67114
rect 294052 67050 294104 67056
rect 293960 64864 294012 64870
rect 293960 64806 294012 64812
rect 294616 57526 294644 572086
rect 295168 460902 295196 580382
rect 295248 577516 295300 577522
rect 295248 577458 295300 577464
rect 295156 460896 295208 460902
rect 295156 460838 295208 460844
rect 295260 455394 295288 577458
rect 295352 459542 295380 580518
rect 295432 580372 295484 580378
rect 295432 580314 295484 580320
rect 297824 580372 297876 580378
rect 297824 580314 297876 580320
rect 295340 459536 295392 459542
rect 295340 459478 295392 459484
rect 295248 455388 295300 455394
rect 295248 455330 295300 455336
rect 295260 333334 295288 455330
rect 295248 333328 295300 333334
rect 295248 333270 295300 333276
rect 295352 329798 295380 459478
rect 295444 458930 295472 580314
rect 295524 580304 295576 580310
rect 295524 580246 295576 580252
rect 295536 460290 295564 580246
rect 296536 461644 296588 461650
rect 296536 461586 296588 461592
rect 295524 460284 295576 460290
rect 295524 460226 295576 460232
rect 295432 458924 295484 458930
rect 295432 458866 295484 458872
rect 296548 329798 296576 461586
rect 296720 460964 296772 460970
rect 296720 460906 296772 460912
rect 296628 460896 296680 460902
rect 296628 460838 296680 460844
rect 296640 332722 296668 460838
rect 296628 332716 296680 332722
rect 296628 332658 296680 332664
rect 295340 329792 295392 329798
rect 295340 329734 295392 329740
rect 296536 329792 296588 329798
rect 296536 329734 296588 329740
rect 296536 315920 296588 315926
rect 296536 315862 296588 315868
rect 295984 315376 296036 315382
rect 295984 315318 296036 315324
rect 295338 186008 295394 186017
rect 295338 185943 295394 185952
rect 295352 77897 295380 185943
rect 295338 77888 295394 77897
rect 295338 77823 295394 77832
rect 295996 60246 296024 315318
rect 296444 313948 296496 313954
rect 296444 313890 296496 313896
rect 296456 206310 296484 313890
rect 296444 206304 296496 206310
rect 296444 206246 296496 206252
rect 296444 201408 296496 201414
rect 296444 201350 296496 201356
rect 295984 60240 296036 60246
rect 295984 60182 296036 60188
rect 294604 57520 294656 57526
rect 294604 57462 294656 57468
rect 294880 56160 294932 56166
rect 294880 56102 294932 56108
rect 294604 56024 294656 56030
rect 294604 55966 294656 55972
rect 294616 54534 294644 55966
rect 294604 54528 294656 54534
rect 294604 54470 294656 54476
rect 292868 52686 293066 52714
rect 294892 52700 294920 56102
rect 296456 54874 296484 201350
rect 296548 188358 296576 315862
rect 296640 200802 296668 332658
rect 296732 331226 296760 460906
rect 297836 460902 297864 580314
rect 297916 577584 297968 577590
rect 297916 577526 297968 577532
rect 297824 460896 297876 460902
rect 297824 460838 297876 460844
rect 297180 444304 297232 444310
rect 297180 444246 297232 444252
rect 297192 444009 297220 444246
rect 297178 444000 297234 444009
rect 297178 443935 297234 443944
rect 297928 442921 297956 577526
rect 298020 458182 298048 582927
rect 299204 580576 299256 580582
rect 299204 580518 299256 580524
rect 299112 577652 299164 577658
rect 299112 577594 299164 577600
rect 298928 459604 298980 459610
rect 298928 459546 298980 459552
rect 298008 458176 298060 458182
rect 298008 458118 298060 458124
rect 297914 442912 297970 442921
rect 297914 442847 297970 442856
rect 296812 442264 296864 442270
rect 296812 442206 296864 442212
rect 296824 333266 296852 442206
rect 296812 333260 296864 333266
rect 296812 333202 296864 333208
rect 296720 331220 296772 331226
rect 296720 331162 296772 331168
rect 297732 329792 297784 329798
rect 297732 329734 297784 329740
rect 297744 329118 297772 329734
rect 297732 329112 297784 329118
rect 297732 329054 297784 329060
rect 297916 329112 297968 329118
rect 297916 329054 297968 329060
rect 297364 315308 297416 315314
rect 297364 315250 297416 315256
rect 296720 314016 296772 314022
rect 296720 313958 296772 313964
rect 296732 202842 296760 313958
rect 296720 202836 296772 202842
rect 296720 202778 296772 202784
rect 296628 200796 296680 200802
rect 296628 200738 296680 200744
rect 296536 188352 296588 188358
rect 296536 188294 296588 188300
rect 296536 187196 296588 187202
rect 296536 187138 296588 187144
rect 296548 70378 296576 187138
rect 297178 76936 297234 76945
rect 297178 76871 297234 76880
rect 297192 76090 297220 76871
rect 297180 76084 297232 76090
rect 297180 76026 297232 76032
rect 296536 70372 296588 70378
rect 296536 70314 296588 70320
rect 296444 54868 296496 54874
rect 296444 54810 296496 54816
rect 297376 54806 297404 315250
rect 297824 314696 297876 314702
rect 297824 314638 297876 314644
rect 297836 204882 297864 314638
rect 297928 205057 297956 329054
rect 298020 315926 298048 458118
rect 298008 315920 298060 315926
rect 298008 315862 298060 315868
rect 298940 315790 298968 459546
rect 299124 456754 299152 577594
rect 299216 459406 299244 580518
rect 299204 459400 299256 459406
rect 299204 459342 299256 459348
rect 299112 456748 299164 456754
rect 299112 456690 299164 456696
rect 299124 332790 299152 456690
rect 299112 332784 299164 332790
rect 299112 332726 299164 332732
rect 299020 331356 299072 331362
rect 299020 331298 299072 331304
rect 298928 315784 298980 315790
rect 298928 315726 298980 315732
rect 298940 314702 298968 315726
rect 298928 314696 298980 314702
rect 298928 314638 298980 314644
rect 297914 205048 297970 205057
rect 297914 204983 297970 204992
rect 297824 204876 297876 204882
rect 297824 204818 297876 204824
rect 298008 204808 298060 204814
rect 298008 204750 298060 204756
rect 297824 187604 297876 187610
rect 297824 187546 297876 187552
rect 297836 77994 297864 187546
rect 297916 186448 297968 186454
rect 297916 186390 297968 186396
rect 297824 77988 297876 77994
rect 297824 77930 297876 77936
rect 297928 63102 297956 186390
rect 297916 63096 297968 63102
rect 297916 63038 297968 63044
rect 297456 60376 297508 60382
rect 297456 60318 297508 60324
rect 297364 54800 297416 54806
rect 297364 54742 297416 54748
rect 297468 54738 297496 60318
rect 298020 56030 298048 204750
rect 299032 204270 299060 331298
rect 299216 330290 299244 459342
rect 299308 459338 299336 583102
rect 299388 580304 299440 580310
rect 299388 580246 299440 580252
rect 299400 461650 299428 580246
rect 300504 470594 300532 583238
rect 300584 583092 300636 583098
rect 300584 583034 300636 583040
rect 300412 470566 300532 470594
rect 299388 461644 299440 461650
rect 299388 461586 299440 461592
rect 300412 460086 300440 470566
rect 300596 460834 300624 583034
rect 300584 460828 300636 460834
rect 300584 460770 300636 460776
rect 300400 460080 300452 460086
rect 300400 460022 300452 460028
rect 300596 459610 300624 460770
rect 300584 459604 300636 459610
rect 300584 459546 300636 459552
rect 299296 459332 299348 459338
rect 299296 459274 299348 459280
rect 299124 330262 299244 330290
rect 299124 329769 299152 330262
rect 299204 329792 299256 329798
rect 299110 329760 299166 329769
rect 299204 329734 299256 329740
rect 299110 329695 299166 329704
rect 299124 329594 299152 329695
rect 299112 329588 299164 329594
rect 299112 329530 299164 329536
rect 299112 314696 299164 314702
rect 299112 314638 299164 314644
rect 299020 204264 299072 204270
rect 299020 204206 299072 204212
rect 299124 186998 299152 314638
rect 299216 201414 299244 329734
rect 299308 325694 299336 459274
rect 300490 458280 300546 458289
rect 300490 458215 300546 458224
rect 300400 457632 300452 457638
rect 300400 457574 300452 457580
rect 300308 443556 300360 443562
rect 300308 443498 300360 443504
rect 300122 331800 300178 331809
rect 300122 331735 300178 331744
rect 299308 325666 299428 325694
rect 299400 315722 299428 325666
rect 299388 315716 299440 315722
rect 299388 315658 299440 315664
rect 299400 204814 299428 315658
rect 299388 204808 299440 204814
rect 299388 204750 299440 204756
rect 299400 204610 299428 204750
rect 299388 204604 299440 204610
rect 299388 204546 299440 204552
rect 299296 204264 299348 204270
rect 299296 204206 299348 204212
rect 299388 204264 299440 204270
rect 299388 204206 299440 204212
rect 299308 204134 299336 204206
rect 299296 204128 299348 204134
rect 299296 204070 299348 204076
rect 299204 201408 299256 201414
rect 299204 201350 299256 201356
rect 299202 201240 299258 201249
rect 299202 201175 299258 201184
rect 299216 200870 299244 201175
rect 299204 200864 299256 200870
rect 299204 200806 299256 200812
rect 298744 186992 298796 186998
rect 298744 186934 298796 186940
rect 299112 186992 299164 186998
rect 299112 186934 299164 186940
rect 298756 60314 298784 186934
rect 299216 76770 299244 200806
rect 299204 76764 299256 76770
rect 299204 76706 299256 76712
rect 299308 62082 299336 204070
rect 299296 62076 299348 62082
rect 299296 62018 299348 62024
rect 299308 60790 299336 62018
rect 298836 60784 298888 60790
rect 298836 60726 298888 60732
rect 299296 60784 299348 60790
rect 299296 60726 299348 60732
rect 298744 60308 298796 60314
rect 298744 60250 298796 60256
rect 298560 56228 298612 56234
rect 298560 56170 298612 56176
rect 298008 56024 298060 56030
rect 298008 55966 298060 55972
rect 297456 54732 297508 54738
rect 297456 54674 297508 54680
rect 296720 53848 296772 53854
rect 296720 53790 296772 53796
rect 296732 52700 296760 53790
rect 298572 52700 298600 56170
rect 298848 53854 298876 60726
rect 299400 56574 299428 204206
rect 300136 76634 300164 331735
rect 300320 315654 300348 443498
rect 300412 332178 300440 457574
rect 300504 333674 300532 458215
rect 300688 458114 300716 583306
rect 300768 583228 300820 583234
rect 300768 583170 300820 583176
rect 300676 458108 300728 458114
rect 300676 458050 300728 458056
rect 300688 345014 300716 458050
rect 300780 444378 300808 583170
rect 301780 460080 301832 460086
rect 301780 460022 301832 460028
rect 300768 444372 300820 444378
rect 300768 444314 300820 444320
rect 300780 443562 300808 444314
rect 300768 443556 300820 443562
rect 300768 443498 300820 443504
rect 300688 344986 300808 345014
rect 300492 333668 300544 333674
rect 300492 333610 300544 333616
rect 300400 332172 300452 332178
rect 300400 332114 300452 332120
rect 300412 325694 300440 332114
rect 300780 329798 300808 344986
rect 301792 329798 301820 460022
rect 301884 459950 301912 585958
rect 301964 583024 302016 583030
rect 301964 582966 302016 582972
rect 301872 459944 301924 459950
rect 301872 459886 301924 459892
rect 301870 459504 301926 459513
rect 301870 459439 301872 459448
rect 301924 459439 301926 459448
rect 301872 459410 301924 459416
rect 301976 457502 302004 582966
rect 302068 459542 302096 586026
rect 318628 586022 318656 587316
rect 318616 586016 318668 586022
rect 318616 585958 318668 585964
rect 323688 585954 323716 587316
rect 303160 585948 303212 585954
rect 303160 585890 303212 585896
rect 323676 585948 323728 585954
rect 323676 585890 323728 585896
rect 302148 585880 302200 585886
rect 302148 585822 302200 585828
rect 302056 459536 302108 459542
rect 302056 459478 302108 459484
rect 301964 457496 302016 457502
rect 301964 457438 302016 457444
rect 301872 456680 301924 456686
rect 301872 456622 301924 456628
rect 301884 332586 301912 456622
rect 301872 332580 301924 332586
rect 301872 332522 301924 332528
rect 302068 332314 302096 459478
rect 302160 457978 302188 585822
rect 302976 580508 303028 580514
rect 302976 580450 303028 580456
rect 302148 457972 302200 457978
rect 302148 457914 302200 457920
rect 302160 332450 302188 457914
rect 302988 456686 303016 580450
rect 303068 459944 303120 459950
rect 303068 459886 303120 459892
rect 303080 459270 303108 459886
rect 303068 459264 303120 459270
rect 303068 459206 303120 459212
rect 302976 456680 303028 456686
rect 302976 456622 303028 456628
rect 303080 332518 303108 459206
rect 303172 459105 303200 585890
rect 328748 585886 328776 587316
rect 328736 585880 328788 585886
rect 328736 585822 328788 585828
rect 333808 585818 333836 587316
rect 303252 585812 303304 585818
rect 303252 585754 303304 585760
rect 333796 585812 333848 585818
rect 333796 585754 333848 585760
rect 303158 459096 303214 459105
rect 303158 459031 303214 459040
rect 303068 332512 303120 332518
rect 303068 332454 303120 332460
rect 302148 332444 302200 332450
rect 302148 332386 302200 332392
rect 302056 332308 302108 332314
rect 302056 332250 302108 332256
rect 301964 331288 302016 331294
rect 301964 331230 302016 331236
rect 300768 329792 300820 329798
rect 300768 329734 300820 329740
rect 301780 329792 301832 329798
rect 301780 329734 301832 329740
rect 300412 325666 300808 325694
rect 300584 316056 300636 316062
rect 300584 315998 300636 316004
rect 300308 315648 300360 315654
rect 300308 315590 300360 315596
rect 300320 314702 300348 315590
rect 300308 314696 300360 314702
rect 300308 314638 300360 314644
rect 300596 204474 300624 315998
rect 300676 313880 300728 313886
rect 300676 313822 300728 313828
rect 300584 204468 300636 204474
rect 300584 204410 300636 204416
rect 300688 201482 300716 313822
rect 300780 204406 300808 325666
rect 301872 313948 301924 313954
rect 301872 313890 301924 313896
rect 301780 204876 301832 204882
rect 301780 204818 301832 204824
rect 301792 204542 301820 204818
rect 301780 204536 301832 204542
rect 301780 204478 301832 204484
rect 300768 204400 300820 204406
rect 300768 204342 300820 204348
rect 300768 204264 300820 204270
rect 300768 204206 300820 204212
rect 300676 201476 300728 201482
rect 300676 201418 300728 201424
rect 300676 188352 300728 188358
rect 300676 188294 300728 188300
rect 300584 185904 300636 185910
rect 300584 185846 300636 185852
rect 300596 78062 300624 185846
rect 300584 78056 300636 78062
rect 300584 77998 300636 78004
rect 300124 76628 300176 76634
rect 300124 76570 300176 76576
rect 300688 61674 300716 188294
rect 300780 69018 300808 204206
rect 301502 203552 301558 203561
rect 301502 203487 301558 203496
rect 301516 76634 301544 203487
rect 301792 200114 301820 204478
rect 301884 204406 301912 313890
rect 301872 204400 301924 204406
rect 301872 204342 301924 204348
rect 301976 203998 302004 331230
rect 301964 203992 302016 203998
rect 301964 203934 302016 203940
rect 301792 200086 301912 200114
rect 301504 76628 301556 76634
rect 301504 76570 301556 76576
rect 301688 75880 301740 75886
rect 301688 75822 301740 75828
rect 301700 75274 301728 75822
rect 301688 75268 301740 75274
rect 301688 75210 301740 75216
rect 301884 73166 301912 200086
rect 301976 75886 302004 203934
rect 302068 203930 302096 332250
rect 302160 331362 302188 332386
rect 302148 331356 302200 331362
rect 302148 331298 302200 331304
rect 303080 331294 303108 332454
rect 303172 332382 303200 459031
rect 303264 458046 303292 585754
rect 338868 583370 338896 587316
rect 338856 583364 338908 583370
rect 338856 583306 338908 583312
rect 343928 583302 343956 587316
rect 343916 583296 343968 583302
rect 343916 583238 343968 583244
rect 348988 583234 349016 587316
rect 348976 583228 349028 583234
rect 348976 583170 349028 583176
rect 354048 583166 354076 587316
rect 354036 583160 354088 583166
rect 354036 583102 354088 583108
rect 359108 583098 359136 587316
rect 359096 583092 359148 583098
rect 359096 583034 359148 583040
rect 364168 583030 364196 587316
rect 364156 583024 364208 583030
rect 369228 583001 369256 587316
rect 364156 582966 364208 582972
rect 369214 582992 369270 583001
rect 369214 582927 369270 582936
rect 374288 580582 374316 587316
rect 374276 580576 374328 580582
rect 374276 580518 374328 580524
rect 379348 580514 379376 587316
rect 379336 580508 379388 580514
rect 379336 580450 379388 580456
rect 384408 580378 384436 587316
rect 384396 580372 384448 580378
rect 384396 580314 384448 580320
rect 389468 580281 389496 587316
rect 394528 580446 394556 587316
rect 394516 580440 394568 580446
rect 394516 580382 394568 580388
rect 399588 580310 399616 587316
rect 404372 587302 404662 587330
rect 408512 587302 409722 587330
rect 414032 587302 414782 587330
rect 419552 587302 419842 587330
rect 399576 580304 399628 580310
rect 389454 580272 389510 580281
rect 399576 580246 399628 580252
rect 389454 580207 389510 580216
rect 404372 571985 404400 587302
rect 408512 577658 408540 587302
rect 408500 577652 408552 577658
rect 408500 577594 408552 577600
rect 414032 577590 414060 587302
rect 414020 577584 414072 577590
rect 414020 577526 414072 577532
rect 419552 577522 419580 587302
rect 424888 586498 424916 587316
rect 429948 586498 429976 587316
rect 434732 587302 435022 587330
rect 424876 586492 424928 586498
rect 424876 586434 424928 586440
rect 429936 586492 429988 586498
rect 429936 586434 429988 586440
rect 424888 585206 424916 586434
rect 424324 585200 424376 585206
rect 424324 585142 424376 585148
rect 424876 585200 424928 585206
rect 424876 585142 424928 585148
rect 419540 577516 419592 577522
rect 419540 577458 419592 577464
rect 404358 571976 404414 571985
rect 404358 571911 404414 571920
rect 424336 570625 424364 585142
rect 434732 571985 434760 587302
rect 440068 580281 440096 587316
rect 444392 587302 445142 587330
rect 440054 580272 440110 580281
rect 440054 580207 440110 580216
rect 444392 572014 444420 587302
rect 450188 580417 450216 587316
rect 450174 580408 450230 580417
rect 450174 580343 450230 580352
rect 455248 580310 455276 587316
rect 460308 580378 460336 587316
rect 465368 583030 465396 587316
rect 469232 587302 470442 587330
rect 465356 583024 465408 583030
rect 465356 582966 465408 582972
rect 460296 580372 460348 580378
rect 460296 580314 460348 580320
rect 455236 580304 455288 580310
rect 455236 580246 455288 580252
rect 469232 572082 469260 587302
rect 475488 580446 475516 587316
rect 480548 585721 480576 587316
rect 485608 585857 485636 587316
rect 485594 585848 485650 585857
rect 485594 585783 485650 585792
rect 480534 585712 480590 585721
rect 480534 585647 480590 585656
rect 490668 583001 490696 587316
rect 495452 587302 495742 587330
rect 490654 582992 490710 583001
rect 490654 582927 490710 582936
rect 475476 580440 475528 580446
rect 475476 580382 475528 580388
rect 495452 572150 495480 587302
rect 500788 583098 500816 587316
rect 505848 583137 505876 587316
rect 510908 583166 510936 587316
rect 515968 583234 515996 587316
rect 521028 585818 521056 587316
rect 525812 587302 526102 587330
rect 521016 585812 521068 585818
rect 521016 585754 521068 585760
rect 515956 583228 516008 583234
rect 515956 583170 516008 583176
rect 510896 583160 510948 583166
rect 505834 583128 505890 583137
rect 500776 583092 500828 583098
rect 510896 583102 510948 583108
rect 505834 583063 505890 583072
rect 500776 583034 500828 583040
rect 525812 572218 525840 587302
rect 531148 585886 531176 587316
rect 536208 585954 536236 587316
rect 541268 586022 541296 587316
rect 546328 586090 546356 587316
rect 546316 586084 546368 586090
rect 546316 586026 546368 586032
rect 541256 586016 541308 586022
rect 541256 585958 541308 585964
rect 536196 585948 536248 585954
rect 536196 585890 536248 585896
rect 531136 585880 531188 585886
rect 531136 585822 531188 585828
rect 551388 585721 551416 587316
rect 556448 585857 556476 587316
rect 556434 585848 556490 585857
rect 556434 585783 556490 585792
rect 551374 585712 551430 585721
rect 551374 585647 551430 585656
rect 561508 585206 561536 587316
rect 561496 585200 561548 585206
rect 566568 585177 566596 587316
rect 568856 586084 568908 586090
rect 568856 586026 568908 586032
rect 567476 586016 567528 586022
rect 567476 585958 567528 585964
rect 561496 585142 561548 585148
rect 566554 585168 566610 585177
rect 566554 585103 566610 585112
rect 525800 572212 525852 572218
rect 525800 572154 525852 572160
rect 495440 572144 495492 572150
rect 495440 572086 495492 572092
rect 469220 572076 469272 572082
rect 469220 572018 469272 572024
rect 444380 572008 444432 572014
rect 434718 571976 434774 571985
rect 444380 571950 444432 571956
rect 434718 571911 434774 571920
rect 424322 570616 424378 570625
rect 424322 570551 424378 570560
rect 303526 461952 303582 461961
rect 303462 461910 303526 461938
rect 303526 461887 303582 461896
rect 305090 461816 305146 461825
rect 305090 461751 305146 461760
rect 305104 460970 305132 461751
rect 399312 461650 399602 461666
rect 399300 461644 399602 461650
rect 399352 461638 399602 461644
rect 399300 461586 399352 461592
rect 305092 460964 305144 460970
rect 305092 460906 305144 460912
rect 303252 458040 303304 458046
rect 303252 457982 303304 457988
rect 303264 457638 303292 457982
rect 303252 457632 303304 457638
rect 303252 457574 303304 457580
rect 303252 457496 303304 457502
rect 303252 457438 303304 457444
rect 303160 332376 303212 332382
rect 303160 332318 303212 332324
rect 303068 331288 303120 331294
rect 303068 331230 303120 331236
rect 302148 329792 302200 329798
rect 302148 329734 302200 329740
rect 302240 329792 302292 329798
rect 302240 329734 302292 329740
rect 302160 204270 302188 329734
rect 302252 329594 302280 329734
rect 302240 329588 302292 329594
rect 302240 329530 302292 329536
rect 303068 318776 303120 318782
rect 303068 318718 303120 318724
rect 302882 313984 302938 313993
rect 302882 313919 302938 313928
rect 302896 204338 302924 313919
rect 303080 307737 303108 318718
rect 303066 307728 303122 307737
rect 303066 307663 303122 307672
rect 302884 204332 302936 204338
rect 302884 204274 302936 204280
rect 302148 204264 302200 204270
rect 302148 204206 302200 204212
rect 303172 204066 303200 332318
rect 303264 315858 303292 457438
rect 305000 456068 305052 456074
rect 305000 456010 305052 456016
rect 305012 455394 305040 456010
rect 305000 455388 305052 455394
rect 305000 455330 305052 455336
rect 305104 451274 305132 460906
rect 308508 459134 308536 461244
rect 313568 459542 313596 461244
rect 313556 459536 313608 459542
rect 313556 459478 313608 459484
rect 318628 459270 318656 461244
rect 318616 459264 318668 459270
rect 318616 459206 318668 459212
rect 323688 459202 323716 461244
rect 313280 459196 313332 459202
rect 313280 459138 313332 459144
rect 323676 459196 323728 459202
rect 323676 459138 323728 459144
rect 308496 459128 308548 459134
rect 313292 459105 313320 459138
rect 308496 459070 308548 459076
rect 313278 459096 313334 459105
rect 313278 459031 313334 459040
rect 328748 457978 328776 461244
rect 333808 458046 333836 461244
rect 338868 458114 338896 461244
rect 343928 460222 343956 461244
rect 347792 461230 349002 461258
rect 343916 460216 343968 460222
rect 343916 460158 343968 460164
rect 338856 458108 338908 458114
rect 338856 458050 338908 458056
rect 333796 458040 333848 458046
rect 333796 457982 333848 457988
rect 328736 457972 328788 457978
rect 328736 457914 328788 457920
rect 305012 451246 305132 451274
rect 305012 442921 305040 451246
rect 347792 444378 347820 461230
rect 354048 459338 354076 461244
rect 359108 460834 359136 461244
rect 359096 460828 359148 460834
rect 359096 460770 359148 460776
rect 354036 459332 354088 459338
rect 354036 459274 354088 459280
rect 364168 457502 364196 461244
rect 369228 458250 369256 461244
rect 374288 459406 374316 461244
rect 374276 459400 374328 459406
rect 374276 459342 374328 459348
rect 369216 458244 369268 458250
rect 369216 458186 369268 458192
rect 364156 457496 364208 457502
rect 364156 457438 364208 457444
rect 379348 456686 379376 461244
rect 384408 460902 384436 461244
rect 384396 460896 384448 460902
rect 384396 460838 384448 460844
rect 389468 459474 389496 461244
rect 391940 461032 391992 461038
rect 391940 460974 391992 460980
rect 391952 460902 391980 460974
rect 394528 460902 394556 461244
rect 404648 460970 404676 461244
rect 404636 460964 404688 460970
rect 404636 460906 404688 460912
rect 391940 460896 391992 460902
rect 391940 460838 391992 460844
rect 394516 460896 394568 460902
rect 394516 460838 394568 460844
rect 389456 459468 389508 459474
rect 389456 459410 389508 459416
rect 409708 456754 409736 461244
rect 414032 461230 414782 461258
rect 409696 456748 409748 456754
rect 409696 456690 409748 456696
rect 379336 456680 379388 456686
rect 379336 456622 379388 456628
rect 347780 444372 347832 444378
rect 347780 444314 347832 444320
rect 414032 443737 414060 461230
rect 419828 456074 419856 461244
rect 424888 459542 424916 461244
rect 429948 459542 429976 461244
rect 435008 459610 435036 461244
rect 434996 459604 435048 459610
rect 434996 459546 435048 459552
rect 438124 459604 438176 459610
rect 438124 459546 438176 459552
rect 424876 459536 424928 459542
rect 424876 459478 424928 459484
rect 429936 459536 429988 459542
rect 429936 459478 429988 459484
rect 424888 458250 424916 459478
rect 424324 458244 424376 458250
rect 424324 458186 424376 458192
rect 424876 458244 424928 458250
rect 424876 458186 424928 458192
rect 419816 456068 419868 456074
rect 419816 456010 419868 456016
rect 414018 443728 414074 443737
rect 414018 443663 414074 443672
rect 424336 443601 424364 458186
rect 438136 444378 438164 459546
rect 440068 455394 440096 461244
rect 445128 460902 445156 461244
rect 445116 460896 445168 460902
rect 445116 460838 445168 460844
rect 450188 459474 450216 461244
rect 455248 460193 455276 461244
rect 455234 460184 455290 460193
rect 455234 460119 455290 460128
rect 450176 459468 450228 459474
rect 450176 459410 450228 459416
rect 460308 459406 460336 461244
rect 460296 459400 460348 459406
rect 460296 459342 460348 459348
rect 465368 459338 465396 461244
rect 470428 460902 470456 461244
rect 474752 461230 475502 461258
rect 470416 460896 470468 460902
rect 470416 460838 470468 460844
rect 465356 459332 465408 459338
rect 465356 459274 465408 459280
rect 440056 455388 440108 455394
rect 440056 455330 440108 455336
rect 438124 444372 438176 444378
rect 438124 444314 438176 444320
rect 474752 444310 474780 461230
rect 480548 458833 480576 461244
rect 485608 458969 485636 461244
rect 485594 458960 485650 458969
rect 485594 458895 485650 458904
rect 480534 458824 480590 458833
rect 480534 458759 480590 458768
rect 490668 458153 490696 461244
rect 495728 460834 495756 461244
rect 495716 460828 495768 460834
rect 495716 460770 495768 460776
rect 500788 458250 500816 461244
rect 500776 458244 500828 458250
rect 500776 458186 500828 458192
rect 490654 458144 490710 458153
rect 505848 458114 505876 461244
rect 490654 458079 490710 458088
rect 505836 458108 505888 458114
rect 505836 458050 505888 458056
rect 510908 458046 510936 461244
rect 510896 458040 510948 458046
rect 510896 457982 510948 457988
rect 515968 457978 515996 461244
rect 521028 460766 521056 461244
rect 521016 460760 521068 460766
rect 521016 460702 521068 460708
rect 526088 460698 526116 461244
rect 526076 460692 526128 460698
rect 526076 460634 526128 460640
rect 531148 459270 531176 461244
rect 536208 460630 536236 461244
rect 536196 460624 536248 460630
rect 536196 460566 536248 460572
rect 531136 459264 531188 459270
rect 531136 459206 531188 459212
rect 515956 457972 516008 457978
rect 515956 457914 516008 457920
rect 541268 457910 541296 461244
rect 546328 459542 546356 461244
rect 546316 459536 546368 459542
rect 546316 459478 546368 459484
rect 551388 458833 551416 461244
rect 556158 459640 556214 459649
rect 556158 459575 556214 459584
rect 556172 459542 556200 459575
rect 556160 459536 556212 459542
rect 556160 459478 556212 459484
rect 556448 458862 556476 461244
rect 561508 459513 561536 461244
rect 565832 461230 566582 461258
rect 565726 461000 565782 461009
rect 565726 460935 565782 460944
rect 564898 460320 564954 460329
rect 564898 460255 564954 460264
rect 561494 459504 561550 459513
rect 561494 459439 561550 459448
rect 564440 459468 564492 459474
rect 564440 459410 564492 459416
rect 564452 459105 564480 459410
rect 564438 459096 564494 459105
rect 564438 459031 564494 459040
rect 556436 458856 556488 458862
rect 551374 458824 551430 458833
rect 556436 458798 556488 458804
rect 551374 458759 551430 458768
rect 541256 457904 541308 457910
rect 541256 457846 541308 457852
rect 564912 455394 564940 460255
rect 564900 455388 564952 455394
rect 564900 455330 564952 455336
rect 564912 454714 564940 455330
rect 564900 454708 564952 454714
rect 564900 454650 564952 454656
rect 565740 451274 565768 460935
rect 565556 451246 565768 451274
rect 565556 444378 565584 451246
rect 565544 444372 565596 444378
rect 565544 444314 565596 444320
rect 474740 444304 474792 444310
rect 474740 444246 474792 444252
rect 424322 443592 424378 443601
rect 424322 443527 424378 443536
rect 565556 443018 565584 444314
rect 565544 443012 565596 443018
rect 565544 442954 565596 442960
rect 565832 442921 565860 461230
rect 565910 458144 565966 458153
rect 565910 458079 565912 458088
rect 565964 458079 565966 458088
rect 565912 458050 565964 458056
rect 567488 457994 567516 585958
rect 568672 585948 568724 585954
rect 568672 585890 568724 585896
rect 567568 585812 567620 585818
rect 567568 585754 567620 585760
rect 567580 460934 567608 585754
rect 567660 583024 567712 583030
rect 567660 582966 567712 582972
rect 567672 480254 567700 582966
rect 567672 480226 567792 480254
rect 567580 460906 567700 460934
rect 567672 460766 567700 460906
rect 567660 460760 567712 460766
rect 567660 460702 567712 460708
rect 567488 457966 567608 457994
rect 567580 457910 567608 457966
rect 567568 457904 567620 457910
rect 567568 457846 567620 457852
rect 304998 442912 305054 442921
rect 304998 442847 305054 442856
rect 565818 442912 565874 442921
rect 565818 442847 565874 442856
rect 304262 333840 304318 333849
rect 304262 333775 304318 333784
rect 565726 333840 565782 333849
rect 565726 333775 565782 333784
rect 303448 332489 303476 333268
rect 303712 332784 303764 332790
rect 303712 332726 303764 332732
rect 303434 332480 303490 332489
rect 303434 332415 303490 332424
rect 303618 330576 303674 330585
rect 303618 330511 303620 330520
rect 303672 330511 303674 330520
rect 303620 330482 303672 330488
rect 303252 315852 303304 315858
rect 303252 315794 303304 315800
rect 303160 204060 303212 204066
rect 303160 204002 303212 204008
rect 302056 203924 302108 203930
rect 302056 203866 302108 203872
rect 301964 75880 302016 75886
rect 301964 75822 302016 75828
rect 302068 74526 302096 203866
rect 302240 200796 302292 200802
rect 302240 200738 302292 200744
rect 302252 187202 302280 200738
rect 302240 187196 302292 187202
rect 302240 187138 302292 187144
rect 303068 186380 303120 186386
rect 303068 186322 303120 186328
rect 302056 74520 302108 74526
rect 302056 74462 302108 74468
rect 301872 73160 301924 73166
rect 301872 73102 301924 73108
rect 300768 69012 300820 69018
rect 300768 68954 300820 68960
rect 303080 63034 303108 186322
rect 303172 74458 303200 204002
rect 303264 187542 303292 315794
rect 303632 313886 303660 330482
rect 303724 318782 303752 332726
rect 303712 318776 303764 318782
rect 303712 318718 303764 318724
rect 304276 318102 304304 333775
rect 305000 333668 305052 333674
rect 305000 333610 305052 333616
rect 304264 318096 304316 318102
rect 304264 318038 304316 318044
rect 305012 314634 305040 333610
rect 305092 333328 305144 333334
rect 501144 333328 501196 333334
rect 305092 333270 305144 333276
rect 305104 332654 305132 333270
rect 305092 332648 305144 332654
rect 305092 332590 305144 332596
rect 305000 314628 305052 314634
rect 305000 314570 305052 314576
rect 305012 313954 305040 314570
rect 305104 314022 305132 332590
rect 306380 332580 306432 332586
rect 306380 332522 306432 332528
rect 305184 318096 305236 318102
rect 305184 318038 305236 318044
rect 305092 314016 305144 314022
rect 305196 313993 305224 318038
rect 306392 316062 306420 332522
rect 308508 332246 308536 333268
rect 311256 332512 311308 332518
rect 311256 332454 311308 332460
rect 308496 332240 308548 332246
rect 308496 332182 308548 332188
rect 311268 332178 311296 332454
rect 313568 332314 313596 333268
rect 318628 332586 318656 333268
rect 318616 332580 318668 332586
rect 318616 332522 318668 332528
rect 323688 332382 323716 333268
rect 328748 332450 328776 333268
rect 333808 332518 333836 333268
rect 333796 332512 333848 332518
rect 333796 332454 333848 332460
rect 328736 332444 328788 332450
rect 328736 332386 328788 332392
rect 323676 332376 323728 332382
rect 323676 332318 323728 332324
rect 313556 332308 313608 332314
rect 313556 332250 313608 332256
rect 311256 332172 311308 332178
rect 311256 332114 311308 332120
rect 338868 329662 338896 333268
rect 343928 329730 343956 333268
rect 347792 333254 349002 333282
rect 343916 329724 343968 329730
rect 343916 329666 343968 329672
rect 338856 329656 338908 329662
rect 338856 329598 338908 329604
rect 306380 316056 306432 316062
rect 306380 315998 306432 316004
rect 347792 315654 347820 333254
rect 354048 331294 354076 333268
rect 358832 333254 359122 333282
rect 362972 333254 364182 333282
rect 368492 333254 369242 333282
rect 374012 333254 374302 333282
rect 378152 333254 379362 333282
rect 384040 333254 384422 333282
rect 389192 333254 389482 333282
rect 352564 331288 352616 331294
rect 352564 331230 352616 331236
rect 354036 331288 354088 331294
rect 354036 331230 354088 331236
rect 352576 315722 352604 331230
rect 358832 315790 358860 333254
rect 362972 315858 363000 333254
rect 368492 315926 368520 333254
rect 374012 331242 374040 333254
rect 373920 331214 374040 331242
rect 373920 329798 373948 331214
rect 373908 329792 373960 329798
rect 373908 329734 373960 329740
rect 378152 315994 378180 333254
rect 384040 332722 384068 333254
rect 384028 332716 384080 332722
rect 384028 332658 384080 332664
rect 378140 315988 378192 315994
rect 378140 315930 378192 315936
rect 368480 315920 368532 315926
rect 368480 315862 368532 315868
rect 362960 315852 363012 315858
rect 362960 315794 363012 315800
rect 358820 315784 358872 315790
rect 358820 315726 358872 315732
rect 352564 315716 352616 315722
rect 352564 315658 352616 315664
rect 347780 315648 347832 315654
rect 347780 315590 347832 315596
rect 389192 314634 389220 333254
rect 394528 331226 394556 333268
rect 394516 331220 394568 331226
rect 394516 331162 394568 331168
rect 399588 329118 399616 333268
rect 404648 331294 404676 333268
rect 408512 333254 409722 333282
rect 404636 331288 404688 331294
rect 404636 331230 404688 331236
rect 405740 331288 405792 331294
rect 405740 331230 405792 331236
rect 399576 329112 399628 329118
rect 399576 329054 399628 329060
rect 405752 318102 405780 331230
rect 408512 318782 408540 333254
rect 414768 330546 414796 333268
rect 419828 332654 419856 333268
rect 419816 332648 419868 332654
rect 419816 332590 419868 332596
rect 424888 332586 424916 333268
rect 429948 332586 429976 333268
rect 424324 332580 424376 332586
rect 424324 332522 424376 332528
rect 424876 332580 424928 332586
rect 424876 332522 424928 332528
rect 429936 332580 429988 332586
rect 429936 332522 429988 332528
rect 414756 330540 414808 330546
rect 414756 330482 414808 330488
rect 424336 319462 424364 332522
rect 435008 331226 435036 333268
rect 440082 333254 440188 333282
rect 440160 331242 440188 333254
rect 445128 332586 445156 333268
rect 449912 333254 450202 333282
rect 454052 333254 455262 333282
rect 459572 333254 460322 333282
rect 445116 332580 445168 332586
rect 445116 332522 445168 332528
rect 434996 331220 435048 331226
rect 440160 331214 440280 331242
rect 434996 331162 435048 331168
rect 440252 329798 440280 331214
rect 440240 329792 440292 329798
rect 440240 329734 440292 329740
rect 424324 319456 424376 319462
rect 424324 319398 424376 319404
rect 449912 318782 449940 333254
rect 408500 318776 408552 318782
rect 408500 318718 408552 318724
rect 449900 318776 449952 318782
rect 449900 318718 449952 318724
rect 405740 318096 405792 318102
rect 405740 318038 405792 318044
rect 454052 314634 454080 333254
rect 459572 318714 459600 333254
rect 465368 331294 465396 333268
rect 469232 333254 470442 333282
rect 475502 333266 475792 333282
rect 475502 333260 475804 333266
rect 475502 333254 475752 333260
rect 465356 331288 465408 331294
rect 465356 331230 465408 331236
rect 467104 331288 467156 331294
rect 467104 331230 467156 331236
rect 459560 318708 459612 318714
rect 459560 318650 459612 318656
rect 389180 314628 389232 314634
rect 389180 314570 389232 314576
rect 454040 314628 454092 314634
rect 454040 314570 454092 314576
rect 467116 314566 467144 331230
rect 469232 318102 469260 333254
rect 475752 333202 475804 333208
rect 480548 329089 480576 333268
rect 485608 331809 485636 333268
rect 489932 333254 490682 333282
rect 495452 333254 495742 333282
rect 500802 333276 501144 333282
rect 500802 333270 501196 333276
rect 500802 333254 501184 333270
rect 505112 333254 505862 333282
rect 510632 333254 510922 333282
rect 514772 333254 515982 333282
rect 520292 333254 521042 333282
rect 525812 333254 526102 333282
rect 529952 333254 531162 333282
rect 485594 331800 485650 331809
rect 485594 331735 485650 331744
rect 480534 329080 480590 329089
rect 480534 329015 480590 329024
rect 489932 318646 489960 333254
rect 489920 318640 489972 318646
rect 489920 318582 489972 318588
rect 469220 318096 469272 318102
rect 469220 318038 469272 318044
rect 495452 316033 495480 333254
rect 495438 316024 495494 316033
rect 505112 315994 505140 333254
rect 495438 315959 495494 315968
rect 505100 315988 505152 315994
rect 505100 315930 505152 315936
rect 510632 315926 510660 333254
rect 510620 315920 510672 315926
rect 510620 315862 510672 315868
rect 514772 315858 514800 333254
rect 514760 315852 514812 315858
rect 514760 315794 514812 315800
rect 520292 315790 520320 333254
rect 520280 315784 520332 315790
rect 520280 315726 520332 315732
rect 525812 315722 525840 333254
rect 525800 315716 525852 315722
rect 525800 315658 525852 315664
rect 529952 315654 529980 333254
rect 536208 332518 536236 333268
rect 536196 332512 536248 332518
rect 536196 332454 536248 332460
rect 541268 332450 541296 333268
rect 541256 332444 541308 332450
rect 541256 332386 541308 332392
rect 546328 332382 546356 333268
rect 546316 332376 546368 332382
rect 546316 332318 546368 332324
rect 551388 331809 551416 333268
rect 556448 331906 556476 333268
rect 561508 331974 561536 333268
rect 561496 331968 561548 331974
rect 561496 331910 561548 331916
rect 556436 331900 556488 331906
rect 556436 331842 556488 331848
rect 551374 331800 551430 331809
rect 551374 331735 551430 331744
rect 529940 315648 529992 315654
rect 529940 315590 529992 315596
rect 565740 314634 565768 333775
rect 566568 331401 566596 333268
rect 567580 332450 567608 457846
rect 567672 451274 567700 460702
rect 567764 459338 567792 480226
rect 568684 460934 568712 585890
rect 568764 585200 568816 585206
rect 568764 585142 568816 585148
rect 568592 460906 568712 460934
rect 568592 460630 568620 460906
rect 568580 460624 568632 460630
rect 568580 460566 568632 460572
rect 567752 459332 567804 459338
rect 567752 459274 567804 459280
rect 567764 458697 567792 459274
rect 567750 458688 567806 458697
rect 567750 458623 567806 458632
rect 567672 451246 567792 451274
rect 567658 433392 567714 433401
rect 567658 433327 567714 433336
rect 567568 332444 567620 332450
rect 567568 332386 567620 332392
rect 566554 331392 566610 331401
rect 566554 331327 566610 331336
rect 566462 331256 566518 331265
rect 565820 331220 565872 331226
rect 566462 331191 566518 331200
rect 565820 331162 565872 331168
rect 565832 330546 565860 331162
rect 565820 330540 565872 330546
rect 565820 330482 565872 330488
rect 566372 315988 566424 315994
rect 566372 315930 566424 315936
rect 566384 315897 566412 315930
rect 566370 315888 566426 315897
rect 566370 315823 566426 315832
rect 565728 314628 565780 314634
rect 565728 314570 565780 314576
rect 467104 314560 467156 314566
rect 467104 314502 467156 314508
rect 565740 314226 565768 314570
rect 565728 314220 565780 314226
rect 565728 314162 565780 314168
rect 566476 313993 566504 331191
rect 567108 315988 567160 315994
rect 567108 315930 567160 315936
rect 567120 314786 567148 315930
rect 567120 314758 567332 314786
rect 567304 314650 567332 314758
rect 567304 314622 567516 314650
rect 305092 313958 305144 313964
rect 305182 313984 305238 313993
rect 305000 313948 305052 313954
rect 305182 313919 305238 313928
rect 566462 313984 566518 313993
rect 566462 313919 566518 313928
rect 305000 313890 305052 313896
rect 303620 313880 303672 313886
rect 303620 313822 303672 313828
rect 303620 205964 303672 205970
rect 303620 205906 303672 205912
rect 303526 205592 303582 205601
rect 303462 205550 303526 205578
rect 303526 205527 303582 205536
rect 303632 202842 303660 205906
rect 303802 205864 303858 205873
rect 303802 205799 303858 205808
rect 565726 205864 565782 205873
rect 565726 205799 565782 205808
rect 303710 205728 303766 205737
rect 303710 205663 303766 205672
rect 303620 202836 303672 202842
rect 303620 202778 303672 202784
rect 303724 202722 303752 205663
rect 303816 202774 303844 205799
rect 564438 205592 564494 205601
rect 564438 205527 564494 205536
rect 305182 205048 305238 205057
rect 305182 204983 305238 204992
rect 305092 204944 305144 204950
rect 305092 204886 305144 204892
rect 303896 204468 303948 204474
rect 303896 204410 303948 204416
rect 303632 202694 303752 202722
rect 303804 202768 303856 202774
rect 303804 202710 303856 202716
rect 303252 187536 303304 187542
rect 303252 187478 303304 187484
rect 303264 186386 303292 187478
rect 303344 186992 303396 186998
rect 303344 186934 303396 186940
rect 303252 186380 303304 186386
rect 303252 186322 303304 186328
rect 303356 186130 303384 186934
rect 303264 186102 303384 186130
rect 303160 74452 303212 74458
rect 303160 74394 303212 74400
rect 303068 63028 303120 63034
rect 303068 62970 303120 62976
rect 300676 61668 300728 61674
rect 300676 61610 300728 61616
rect 299388 56568 299440 56574
rect 299388 56510 299440 56516
rect 299400 56234 299428 56510
rect 299388 56228 299440 56234
rect 299388 56170 299440 56176
rect 303264 56098 303292 186102
rect 303632 185881 303660 202694
rect 303908 200114 303936 204410
rect 305000 204400 305052 204406
rect 305000 204342 305052 204348
rect 303724 200086 303936 200114
rect 303724 186454 303752 200086
rect 303712 186448 303764 186454
rect 303712 186390 303764 186396
rect 305012 185910 305040 204342
rect 305104 187610 305132 204886
rect 305196 187649 305224 204983
rect 308508 204241 308536 205292
rect 308494 204232 308550 204241
rect 308494 204167 308550 204176
rect 313568 203930 313596 205292
rect 318628 203998 318656 205292
rect 323688 204066 323716 205292
rect 328748 204134 328776 205292
rect 333808 204202 333836 205292
rect 333796 204196 333848 204202
rect 333796 204138 333848 204144
rect 328736 204128 328788 204134
rect 328736 204070 328788 204076
rect 323676 204060 323728 204066
rect 323676 204002 323728 204008
rect 318616 203992 318668 203998
rect 318616 203934 318668 203940
rect 313556 203924 313608 203930
rect 313556 203866 313608 203872
rect 338868 201414 338896 205292
rect 343928 204270 343956 205292
rect 347792 205278 349002 205306
rect 343916 204264 343968 204270
rect 343916 204206 343968 204212
rect 338856 201408 338908 201414
rect 338856 201350 338908 201356
rect 305736 187672 305788 187678
rect 305182 187640 305238 187649
rect 305092 187604 305144 187610
rect 305182 187575 305238 187584
rect 305734 187640 305736 187649
rect 305788 187640 305790 187649
rect 305734 187575 305790 187584
rect 305092 187546 305144 187552
rect 347792 186998 347820 205278
rect 354048 204610 354076 205292
rect 354036 204604 354088 204610
rect 354036 204546 354088 204552
rect 359108 204542 359136 205292
rect 362972 205278 364182 205306
rect 368492 205278 369242 205306
rect 359096 204536 359148 204542
rect 359096 204478 359148 204484
rect 362972 187542 363000 205278
rect 368492 188358 368520 205278
rect 374288 200870 374316 205292
rect 379348 204474 379376 205292
rect 379336 204468 379388 204474
rect 379336 204410 379388 204416
rect 384408 204134 384436 205292
rect 389468 204406 389496 205292
rect 393332 205278 394542 205306
rect 398852 205278 399602 205306
rect 389456 204400 389508 204406
rect 389456 204342 389508 204348
rect 382280 204128 382332 204134
rect 382280 204070 382332 204076
rect 384396 204128 384448 204134
rect 384396 204070 384448 204076
rect 374276 200864 374328 200870
rect 374276 200806 374328 200812
rect 382292 200802 382320 204070
rect 382280 200796 382332 200802
rect 382280 200738 382332 200744
rect 368480 188352 368532 188358
rect 368480 188294 368532 188300
rect 393332 187610 393360 205278
rect 398852 187678 398880 205278
rect 404648 204270 404676 205292
rect 404636 204264 404688 204270
rect 404636 204206 404688 204212
rect 405924 204264 405976 204270
rect 405924 204206 405976 204212
rect 405936 202162 405964 204206
rect 409708 202774 409736 205292
rect 414768 202910 414796 205292
rect 419552 205278 419842 205306
rect 413560 202904 413612 202910
rect 413560 202846 413612 202852
rect 414756 202904 414808 202910
rect 414756 202846 414808 202852
rect 408500 202768 408552 202774
rect 408500 202710 408552 202716
rect 409696 202768 409748 202774
rect 409696 202710 409748 202716
rect 405924 202156 405976 202162
rect 405924 202098 405976 202104
rect 408512 198014 408540 202710
rect 413572 201482 413600 202846
rect 419552 202842 419580 205278
rect 424888 204270 424916 205292
rect 429948 204270 429976 205292
rect 434732 205278 435022 205306
rect 424324 204264 424376 204270
rect 424324 204206 424376 204212
rect 424876 204264 424928 204270
rect 424876 204206 424928 204212
rect 429936 204264 429988 204270
rect 429936 204206 429988 204212
rect 419540 202836 419592 202842
rect 419540 202778 419592 202784
rect 413284 201476 413336 201482
rect 413284 201418 413336 201424
rect 413560 201476 413612 201482
rect 413560 201418 413612 201424
rect 408500 198008 408552 198014
rect 408500 197950 408552 197956
rect 398840 187672 398892 187678
rect 398840 187614 398892 187620
rect 393320 187604 393372 187610
rect 393320 187546 393372 187552
rect 362960 187536 363012 187542
rect 362960 187478 363012 187484
rect 413296 186998 413324 201418
rect 347780 186992 347832 186998
rect 347780 186934 347832 186940
rect 413284 186992 413336 186998
rect 413284 186934 413336 186940
rect 419552 185910 419580 202778
rect 424336 189786 424364 204206
rect 424324 189780 424376 189786
rect 424324 189722 424376 189728
rect 434732 189038 434760 205278
rect 440068 202910 440096 205292
rect 445128 202910 445156 205292
rect 450188 204377 450216 205292
rect 450174 204368 450230 204377
rect 450174 204303 450230 204312
rect 440056 202904 440108 202910
rect 440056 202846 440108 202852
rect 440884 202904 440936 202910
rect 440884 202846 440936 202852
rect 445116 202904 445168 202910
rect 445116 202846 445168 202852
rect 446404 202904 446456 202910
rect 446404 202846 446456 202852
rect 440896 198694 440924 202846
rect 440884 198688 440936 198694
rect 440884 198630 440936 198636
rect 446416 198626 446444 202846
rect 455248 202230 455276 205292
rect 455236 202224 455288 202230
rect 455236 202166 455288 202172
rect 460308 200802 460336 205292
rect 465368 203250 465396 205292
rect 470428 204134 470456 205292
rect 475502 205278 476068 205306
rect 470416 204128 470468 204134
rect 470416 204070 470468 204076
rect 471336 204128 471388 204134
rect 471336 204070 471388 204076
rect 465356 203244 465408 203250
rect 465356 203186 465408 203192
rect 467748 203244 467800 203250
rect 467748 203186 467800 203192
rect 467760 201482 467788 203186
rect 467748 201476 467800 201482
rect 467748 201418 467800 201424
rect 471348 201414 471376 204070
rect 476040 203402 476068 205278
rect 476040 203374 476160 203402
rect 471336 201408 471388 201414
rect 471336 201350 471388 201356
rect 476132 201346 476160 203374
rect 476120 201340 476172 201346
rect 476120 201282 476172 201288
rect 460296 200796 460348 200802
rect 460296 200738 460348 200744
rect 480548 200705 480576 205292
rect 485608 203561 485636 205292
rect 489932 205278 490682 205306
rect 485594 203552 485650 203561
rect 485594 203487 485650 203496
rect 480534 200696 480590 200705
rect 480534 200631 480590 200640
rect 446404 198620 446456 198626
rect 446404 198562 446456 198568
rect 434720 189032 434772 189038
rect 434720 188974 434772 188980
rect 489932 188970 489960 205278
rect 495728 202910 495756 205292
rect 500788 203114 500816 205292
rect 505848 204338 505876 205292
rect 510908 204406 510936 205292
rect 515968 204474 515996 205292
rect 521042 205278 521700 205306
rect 526102 205278 526392 205306
rect 531162 205278 531544 205306
rect 521672 204542 521700 205278
rect 526364 204950 526392 205278
rect 526352 204944 526404 204950
rect 526352 204886 526404 204892
rect 531516 204610 531544 205278
rect 531504 204604 531556 204610
rect 531504 204546 531556 204552
rect 521660 204536 521712 204542
rect 521660 204478 521712 204484
rect 515956 204468 516008 204474
rect 515956 204410 516008 204416
rect 510896 204400 510948 204406
rect 510896 204342 510948 204348
rect 505836 204332 505888 204338
rect 505836 204274 505888 204280
rect 536208 204105 536236 205292
rect 541268 204270 541296 205292
rect 541256 204264 541308 204270
rect 541256 204206 541308 204212
rect 546328 204202 546356 205292
rect 546316 204196 546368 204202
rect 546316 204138 546368 204144
rect 536194 204096 536250 204105
rect 536194 204031 536250 204040
rect 551388 203590 551416 205292
rect 556448 203658 556476 205292
rect 561508 204134 561536 205292
rect 561496 204128 561548 204134
rect 561496 204070 561548 204076
rect 556436 203652 556488 203658
rect 556436 203594 556488 203600
rect 551376 203584 551428 203590
rect 551376 203526 551428 203532
rect 500776 203108 500828 203114
rect 500776 203050 500828 203056
rect 503628 203108 503680 203114
rect 503628 203050 503680 203056
rect 495716 202904 495768 202910
rect 495716 202846 495768 202852
rect 498568 202904 498620 202910
rect 498568 202846 498620 202852
rect 498580 201278 498608 202846
rect 498568 201272 498620 201278
rect 498568 201214 498620 201220
rect 503640 201210 503668 203050
rect 564452 202586 564480 205527
rect 564360 202558 564480 202586
rect 564360 202230 564388 202558
rect 564348 202224 564400 202230
rect 564348 202166 564400 202172
rect 560944 202156 560996 202162
rect 560944 202098 560996 202104
rect 503628 201204 503680 201210
rect 503628 201146 503680 201152
rect 489920 188964 489972 188970
rect 489920 188906 489972 188912
rect 560956 188358 560984 202098
rect 560944 188352 560996 188358
rect 560944 188294 560996 188300
rect 564360 187649 564388 202166
rect 565740 189038 565768 205799
rect 566568 203454 566596 205292
rect 567488 204338 567516 314622
rect 567476 204332 567528 204338
rect 567476 204274 567528 204280
rect 567580 204270 567608 332386
rect 567672 318782 567700 433327
rect 567660 318776 567712 318782
rect 567660 318718 567712 318724
rect 567672 306374 567700 318718
rect 567764 315790 567792 451246
rect 568592 332518 568620 460566
rect 568670 459640 568726 459649
rect 568670 459575 568726 459584
rect 568580 332512 568632 332518
rect 568580 332454 568632 332460
rect 567752 315784 567804 315790
rect 567752 315726 567804 315732
rect 567764 314702 567792 315726
rect 567752 314696 567804 314702
rect 567752 314638 567804 314644
rect 567672 306346 567884 306374
rect 567856 209774 567884 306346
rect 567856 209746 568068 209774
rect 568040 205698 568068 209746
rect 568028 205692 568080 205698
rect 568028 205634 568080 205640
rect 567660 204536 567712 204542
rect 567660 204478 567712 204484
rect 567568 204264 567620 204270
rect 567568 204206 567620 204212
rect 566556 203448 566608 203454
rect 566556 203390 566608 203396
rect 565728 189032 565780 189038
rect 565728 188974 565780 188980
rect 565740 188426 565768 188974
rect 565728 188420 565780 188426
rect 565728 188362 565780 188368
rect 564346 187640 564402 187649
rect 564346 187575 564402 187584
rect 305000 185904 305052 185910
rect 303618 185872 303674 185881
rect 305000 185846 305052 185852
rect 419540 185904 419592 185910
rect 419540 185846 419592 185852
rect 303618 185807 303674 185816
rect 332600 77920 332652 77926
rect 303526 77888 303582 77897
rect 303462 77846 303526 77874
rect 332600 77862 332652 77868
rect 336738 77888 336794 77897
rect 303526 77823 303582 77832
rect 308508 75857 308536 77316
rect 313292 77302 313582 77330
rect 308494 75848 308550 75857
rect 308494 75783 308550 75792
rect 308404 75472 308456 75478
rect 308404 75414 308456 75420
rect 307944 75268 307996 75274
rect 307944 75210 307996 75216
rect 307956 74534 307984 75210
rect 307864 74506 307984 74534
rect 307864 74458 307892 74506
rect 307852 74452 307904 74458
rect 307852 74394 307904 74400
rect 303712 71052 303764 71058
rect 303712 70994 303764 71000
rect 303252 56092 303304 56098
rect 303252 56034 303304 56040
rect 300400 54800 300452 54806
rect 300400 54742 300452 54748
rect 298836 53848 298888 53854
rect 298836 53790 298888 53796
rect 300412 52700 300440 54742
rect 303724 52714 303752 70994
rect 307760 61396 307812 61402
rect 307760 61338 307812 61344
rect 305920 57384 305972 57390
rect 305920 57326 305972 57332
rect 303724 52686 304106 52714
rect 305932 52700 305960 57326
rect 307772 52700 307800 61338
rect 307864 56166 307892 74394
rect 308416 61606 308444 75414
rect 313292 74526 313320 77302
rect 318628 75886 318656 77316
rect 318616 75880 318668 75886
rect 318616 75822 318668 75828
rect 319444 75336 319496 75342
rect 319444 75278 319496 75284
rect 313280 74520 313332 74526
rect 313280 74462 313332 74468
rect 308404 61600 308456 61606
rect 308404 61542 308456 61548
rect 309232 61532 309284 61538
rect 309232 61474 309284 61480
rect 309784 61532 309836 61538
rect 309784 61474 309836 61480
rect 307852 56160 307904 56166
rect 307852 56102 307904 56108
rect 309244 52714 309272 61474
rect 309796 54806 309824 61474
rect 311072 61464 311124 61470
rect 311072 61406 311124 61412
rect 309784 54800 309836 54806
rect 309784 54742 309836 54748
rect 311084 52714 311112 61406
rect 313292 60382 313320 74462
rect 317328 69896 317380 69902
rect 317328 69838 317380 69844
rect 313372 69760 313424 69766
rect 313372 69702 313424 69708
rect 313280 60376 313332 60382
rect 313280 60318 313332 60324
rect 313384 52714 313412 69702
rect 317340 69018 317368 69838
rect 316592 69012 316644 69018
rect 316592 68954 316644 68960
rect 317328 69012 317380 69018
rect 317328 68954 317380 68960
rect 309244 52686 309626 52714
rect 311084 52686 311466 52714
rect 313306 52686 313412 52714
rect 316604 52714 316632 68954
rect 319456 56574 319484 75278
rect 323688 75274 323716 77316
rect 328472 77302 328762 77330
rect 323676 75268 323728 75274
rect 323676 75210 323728 75216
rect 322204 73976 322256 73982
rect 322204 73918 322256 73924
rect 322296 73976 322348 73982
rect 322296 73918 322348 73924
rect 322112 73160 322164 73166
rect 322112 73102 322164 73108
rect 319444 56568 319496 56574
rect 319444 56510 319496 56516
rect 318800 56160 318852 56166
rect 318800 56102 318852 56108
rect 316604 52686 316986 52714
rect 318812 52700 318840 56102
rect 320640 56092 320692 56098
rect 320640 56034 320692 56040
rect 320652 52700 320680 56034
rect 322124 52714 322152 73102
rect 322216 54806 322244 73918
rect 322308 73166 322336 73918
rect 322296 73160 322348 73166
rect 322296 73102 322348 73108
rect 324320 63028 324372 63034
rect 324320 62970 324372 62976
rect 322204 54800 322256 54806
rect 322204 54742 322256 54748
rect 322124 52686 322506 52714
rect 324332 52700 324360 62970
rect 328472 62082 328500 77302
rect 329104 76764 329156 76770
rect 329104 76706 329156 76712
rect 329116 62082 329144 76706
rect 332612 75886 332640 77862
rect 336004 77852 336056 77858
rect 336738 77823 336794 77832
rect 454038 77888 454094 77897
rect 455326 77888 455382 77897
rect 455262 77846 455326 77874
rect 454038 77823 454094 77832
rect 455326 77823 455382 77832
rect 336004 77794 336056 77800
rect 332600 75880 332652 75886
rect 332600 75822 332652 75828
rect 332612 74534 332640 75822
rect 333808 75342 333836 77316
rect 333796 75336 333848 75342
rect 333796 75278 333848 75284
rect 332612 74506 333192 74534
rect 331220 71052 331272 71058
rect 331220 70994 331272 71000
rect 331232 70378 331260 70994
rect 331220 70372 331272 70378
rect 331220 70314 331272 70320
rect 331232 64874 331260 70314
rect 331232 64846 331352 64874
rect 329840 63096 329892 63102
rect 329840 63038 329892 63044
rect 328460 62076 328512 62082
rect 328460 62018 328512 62024
rect 329104 62076 329156 62082
rect 329104 62018 329156 62024
rect 325884 61668 325936 61674
rect 325884 61610 325936 61616
rect 325896 61402 325924 61610
rect 325884 61396 325936 61402
rect 325884 61338 325936 61344
rect 325896 52714 325924 61338
rect 329116 53854 329144 62018
rect 329852 57934 329880 63038
rect 329840 57928 329892 57934
rect 329840 57870 329892 57876
rect 328000 53848 328052 53854
rect 328000 53790 328052 53796
rect 329104 53848 329156 53854
rect 329104 53790 329156 53796
rect 325896 52686 326186 52714
rect 328012 52700 328040 53790
rect 329852 52700 329880 57870
rect 331324 52714 331352 64846
rect 333164 52714 333192 74506
rect 336016 67590 336044 77794
rect 336004 67584 336056 67590
rect 336004 67526 336056 67532
rect 336016 66842 336044 67526
rect 335360 66836 335412 66842
rect 335360 66778 335412 66784
rect 336004 66836 336056 66842
rect 336004 66778 336056 66784
rect 331324 52686 331706 52714
rect 333164 52686 333546 52714
rect 335372 52700 335400 66778
rect 336752 59362 336780 77823
rect 338224 77302 338882 77330
rect 338120 69760 338172 69766
rect 338120 69702 338172 69708
rect 336740 59356 336792 59362
rect 336740 59298 336792 59304
rect 336752 55214 336780 59298
rect 338132 55214 338160 69702
rect 338224 61538 338252 77302
rect 342352 74044 342404 74050
rect 342352 73986 342404 73992
rect 338212 61532 338264 61538
rect 338212 61474 338264 61480
rect 340880 60376 340932 60382
rect 340880 60318 340932 60324
rect 336752 55186 336872 55214
rect 338132 55186 338712 55214
rect 336844 52714 336872 55186
rect 338684 52714 338712 55186
rect 336844 52686 337226 52714
rect 338684 52686 339066 52714
rect 340892 52700 340920 60318
rect 342364 52714 342392 73986
rect 343928 69902 343956 77316
rect 347792 77302 349002 77330
rect 353312 77302 354062 77330
rect 343916 69896 343968 69902
rect 343916 69838 343968 69844
rect 346400 57316 346452 57322
rect 346400 57258 346452 57264
rect 344560 56024 344612 56030
rect 344560 55966 344612 55972
rect 342364 52686 342746 52714
rect 344572 52700 344600 55966
rect 346412 52700 346440 57258
rect 347792 56166 347820 77302
rect 349712 66972 349764 66978
rect 349712 66914 349764 66920
rect 347872 58676 347924 58682
rect 347872 58618 347924 58624
rect 347780 56160 347832 56166
rect 347780 56102 347832 56108
rect 347884 52714 347912 58618
rect 349724 52714 349752 66914
rect 353312 56098 353340 77302
rect 359108 73982 359136 77316
rect 362972 77302 364182 77330
rect 368584 77302 369242 77330
rect 374012 77302 374302 77330
rect 378152 77302 379362 77330
rect 359096 73976 359148 73982
rect 359096 73918 359148 73924
rect 357440 71120 357492 71126
rect 357440 71062 357492 71068
rect 353392 68400 353444 68406
rect 353392 68342 353444 68348
rect 353300 56092 353352 56098
rect 353300 56034 353352 56040
rect 351920 54800 351972 54806
rect 351920 54742 351972 54748
rect 347884 52686 348266 52714
rect 349724 52686 350106 52714
rect 351932 52700 351960 54742
rect 353404 52714 353432 68342
rect 355232 58744 355284 58750
rect 355232 58686 355284 58692
rect 355324 58744 355376 58750
rect 355324 58686 355376 58692
rect 355244 52714 355272 58686
rect 355336 54602 355364 58686
rect 355324 54596 355376 54602
rect 355324 54538 355376 54544
rect 353404 52686 353786 52714
rect 355244 52686 355626 52714
rect 357452 52700 357480 71062
rect 362972 63034 363000 77302
rect 366272 73908 366324 73914
rect 366272 73850 366324 73856
rect 364432 71188 364484 71194
rect 364432 71130 364484 71136
rect 362960 63028 363012 63034
rect 362960 62970 363012 62976
rect 362960 60172 363012 60178
rect 362960 60114 363012 60120
rect 360752 60104 360804 60110
rect 360752 60046 360804 60052
rect 358912 60036 358964 60042
rect 358912 59978 358964 59984
rect 358924 52714 358952 59978
rect 360764 52714 360792 60046
rect 358924 52686 359306 52714
rect 360764 52686 361146 52714
rect 362972 52700 363000 60114
rect 364444 52714 364472 71130
rect 366284 52714 366312 73850
rect 368480 69828 368532 69834
rect 368480 69770 368532 69776
rect 364444 52686 364826 52714
rect 366284 52686 366666 52714
rect 368492 52700 368520 69770
rect 368584 61402 368612 77302
rect 371792 72616 371844 72622
rect 371792 72558 371844 72564
rect 368572 61396 368624 61402
rect 368572 61338 368624 61344
rect 370320 57452 370372 57458
rect 370320 57394 370372 57400
rect 370332 52700 370360 57394
rect 371804 52714 371832 72558
rect 374012 62082 374040 77302
rect 376760 76628 376812 76634
rect 376760 76570 376812 76576
rect 376772 74534 376800 76570
rect 376772 74506 377352 74534
rect 375472 68536 375524 68542
rect 375472 68478 375524 68484
rect 374000 62076 374052 62082
rect 374000 62018 374052 62024
rect 374000 58812 374052 58818
rect 374000 58754 374052 58760
rect 371804 52686 372186 52714
rect 374012 52700 374040 58754
rect 375484 52714 375512 68478
rect 377324 52714 377352 74506
rect 378152 57934 378180 77302
rect 384408 71058 384436 77316
rect 386418 76664 386474 76673
rect 386418 76599 386474 76608
rect 385040 76016 385092 76022
rect 385040 75958 385092 75964
rect 384396 71052 384448 71058
rect 384396 70994 384448 71000
rect 378140 57928 378192 57934
rect 378140 57870 378192 57876
rect 383200 57520 383252 57526
rect 383200 57462 383252 57468
rect 381358 57352 381414 57361
rect 381358 57287 381414 57296
rect 379520 54732 379572 54738
rect 379520 54674 379572 54680
rect 375484 52686 375866 52714
rect 377324 52686 377706 52714
rect 379532 52700 379560 54674
rect 381372 52700 381400 57287
rect 383212 52700 383240 57462
rect 385052 52700 385080 75958
rect 386432 74534 386460 76599
rect 387798 76528 387854 76537
rect 387798 76463 387854 76472
rect 387812 74534 387840 76463
rect 389468 75886 389496 77316
rect 393332 77302 394542 77330
rect 398944 77302 399602 77330
rect 404464 77302 404662 77330
rect 409156 77302 409722 77330
rect 389456 75880 389508 75886
rect 389456 75822 389508 75828
rect 386432 74506 386552 74534
rect 387812 74506 388392 74534
rect 386524 52714 386552 74506
rect 388364 52714 388392 74506
rect 390560 73908 390612 73914
rect 390560 73850 390612 73856
rect 386524 52686 386906 52714
rect 388364 52686 388746 52714
rect 390572 52700 390600 73850
rect 393332 67590 393360 77302
rect 398838 76800 398894 76809
rect 398838 76735 398894 76744
rect 393320 67584 393372 67590
rect 393320 67526 393372 67532
rect 396080 60308 396132 60314
rect 396080 60250 396132 60256
rect 392032 58676 392084 58682
rect 392032 58618 392084 58624
rect 392044 52714 392072 58618
rect 394240 54664 394292 54670
rect 394240 54606 394292 54612
rect 392044 52686 392426 52714
rect 394252 52700 394280 54606
rect 396092 52700 396120 60250
rect 397552 60240 397604 60246
rect 397552 60182 397604 60188
rect 397564 52714 397592 60182
rect 398852 55214 398880 76735
rect 398944 59362 398972 77302
rect 404360 76628 404412 76634
rect 404360 76570 404412 76576
rect 403070 73808 403126 73817
rect 403070 73743 403126 73752
rect 401598 59936 401654 59945
rect 401598 59871 401654 59880
rect 398932 59356 398984 59362
rect 398932 59298 398984 59304
rect 398852 55186 399432 55214
rect 399404 52714 399432 55186
rect 397564 52686 397946 52714
rect 399404 52686 399786 52714
rect 401612 52700 401640 59871
rect 403084 52714 403112 73743
rect 404372 64874 404400 76570
rect 404464 69766 404492 77302
rect 408592 73976 408644 73982
rect 407118 73944 407174 73953
rect 408592 73918 408644 73924
rect 407118 73879 407174 73888
rect 405648 70372 405700 70378
rect 405648 70314 405700 70320
rect 405660 69766 405688 70314
rect 404452 69760 404504 69766
rect 404452 69702 404504 69708
rect 405648 69760 405700 69766
rect 405648 69702 405700 69708
rect 404372 64846 404952 64874
rect 404924 52714 404952 64846
rect 403084 52686 403466 52714
rect 404924 52686 405306 52714
rect 407132 52700 407160 73879
rect 408604 52714 408632 73918
rect 409156 69018 409184 77302
rect 414768 74594 414796 77316
rect 419842 77302 420224 77330
rect 418160 76696 418212 76702
rect 418160 76638 418212 76644
rect 414020 74588 414072 74594
rect 414020 74530 414072 74536
rect 414756 74588 414808 74594
rect 414756 74530 414808 74536
rect 414032 74050 414060 74530
rect 414020 74044 414072 74050
rect 414020 73986 414072 73992
rect 410432 69760 410484 69766
rect 410432 69702 410484 69708
rect 409144 69012 409196 69018
rect 409144 68954 409196 68960
rect 409156 60382 409184 68954
rect 409144 60376 409196 60382
rect 409144 60318 409196 60324
rect 410444 52714 410472 69702
rect 415952 61600 416004 61606
rect 415952 61542 416004 61548
rect 412640 61396 412692 61402
rect 412640 61338 412692 61344
rect 408604 52686 408986 52714
rect 410444 52686 410826 52714
rect 412652 52700 412680 61338
rect 414480 54528 414532 54534
rect 414480 54470 414532 54476
rect 414492 52700 414520 54470
rect 415964 52714 415992 61542
rect 415964 52686 416346 52714
rect 418172 52700 418200 76638
rect 420196 68921 420224 77302
rect 424888 75886 424916 77316
rect 429948 75886 429976 77316
rect 435022 77302 435404 77330
rect 430580 76696 430632 76702
rect 430580 76638 430632 76644
rect 423680 75880 423732 75886
rect 423680 75822 423732 75828
rect 424876 75880 424928 75886
rect 424876 75822 424928 75828
rect 429936 75880 429988 75886
rect 429936 75822 429988 75828
rect 423692 71262 423720 75822
rect 430592 74534 430620 76638
rect 430592 74506 430712 74534
rect 423680 71256 423732 71262
rect 423680 71198 423732 71204
rect 420182 68912 420238 68921
rect 420182 68847 420238 68856
rect 419998 57216 420054 57225
rect 419998 57151 420054 57160
rect 420012 52700 420040 57151
rect 420196 56030 420224 68847
rect 420184 56024 420236 56030
rect 420184 55966 420236 55972
rect 421838 54632 421894 54641
rect 421838 54567 421894 54576
rect 429200 54596 429252 54602
rect 421852 52700 421880 54567
rect 429200 54538 429252 54544
rect 427360 54528 427412 54534
rect 423678 54496 423734 54505
rect 423678 54431 423734 54440
rect 425518 54496 425574 54505
rect 427360 54470 427412 54476
rect 425518 54431 425574 54440
rect 423692 52700 423720 54431
rect 425532 52700 425560 54431
rect 427372 52700 427400 54470
rect 429212 52700 429240 54538
rect 430684 52714 430712 74506
rect 435376 73166 435404 77302
rect 439608 77302 440082 77330
rect 445036 77302 445142 77330
rect 450202 77302 450584 77330
rect 435364 73160 435416 73166
rect 435364 73102 435416 73108
rect 435376 62898 435404 73102
rect 439608 71738 439636 77302
rect 445036 73098 445064 77302
rect 445024 73092 445076 73098
rect 445024 73034 445076 73040
rect 439596 71732 439648 71738
rect 439596 71674 439648 71680
rect 435364 62892 435416 62898
rect 435364 62834 435416 62840
rect 439608 62830 439636 71674
rect 445036 62966 445064 73034
rect 450556 73030 450584 77302
rect 450544 73024 450596 73030
rect 450544 72966 450596 72972
rect 445024 62960 445076 62966
rect 445024 62902 445076 62908
rect 439596 62824 439648 62830
rect 439502 62792 439558 62801
rect 439596 62766 439648 62772
rect 439502 62727 439558 62736
rect 432512 58812 432564 58818
rect 432512 58754 432564 58760
rect 432524 52714 432552 58754
rect 439516 54602 439544 62727
rect 450556 55962 450584 72966
rect 450544 55956 450596 55962
rect 450544 55898 450596 55904
rect 454052 55894 454080 77823
rect 460308 72962 460336 77316
rect 465382 77302 465764 77330
rect 459560 72956 459612 72962
rect 459560 72898 459612 72904
rect 460296 72956 460348 72962
rect 460296 72898 460348 72904
rect 459572 72486 459600 72898
rect 459560 72480 459612 72486
rect 459560 72422 459612 72428
rect 465736 71777 465764 77302
rect 465722 71768 465778 71777
rect 465722 71703 465778 71712
rect 465736 64326 465764 71703
rect 470428 71670 470456 77316
rect 475396 77302 475502 77330
rect 480272 77302 480562 77330
rect 469864 71664 469916 71670
rect 469864 71606 469916 71612
rect 470416 71664 470468 71670
rect 470416 71606 470468 71612
rect 465724 64320 465776 64326
rect 465724 64262 465776 64268
rect 469876 64258 469904 71606
rect 475396 71602 475424 77302
rect 475384 71596 475436 71602
rect 475384 71538 475436 71544
rect 469864 64252 469916 64258
rect 469864 64194 469916 64200
rect 475396 64190 475424 71538
rect 480272 65686 480300 77302
rect 485608 73846 485636 77316
rect 490576 77302 490682 77330
rect 495742 77302 496124 77330
rect 485596 73840 485648 73846
rect 485596 73782 485648 73788
rect 490576 72894 490604 77302
rect 490564 72888 490616 72894
rect 490564 72830 490616 72836
rect 480260 65680 480312 65686
rect 480260 65622 480312 65628
rect 490576 65618 490604 72830
rect 496096 71534 496124 77302
rect 496084 71528 496136 71534
rect 496084 71470 496136 71476
rect 490564 65612 490616 65618
rect 490564 65554 490616 65560
rect 496096 65550 496124 71470
rect 500788 71466 500816 77316
rect 505848 75886 505876 77316
rect 510922 77302 511304 77330
rect 505836 75880 505888 75886
rect 505836 75822 505888 75828
rect 505848 75177 505876 75822
rect 511276 75818 511304 77302
rect 511264 75812 511316 75818
rect 511264 75754 511316 75760
rect 505834 75168 505890 75177
rect 505834 75103 505890 75112
rect 507032 74588 507084 74594
rect 507032 74530 507084 74536
rect 507044 73846 507072 74530
rect 507032 73840 507084 73846
rect 507032 73782 507084 73788
rect 500776 71460 500828 71466
rect 500776 71402 500828 71408
rect 500788 67046 500816 71402
rect 500776 67040 500828 67046
rect 500776 66982 500828 66988
rect 496084 65544 496136 65550
rect 496084 65486 496136 65492
rect 475384 64184 475436 64190
rect 475384 64126 475436 64132
rect 511276 58750 511304 75754
rect 515968 75750 515996 77316
rect 515956 75744 516008 75750
rect 515956 75686 516008 75692
rect 515968 75206 515996 75686
rect 521028 75682 521056 77316
rect 520280 75676 520332 75682
rect 520280 75618 520332 75624
rect 521016 75676 521068 75682
rect 521016 75618 521068 75624
rect 515956 75200 516008 75206
rect 515956 75142 516008 75148
rect 520292 68474 520320 75618
rect 526088 75614 526116 77316
rect 526076 75608 526128 75614
rect 526076 75550 526128 75556
rect 526088 69698 526116 75550
rect 531148 75546 531176 77316
rect 536116 77302 536222 77330
rect 529940 75540 529992 75546
rect 529940 75482 529992 75488
rect 531136 75540 531188 75546
rect 531136 75482 531188 75488
rect 529952 72554 529980 75482
rect 536116 74526 536144 77302
rect 536104 74520 536156 74526
rect 536104 74462 536156 74468
rect 534080 73840 534132 73846
rect 534080 73782 534132 73788
rect 534092 72826 534120 73782
rect 534080 72820 534132 72826
rect 534080 72762 534132 72768
rect 529940 72548 529992 72554
rect 529940 72490 529992 72496
rect 526076 69692 526128 69698
rect 526076 69634 526128 69640
rect 520280 68468 520332 68474
rect 520280 68410 520332 68416
rect 536116 66910 536144 74462
rect 541268 74458 541296 77316
rect 545776 77302 546342 77330
rect 550652 77302 551402 77330
rect 541256 74452 541308 74458
rect 541256 74394 541308 74400
rect 541268 68338 541296 74394
rect 545776 74390 545804 77302
rect 545764 74384 545816 74390
rect 545764 74326 545816 74332
rect 541256 68332 541308 68338
rect 541256 68274 541308 68280
rect 536104 66904 536156 66910
rect 536104 66846 536156 66852
rect 511264 58744 511316 58750
rect 511264 58686 511316 58692
rect 545776 57254 545804 74326
rect 550652 58682 550680 77302
rect 556448 69766 556476 77316
rect 561140 77302 561522 77330
rect 566108 77302 566582 77330
rect 561140 74534 561168 77302
rect 560956 74506 561168 74534
rect 560956 74322 560984 74506
rect 560944 74316 560996 74322
rect 560944 74258 560996 74264
rect 556436 69760 556488 69766
rect 556436 69702 556488 69708
rect 558182 69728 558238 69737
rect 558182 69663 558238 69672
rect 550640 58676 550692 58682
rect 550640 58618 550692 58624
rect 545764 57248 545816 57254
rect 545764 57190 545816 57196
rect 454040 55888 454092 55894
rect 454040 55830 454092 55836
rect 439504 54596 439556 54602
rect 439504 54538 439556 54544
rect 558196 54534 558224 69663
rect 560956 61402 560984 74258
rect 566108 64874 566136 77302
rect 567580 74458 567608 204206
rect 567672 75682 567700 204478
rect 568040 204377 568068 205634
rect 568026 204368 568082 204377
rect 567752 204332 567804 204338
rect 568026 204303 568082 204312
rect 567752 204274 567804 204280
rect 567764 75886 567792 204274
rect 568592 204105 568620 332454
rect 568684 332382 568712 459575
rect 568776 459513 568804 585142
rect 568868 459649 568896 586026
rect 569960 585880 570012 585886
rect 569960 585822 570012 585828
rect 571338 585848 571394 585857
rect 568948 583092 569000 583098
rect 568948 583034 569000 583040
rect 568854 459640 568910 459649
rect 568854 459575 568910 459584
rect 568762 459504 568818 459513
rect 568762 459439 568818 459448
rect 568672 332376 568724 332382
rect 568672 332318 568724 332324
rect 568684 204202 568712 332318
rect 568776 331974 568804 459439
rect 568960 458182 568988 583034
rect 569972 459270 570000 585822
rect 571338 585783 571394 585792
rect 570328 583228 570380 583234
rect 570328 583170 570380 583176
rect 570144 583160 570196 583166
rect 570144 583102 570196 583108
rect 570052 459808 570104 459814
rect 570052 459750 570104 459756
rect 569960 459264 570012 459270
rect 569960 459206 570012 459212
rect 569972 458250 570000 459206
rect 569960 458244 570012 458250
rect 569960 458186 570012 458192
rect 568948 458176 569000 458182
rect 568948 458118 569000 458124
rect 568856 443012 568908 443018
rect 568856 442954 568908 442960
rect 568764 331968 568816 331974
rect 568764 331910 568816 331916
rect 568868 330546 568896 442954
rect 569960 331900 570012 331906
rect 569960 331842 570012 331848
rect 568856 330540 568908 330546
rect 568856 330482 568908 330488
rect 568764 314696 568816 314702
rect 568764 314638 568816 314644
rect 568854 314664 568910 314673
rect 568776 204542 568804 314638
rect 568854 314599 568910 314608
rect 568868 314566 568896 314599
rect 568856 314560 568908 314566
rect 568856 314502 568908 314508
rect 568856 314220 568908 314226
rect 568856 314162 568908 314168
rect 568868 205601 568896 314162
rect 568854 205592 568910 205601
rect 568854 205527 568910 205536
rect 568764 204536 568816 204542
rect 568764 204478 568816 204484
rect 568672 204196 568724 204202
rect 568672 204138 568724 204144
rect 568578 204096 568634 204105
rect 568578 204031 568634 204040
rect 567752 75880 567804 75886
rect 567752 75822 567804 75828
rect 567660 75676 567712 75682
rect 567660 75618 567712 75624
rect 568592 74526 568620 204031
rect 568580 74520 568632 74526
rect 568580 74462 568632 74468
rect 567568 74452 567620 74458
rect 567568 74394 567620 74400
rect 568684 74390 568712 204138
rect 568764 203652 568816 203658
rect 568764 203594 568816 203600
rect 568672 74384 568724 74390
rect 568672 74326 568724 74332
rect 568776 73982 568804 203594
rect 568856 203448 568908 203454
rect 568856 203390 568908 203396
rect 568868 76702 568896 203390
rect 568856 76696 568908 76702
rect 568856 76638 568908 76644
rect 568764 73976 568816 73982
rect 569972 73953 570000 331842
rect 570064 315722 570092 459750
rect 570156 458046 570184 583102
rect 570236 572212 570288 572218
rect 570236 572154 570288 572160
rect 570248 460698 570276 572154
rect 570236 460692 570288 460698
rect 570236 460634 570288 460640
rect 570248 459814 570276 460634
rect 570236 459808 570288 459814
rect 570236 459750 570288 459756
rect 570144 458040 570196 458046
rect 570144 457982 570196 457988
rect 570156 315926 570184 457982
rect 570340 457978 570368 583170
rect 570604 458176 570656 458182
rect 570604 458118 570656 458124
rect 570328 457972 570380 457978
rect 570328 457914 570380 457920
rect 570340 456822 570368 457914
rect 570328 456816 570380 456822
rect 570328 456758 570380 456764
rect 570616 334014 570644 458118
rect 570604 334008 570656 334014
rect 570604 333950 570656 333956
rect 570616 333334 570644 333950
rect 570604 333328 570656 333334
rect 570604 333270 570656 333276
rect 570236 331968 570288 331974
rect 570236 331910 570288 331916
rect 570144 315920 570196 315926
rect 570144 315862 570196 315868
rect 570052 315716 570104 315722
rect 570052 315658 570104 315664
rect 570064 204950 570092 315658
rect 570156 314702 570184 315862
rect 570144 314696 570196 314702
rect 570144 314638 570196 314644
rect 570052 204944 570104 204950
rect 570052 204886 570104 204892
rect 570248 204134 570276 331910
rect 570328 314560 570380 314566
rect 570328 314502 570380 314508
rect 570236 204128 570288 204134
rect 570236 204070 570288 204076
rect 570052 203584 570104 203590
rect 570052 203526 570104 203532
rect 568764 73918 568816 73924
rect 569958 73944 570014 73953
rect 570064 73914 570092 203526
rect 570248 200114 570276 204070
rect 570340 201482 570368 314502
rect 570328 201476 570380 201482
rect 570328 201418 570380 201424
rect 570340 201385 570368 201418
rect 570326 201376 570382 201385
rect 570326 201311 570382 201320
rect 570156 200086 570276 200114
rect 570156 74322 570184 200086
rect 570236 185904 570288 185910
rect 570236 185846 570288 185852
rect 570248 79393 570276 185846
rect 570234 79384 570290 79393
rect 570234 79319 570290 79328
rect 570144 74316 570196 74322
rect 570144 74258 570196 74264
rect 569958 73879 570014 73888
rect 570052 73908 570104 73914
rect 570052 73850 570104 73856
rect 571352 73817 571380 585783
rect 574192 580440 574244 580446
rect 574192 580382 574244 580388
rect 572720 580372 572772 580378
rect 572720 580314 572772 580320
rect 571432 580304 571484 580310
rect 571432 580246 571484 580252
rect 571444 459649 571472 580246
rect 571524 572144 571576 572150
rect 571524 572086 571576 572092
rect 571536 460834 571564 572086
rect 571524 460828 571576 460834
rect 571524 460770 571576 460776
rect 571430 459640 571486 459649
rect 571536 459610 571564 460770
rect 571430 459575 571486 459584
rect 571524 459604 571576 459610
rect 571524 459546 571576 459552
rect 572732 459406 572760 580314
rect 572812 572076 572864 572082
rect 572812 572018 572864 572024
rect 572824 460902 572852 572018
rect 572812 460896 572864 460902
rect 572812 460838 572864 460844
rect 572824 459678 572852 460838
rect 572812 459672 572864 459678
rect 572812 459614 572864 459620
rect 574100 459672 574152 459678
rect 574100 459614 574152 459620
rect 572996 459604 573048 459610
rect 572996 459546 573048 459552
rect 572720 459400 572772 459406
rect 572720 459342 572772 459348
rect 571432 458856 571484 458862
rect 571432 458798 571484 458804
rect 571444 76634 571472 458798
rect 572732 458250 572760 459342
rect 571524 458244 571576 458250
rect 571524 458186 571576 458192
rect 572720 458244 572772 458250
rect 572720 458186 572772 458192
rect 571536 316062 571564 458186
rect 572812 456816 572864 456822
rect 572812 456758 572864 456764
rect 571616 454708 571668 454714
rect 571616 454650 571668 454656
rect 571628 329798 571656 454650
rect 571616 329792 571668 329798
rect 571616 329734 571668 329740
rect 571524 316056 571576 316062
rect 571524 315998 571576 316004
rect 571524 315920 571576 315926
rect 571524 315862 571576 315868
rect 571536 315654 571564 315862
rect 571524 315648 571576 315654
rect 571524 315590 571576 315596
rect 571524 314696 571576 314702
rect 571524 314638 571576 314644
rect 571536 204406 571564 314638
rect 571524 204400 571576 204406
rect 571524 204342 571576 204348
rect 571432 76628 571484 76634
rect 571432 76570 571484 76576
rect 571430 76120 571486 76129
rect 571430 76055 571486 76064
rect 571444 76022 571472 76055
rect 571432 76016 571484 76022
rect 571432 75958 571484 75964
rect 571536 75818 571564 204342
rect 571628 198694 571656 329734
rect 572824 325694 572852 456758
rect 572904 330540 572956 330546
rect 572904 330482 572956 330488
rect 572732 325666 572852 325694
rect 572732 315858 572760 325666
rect 572812 315988 572864 315994
rect 572812 315930 572864 315936
rect 572720 315852 572772 315858
rect 572720 315794 572772 315800
rect 572732 204814 572760 315794
rect 572720 204808 572772 204814
rect 572720 204750 572772 204756
rect 572732 204474 572760 204750
rect 572824 204610 572852 315930
rect 572916 205873 572944 330482
rect 573008 316033 573036 459546
rect 573364 318096 573416 318102
rect 573364 318038 573416 318044
rect 573376 317422 573404 318038
rect 574112 317422 574140 459614
rect 574204 444310 574232 580382
rect 575480 572008 575532 572014
rect 575480 571950 575532 571956
rect 575492 460970 575520 571950
rect 579618 524512 579674 524521
rect 577688 524476 577740 524482
rect 579618 524447 579620 524456
rect 577688 524418 577740 524424
rect 579672 524447 579674 524456
rect 579620 524418 579672 524424
rect 577504 484628 577556 484634
rect 577504 484570 577556 484576
rect 575480 460964 575532 460970
rect 575532 460912 575704 460934
rect 575480 460906 575704 460912
rect 575480 458244 575532 458250
rect 575480 458186 575532 458192
rect 574192 444304 574244 444310
rect 574192 444246 574244 444252
rect 574204 333266 574232 444246
rect 574468 334008 574520 334014
rect 574468 333950 574520 333956
rect 574192 333260 574244 333266
rect 574192 333202 574244 333208
rect 574204 332722 574232 333202
rect 574192 332716 574244 332722
rect 574192 332658 574244 332664
rect 573364 317416 573416 317422
rect 573364 317358 573416 317364
rect 574100 317416 574152 317422
rect 574100 317358 574152 317364
rect 572994 316024 573050 316033
rect 572994 315959 573050 315968
rect 573008 314809 573036 315959
rect 572994 314800 573050 314809
rect 572994 314735 573050 314744
rect 572902 205864 572958 205873
rect 572902 205799 572958 205808
rect 572904 204944 572956 204950
rect 572904 204886 572956 204892
rect 572812 204604 572864 204610
rect 572812 204546 572864 204552
rect 572720 204468 572772 204474
rect 572720 204410 572772 204416
rect 572720 201476 572772 201482
rect 572720 201418 572772 201424
rect 571616 198688 571668 198694
rect 571616 198630 571668 198636
rect 571524 75812 571576 75818
rect 571524 75754 571576 75760
rect 571338 73808 571394 73817
rect 571338 73743 571394 73752
rect 571628 71738 571656 198630
rect 571616 71732 571668 71738
rect 571616 71674 571668 71680
rect 572732 71670 572760 201418
rect 572824 75546 572852 204546
rect 572916 75614 572944 204886
rect 573376 201482 573404 317358
rect 574098 314800 574154 314809
rect 574098 314735 574154 314744
rect 573364 201476 573416 201482
rect 573364 201418 573416 201424
rect 574112 201278 574140 314735
rect 574284 204808 574336 204814
rect 574284 204750 574336 204756
rect 574100 201272 574152 201278
rect 574100 201214 574152 201220
rect 572996 188420 573048 188426
rect 572996 188362 573048 188368
rect 572904 75608 572956 75614
rect 572904 75550 572956 75556
rect 572812 75540 572864 75546
rect 572812 75482 572864 75488
rect 573008 73166 573036 188362
rect 572996 73160 573048 73166
rect 572996 73102 573048 73108
rect 572720 71664 572772 71670
rect 572720 71606 572772 71612
rect 574112 71534 574140 201214
rect 574192 198008 574244 198014
rect 574192 197950 574244 197956
rect 574204 79354 574232 197950
rect 574192 79348 574244 79354
rect 574192 79290 574244 79296
rect 574190 76528 574246 76537
rect 574190 76463 574246 76472
rect 574204 75954 574232 76463
rect 574192 75948 574244 75954
rect 574192 75890 574244 75896
rect 574296 75750 574324 204750
rect 574376 201476 574428 201482
rect 574376 201418 574428 201424
rect 574388 200802 574416 201418
rect 574480 201210 574508 333950
rect 575492 318714 575520 458186
rect 575570 457464 575626 457473
rect 575570 457399 575626 457408
rect 575480 318708 575532 318714
rect 575480 318650 575532 318656
rect 575492 201482 575520 318650
rect 575584 318646 575612 457399
rect 575676 332654 575704 460906
rect 575756 332716 575808 332722
rect 575756 332658 575808 332664
rect 575664 332648 575716 332654
rect 575664 332590 575716 332596
rect 575572 318640 575624 318646
rect 575572 318582 575624 318588
rect 575480 201476 575532 201482
rect 575480 201418 575532 201424
rect 574468 201204 574520 201210
rect 574468 201146 574520 201152
rect 574480 201074 574508 201146
rect 574468 201068 574520 201074
rect 574468 201010 574520 201016
rect 574376 200796 574428 200802
rect 574376 200738 574428 200744
rect 574284 75744 574336 75750
rect 574284 75686 574336 75692
rect 574388 72962 574416 200738
rect 575584 188970 575612 318582
rect 575676 198626 575704 332590
rect 575768 201346 575796 332658
rect 575756 201340 575808 201346
rect 575756 201282 575808 201288
rect 575768 200114 575796 201282
rect 575940 201068 575992 201074
rect 575940 201010 575992 201016
rect 575768 200086 575888 200114
rect 575664 198620 575716 198626
rect 575664 198562 575716 198568
rect 575572 188964 575624 188970
rect 575572 188906 575624 188912
rect 575584 187746 575612 188906
rect 575572 187740 575624 187746
rect 575572 187682 575624 187688
rect 574468 79348 574520 79354
rect 574468 79290 574520 79296
rect 574376 72956 574428 72962
rect 574376 72898 574428 72904
rect 574100 71528 574152 71534
rect 574100 71470 574152 71476
rect 574480 69018 574508 79290
rect 575676 73098 575704 198562
rect 575756 187740 575808 187746
rect 575756 187682 575808 187688
rect 575664 73092 575716 73098
rect 575664 73034 575716 73040
rect 575768 72894 575796 187682
rect 575756 72888 575808 72894
rect 575756 72830 575808 72836
rect 575860 71602 575888 200086
rect 575848 71596 575900 71602
rect 575848 71538 575900 71544
rect 575952 71466 575980 201010
rect 575940 71460 575992 71466
rect 575940 71402 575992 71408
rect 574468 69012 574520 69018
rect 574468 68954 574520 68960
rect 565832 64846 566136 64874
rect 560944 61396 560996 61402
rect 560944 61338 560996 61344
rect 565832 58818 565860 64846
rect 565820 58812 565872 58818
rect 565820 58754 565872 58760
rect 558184 54528 558236 54534
rect 558184 54470 558236 54476
rect 577516 53106 577544 484570
rect 577596 364744 577648 364750
rect 577596 364686 577648 364692
rect 577608 75857 577636 364686
rect 577700 318073 577728 524418
rect 580276 459134 580304 683839
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580264 459128 580316 459134
rect 580264 459070 580316 459076
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 577686 318064 577742 318073
rect 577686 317999 577742 318008
rect 578240 205692 578292 205698
rect 578240 205634 578292 205640
rect 577594 75848 577650 75857
rect 577594 75783 577650 75792
rect 578252 73030 578280 205634
rect 578332 188352 578384 188358
rect 578332 188294 578384 188300
rect 578240 73024 578292 73030
rect 578240 72966 578292 72972
rect 578344 70378 578372 188294
rect 579620 186992 579672 186998
rect 579620 186934 579672 186940
rect 579632 72826 579660 186934
rect 580276 76566 580304 378383
rect 580368 332489 580396 630799
rect 580920 591025 580948 643991
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580538 577688 580594 577697
rect 580538 577623 580594 577632
rect 580446 471472 580502 471481
rect 580446 471407 580502 471416
rect 580354 332480 580410 332489
rect 580354 332415 580410 332424
rect 580460 204241 580488 471407
rect 580552 332246 580580 577623
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 484673 580948 537775
rect 580630 484664 580686 484673
rect 580630 484599 580632 484608
rect 580684 484599 580686 484608
rect 580906 484664 580962 484673
rect 580906 484599 580962 484608
rect 580632 484570 580684 484576
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 378457 580948 431559
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580630 365120 580686 365129
rect 580630 365055 580686 365064
rect 580644 364750 580672 365055
rect 580632 364744 580684 364750
rect 580632 364686 580684 364692
rect 580540 332240 580592 332246
rect 580540 332182 580592 332188
rect 580446 204232 580502 204241
rect 580446 204167 580502 204176
rect 580264 76560 580316 76566
rect 580264 76502 580316 76508
rect 579620 72820 579672 72826
rect 579620 72762 579672 72768
rect 578332 70372 578384 70378
rect 578332 70314 578384 70320
rect 577504 53100 577556 53106
rect 577504 53042 577556 53048
rect 430684 52686 431066 52714
rect 432524 52686 432906 52714
rect 153106 38720 153162 38729
rect 153106 38655 153162 38664
rect 151726 38176 151782 38185
rect 151726 38111 151782 38120
rect 437386 37632 437442 37641
rect 437386 37567 437442 37576
rect 437400 37330 437428 37567
rect 437388 37324 437440 37330
rect 437388 37266 437440 37272
rect 565084 37324 565136 37330
rect 565084 37266 565136 37272
rect 151634 37224 151690 37233
rect 151634 37159 151690 37168
rect 151174 33144 151230 33153
rect 151174 33079 151230 33088
rect 151082 28520 151138 28529
rect 151082 28455 151138 28464
rect 151082 26480 151138 26489
rect 151082 26415 151138 26424
rect 3608 26240 3660 26246
rect 150440 26240 150492 26246
rect 3608 26182 3660 26188
rect 150438 26208 150440 26217
rect 150492 26208 150494 26217
rect 150438 26143 150494 26152
rect 127624 21412 127676 21418
rect 127624 21354 127676 21360
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 127636 2990 127664 21354
rect 138020 20052 138072 20058
rect 138020 19994 138072 20000
rect 135260 18896 135312 18902
rect 135260 18838 135312 18844
rect 131120 17468 131172 17474
rect 131120 17410 131172 17416
rect 131132 16574 131160 17410
rect 131132 16546 131344 16574
rect 129372 8968 129424 8974
rect 129372 8910 129424 8916
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 125876 2984 125928 2990
rect 125876 2926 125928 2932
rect 127624 2984 127676 2990
rect 127624 2926 127676 2932
rect 125888 480 125916 2926
rect 128188 480 128216 3402
rect 129384 480 129412 8910
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132960 7608 133012 7614
rect 132960 7550 133012 7556
rect 132972 480 133000 7550
rect 135272 480 135300 18838
rect 138032 16574 138060 19994
rect 142160 17536 142212 17542
rect 142160 17478 142212 17484
rect 138032 16546 138888 16574
rect 136456 9036 136508 9042
rect 136456 8978 136508 8984
rect 136468 480 136496 8978
rect 138860 480 138888 16546
rect 141424 10328 141476 10334
rect 141424 10270 141476 10276
rect 141436 3534 141464 10270
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 141424 3528 141476 3534
rect 141424 3470 141476 3476
rect 140056 480 140084 3470
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 17478
rect 145472 16244 145524 16250
rect 145472 16186 145524 16192
rect 143540 10396 143592 10402
rect 143540 10338 143592 10344
rect 143552 480 143580 10338
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16186
rect 151096 6866 151124 26415
rect 299584 23854 300518 23882
rect 214840 23792 214892 23798
rect 214498 23740 214840 23746
rect 214498 23734 214892 23740
rect 214498 23718 214880 23734
rect 243846 23730 244136 23746
rect 243846 23724 244148 23730
rect 243846 23718 244096 23724
rect 244096 23666 244148 23672
rect 266268 23656 266320 23662
rect 266110 23604 266268 23610
rect 266110 23598 266320 23604
rect 266110 23582 266308 23598
rect 267122 23594 267412 23610
rect 267122 23588 267424 23594
rect 267122 23582 267372 23588
rect 267372 23530 267424 23536
rect 269488 23520 269540 23526
rect 269146 23468 269488 23474
rect 277306 23488 277362 23497
rect 269146 23462 269540 23468
rect 269146 23446 269528 23462
rect 277242 23446 277306 23474
rect 277306 23423 277362 23432
rect 164332 21548 164384 21554
rect 164332 21490 164384 21496
rect 164344 16574 164372 21490
rect 164896 21418 164924 23324
rect 165724 23310 165922 23338
rect 166552 23310 166934 23338
rect 167012 23310 167946 23338
rect 168392 23310 168958 23338
rect 164884 21412 164936 21418
rect 164884 21354 164936 21360
rect 165620 19984 165672 19990
rect 165620 19926 165672 19932
rect 164344 16546 164464 16574
rect 163686 13016 163742 13025
rect 163686 12951 163742 12960
rect 151820 11960 151872 11966
rect 151820 11902 151872 11908
rect 151084 6860 151136 6866
rect 151084 6802 151136 6808
rect 150624 6248 150676 6254
rect 150624 6190 150676 6196
rect 147680 4820 147732 4826
rect 147680 4762 147732 4768
rect 147692 2802 147720 4762
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 147600 2774 147720 2802
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 354 147210 480
rect 147600 354 147628 2774
rect 149532 480 149560 3470
rect 150636 480 150664 6190
rect 151832 3602 151860 11902
rect 157800 11756 157852 11762
rect 157800 11698 157852 11704
rect 154212 7676 154264 7682
rect 154212 7618 154264 7624
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 153028 480 153056 3538
rect 154224 480 154252 7618
rect 156602 3360 156658 3369
rect 156602 3295 156658 3304
rect 156616 480 156644 3295
rect 157812 480 157840 11698
rect 160100 6180 160152 6186
rect 160100 6122 160152 6128
rect 160112 480 160140 6122
rect 161296 4888 161348 4894
rect 161296 4830 161348 4836
rect 161308 480 161336 4830
rect 163700 480 163728 12951
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 165632 7614 165660 19926
rect 165724 8974 165752 23310
rect 166552 19990 166580 23310
rect 166540 19984 166592 19990
rect 166540 19926 166592 19932
rect 167012 9042 167040 23310
rect 168392 10334 168420 23310
rect 169760 20120 169812 20126
rect 169760 20062 169812 20068
rect 168380 10328 168432 10334
rect 168380 10270 168432 10276
rect 167000 9036 167052 9042
rect 167000 8978 167052 8984
rect 165712 8968 165764 8974
rect 165712 8910 165764 8916
rect 165620 7608 165672 7614
rect 165620 7550 165672 7556
rect 168380 3936 168432 3942
rect 168380 3878 168432 3884
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 167196 480 167224 3538
rect 168392 480 168420 3878
rect 169772 490 169800 20062
rect 169852 19984 169904 19990
rect 169852 19926 169904 19932
rect 169864 4826 169892 19926
rect 169956 10402 169984 23324
rect 170600 23310 170982 23338
rect 171152 23310 171994 23338
rect 172532 23310 173006 23338
rect 170600 19990 170628 23310
rect 170588 19984 170640 19990
rect 170588 19926 170640 19932
rect 169944 10396 169996 10402
rect 169944 10338 169996 10344
rect 171152 6254 171180 23310
rect 171784 20732 171836 20738
rect 171784 20674 171836 20680
rect 171140 6248 171192 6254
rect 171140 6190 171192 6196
rect 169852 4820 169904 4826
rect 169852 4762 169904 4768
rect 171796 3942 171824 20674
rect 172532 7682 172560 23310
rect 173900 19984 173952 19990
rect 173900 19926 173952 19932
rect 172520 7676 172572 7682
rect 172520 7618 172572 7624
rect 173912 4894 173940 19926
rect 174004 11762 174032 23324
rect 174648 23310 175030 23338
rect 174544 20936 174596 20942
rect 174544 20878 174596 20884
rect 173992 11756 174044 11762
rect 173992 11698 174044 11704
rect 174268 9172 174320 9178
rect 174268 9114 174320 9120
rect 173900 4888 173952 4894
rect 173900 4830 173952 4836
rect 171784 3936 171836 3942
rect 171784 3878 171836 3884
rect 171968 3052 172020 3058
rect 171968 2994 172020 3000
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 169772 462 170352 490
rect 171980 480 172008 2994
rect 174280 480 174308 9114
rect 174556 3058 174584 20878
rect 174648 19990 174676 23310
rect 176028 21554 176056 23324
rect 176016 21548 176068 21554
rect 176016 21490 176068 21496
rect 177040 20738 177068 23324
rect 178052 20942 178080 23324
rect 178040 20936 178092 20942
rect 178040 20878 178092 20884
rect 178040 20800 178092 20806
rect 178040 20742 178092 20748
rect 177028 20732 177080 20738
rect 177028 20674 177080 20680
rect 177304 20732 177356 20738
rect 177304 20674 177356 20680
rect 176660 20188 176712 20194
rect 176660 20130 176712 20136
rect 174636 19984 174688 19990
rect 174636 19926 174688 19932
rect 175464 3664 175516 3670
rect 175464 3606 175516 3612
rect 174544 3052 174596 3058
rect 174544 2994 174596 3000
rect 175476 480 175504 3606
rect 176672 3398 176700 20130
rect 177316 3670 177344 20674
rect 178052 16574 178080 20742
rect 179064 20738 179092 23324
rect 180076 20806 180104 23324
rect 180064 20800 180116 20806
rect 180064 20742 180116 20748
rect 181088 20738 181116 23324
rect 182100 20806 182128 23324
rect 182088 20800 182140 20806
rect 182088 20742 182140 20748
rect 183112 20738 183140 23324
rect 184124 20874 184152 23324
rect 185044 23310 185150 23338
rect 185228 23310 186162 23338
rect 186332 23310 187174 23338
rect 187712 23310 188186 23338
rect 184112 20868 184164 20874
rect 184112 20810 184164 20816
rect 184204 20800 184256 20806
rect 184204 20742 184256 20748
rect 179052 20732 179104 20738
rect 179052 20674 179104 20680
rect 181076 20732 181128 20738
rect 181076 20674 181128 20680
rect 182180 20732 182232 20738
rect 182180 20674 182232 20680
rect 183100 20732 183152 20738
rect 183100 20674 183152 20680
rect 178052 16546 178632 16574
rect 177304 3664 177356 3670
rect 177304 3606 177356 3612
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177868 480 177896 3334
rect 170324 354 170352 462
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 181444 9104 181496 9110
rect 181444 9046 181496 9052
rect 181456 480 181484 9046
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 20674
rect 184216 3058 184244 20742
rect 184296 20732 184348 20738
rect 184296 20674 184348 20680
rect 184308 3330 184336 20674
rect 185044 7682 185072 23310
rect 185228 19938 185256 23310
rect 185584 20868 185636 20874
rect 185584 20810 185636 20816
rect 185136 19910 185256 19938
rect 185032 7676 185084 7682
rect 185032 7618 185084 7624
rect 185136 7614 185164 19910
rect 185216 18964 185268 18970
rect 185216 18906 185268 18912
rect 185124 7608 185176 7614
rect 185124 7550 185176 7556
rect 185228 6914 185256 18906
rect 184952 6886 185256 6914
rect 184296 3324 184348 3330
rect 184296 3266 184348 3272
rect 184204 3052 184256 3058
rect 184204 2994 184256 3000
rect 184952 480 184980 6886
rect 185596 4826 185624 20810
rect 186332 10402 186360 23310
rect 186320 10396 186372 10402
rect 186320 10338 186372 10344
rect 187712 10334 187740 23310
rect 189080 19984 189132 19990
rect 189080 19926 189132 19932
rect 189092 11762 189120 19926
rect 189184 11830 189212 23324
rect 189920 23310 190210 23338
rect 190472 23310 191222 23338
rect 191852 23310 192234 23338
rect 189920 19990 189948 23310
rect 189908 19984 189960 19990
rect 189908 19926 189960 19932
rect 190472 14618 190500 23310
rect 190460 14612 190512 14618
rect 190460 14554 190512 14560
rect 189172 11824 189224 11830
rect 189172 11766 189224 11772
rect 189080 11756 189132 11762
rect 189080 11698 189132 11704
rect 191852 10538 191880 23310
rect 193232 21554 193260 23324
rect 193324 23310 194258 23338
rect 194612 23310 195270 23338
rect 196084 23310 196282 23338
rect 196912 23310 197294 23338
rect 193220 21548 193272 21554
rect 193220 21490 193272 21496
rect 193324 13122 193352 23310
rect 194612 14550 194640 23310
rect 195980 19984 196032 19990
rect 195980 19926 196032 19932
rect 194600 14544 194652 14550
rect 194600 14486 194652 14492
rect 195992 14482 196020 19926
rect 196084 15978 196112 23310
rect 196912 19990 196940 23310
rect 196900 19984 196952 19990
rect 196900 19926 196952 19932
rect 198292 17338 198320 23324
rect 199304 21486 199332 23324
rect 200132 23310 200330 23338
rect 199292 21480 199344 21486
rect 199292 21422 199344 21428
rect 198280 17332 198332 17338
rect 198280 17274 198332 17280
rect 198740 16176 198792 16182
rect 198740 16118 198792 16124
rect 196072 15972 196124 15978
rect 196072 15914 196124 15920
rect 195980 14476 196032 14482
rect 195980 14418 196032 14424
rect 193312 13116 193364 13122
rect 193312 13058 193364 13064
rect 191840 10532 191892 10538
rect 191840 10474 191892 10480
rect 187700 10328 187752 10334
rect 187700 10270 187752 10276
rect 195612 9240 195664 9246
rect 195612 9182 195664 9188
rect 188528 6384 188580 6390
rect 188528 6326 188580 6332
rect 185584 4820 185636 4826
rect 185584 4762 185636 4768
rect 186136 3052 186188 3058
rect 186136 2994 186188 3000
rect 186148 480 186176 2994
rect 188540 480 188568 6326
rect 192024 5024 192076 5030
rect 192024 4966 192076 4972
rect 189724 3324 189776 3330
rect 189724 3266 189776 3272
rect 189736 480 189764 3266
rect 192036 480 192064 4966
rect 193220 4820 193272 4826
rect 193220 4762 193272 4768
rect 193232 480 193260 4762
rect 195624 480 195652 9182
rect 196808 7676 196860 7682
rect 196808 7618 196860 7624
rect 196820 480 196848 7618
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 16118
rect 200132 15910 200160 23310
rect 201328 17270 201356 23324
rect 201500 20256 201552 20262
rect 201500 20198 201552 20204
rect 201316 17264 201368 17270
rect 201316 17206 201368 17212
rect 200120 15904 200172 15910
rect 200120 15846 200172 15852
rect 200304 7608 200356 7614
rect 200304 7550 200356 7556
rect 200316 480 200344 7550
rect 201512 3398 201540 20198
rect 202340 18698 202368 23324
rect 202328 18692 202380 18698
rect 202328 18634 202380 18640
rect 203352 18630 203380 23324
rect 203340 18624 203392 18630
rect 203340 18566 203392 18572
rect 204260 16720 204312 16726
rect 204260 16662 204312 16668
rect 203432 10396 203484 10402
rect 203432 10338 203484 10344
rect 201500 3392 201552 3398
rect 201500 3334 201552 3340
rect 202696 3392 202748 3398
rect 202696 3334 202748 3340
rect 202708 480 202736 3334
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 10338
rect 204272 4826 204300 16662
rect 204364 4894 204392 23324
rect 205008 23310 205390 23338
rect 205652 23310 206402 23338
rect 207032 23310 207414 23338
rect 208426 23310 208532 23338
rect 205008 16726 205036 23310
rect 204996 16720 205048 16726
rect 204996 16662 205048 16668
rect 205652 6254 205680 23310
rect 206284 21412 206336 21418
rect 206284 21354 206336 21360
rect 206192 7812 206244 7818
rect 206192 7754 206244 7760
rect 205640 6248 205692 6254
rect 205640 6190 205692 6196
rect 204352 4888 204404 4894
rect 204352 4830 204404 4836
rect 204260 4820 204312 4826
rect 204260 4762 204312 4768
rect 206204 480 206232 7754
rect 206296 6186 206324 21354
rect 207032 7954 207060 23310
rect 208400 19984 208452 19990
rect 208400 19926 208452 19932
rect 207112 10328 207164 10334
rect 207112 10270 207164 10276
rect 207020 7948 207072 7954
rect 207020 7890 207072 7896
rect 206284 6180 206336 6186
rect 206284 6122 206336 6128
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 10270
rect 208412 7614 208440 19926
rect 208504 7682 208532 23310
rect 209056 23310 209438 23338
rect 209056 19990 209084 23310
rect 210332 21548 210384 21554
rect 210332 21490 210384 21496
rect 209044 19984 209096 19990
rect 209044 19926 209096 19932
rect 210344 12034 210372 21490
rect 210436 20738 210464 23324
rect 211448 21554 211476 23324
rect 211632 23310 212474 23338
rect 212552 23310 213486 23338
rect 211436 21548 211488 21554
rect 211436 21490 211488 21496
rect 210424 20732 210476 20738
rect 210424 20674 210476 20680
rect 210332 12028 210384 12034
rect 210332 11970 210384 11976
rect 209780 11824 209832 11830
rect 209780 11766 209832 11772
rect 209792 9674 209820 11766
rect 209872 10328 209924 10334
rect 209872 10270 209924 10276
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 208492 7676 208544 7682
rect 208492 7618 208544 7624
rect 208400 7608 208452 7614
rect 208400 7550 208452 7556
rect 209884 6914 209912 10270
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 211632 9314 211660 23310
rect 211804 20732 211856 20738
rect 211804 20674 211856 20680
rect 211620 9308 211672 9314
rect 211620 9250 211672 9256
rect 211816 5166 211844 20674
rect 212552 6186 212580 23310
rect 215496 22506 215524 23324
rect 215864 23310 216522 23338
rect 215484 22500 215536 22506
rect 215484 22442 215536 22448
rect 213368 14748 213420 14754
rect 213368 14690 213420 14696
rect 212540 6180 212592 6186
rect 212540 6122 212592 6128
rect 211804 5160 211856 5166
rect 211804 5102 211856 5108
rect 213380 480 213408 14690
rect 214472 11756 214524 11762
rect 214472 11698 214524 11704
rect 214484 480 214512 11698
rect 215864 6914 215892 23310
rect 217520 22438 217548 23324
rect 218164 23310 218546 23338
rect 217508 22432 217560 22438
rect 217508 22374 217560 22380
rect 218060 14612 218112 14618
rect 218060 14554 218112 14560
rect 215312 6886 215892 6914
rect 215312 2446 215340 6886
rect 216864 6452 216916 6458
rect 216864 6394 216916 6400
rect 215300 2440 215352 2446
rect 215300 2382 215352 2388
rect 216876 480 216904 6394
rect 218072 480 218100 14554
rect 218164 10470 218192 23310
rect 218152 10464 218204 10470
rect 218152 10406 218204 10412
rect 219544 10402 219572 23324
rect 220556 22370 220584 23324
rect 220832 23310 221582 23338
rect 222212 23310 222594 23338
rect 220544 22364 220596 22370
rect 220544 22306 220596 22312
rect 219992 13388 220044 13394
rect 219992 13330 220044 13336
rect 219532 10396 219584 10402
rect 219532 10338 219584 10344
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 13330
rect 220832 2378 220860 23310
rect 221096 10532 221148 10538
rect 221096 10474 221148 10480
rect 220820 2372 220872 2378
rect 220820 2314 220872 2320
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 10474
rect 222212 2310 222240 23310
rect 223592 11898 223620 23324
rect 223684 23310 224618 23338
rect 225064 23310 225630 23338
rect 223580 11892 223632 11898
rect 223580 11834 223632 11840
rect 223684 11830 223712 23310
rect 223672 11824 223724 11830
rect 223672 11766 223724 11772
rect 225064 11762 225092 23310
rect 226628 21690 226656 23324
rect 226904 23310 227654 23338
rect 226616 21684 226668 21690
rect 226616 21626 226668 21632
rect 225144 12028 225196 12034
rect 225144 11970 225196 11976
rect 225052 11756 225104 11762
rect 225052 11698 225104 11704
rect 223948 5092 224000 5098
rect 223948 5034 224000 5040
rect 222200 2304 222252 2310
rect 222200 2246 222252 2252
rect 223960 480 223988 5034
rect 225156 480 225184 11970
rect 226904 10305 226932 23310
rect 228652 22302 228680 23324
rect 229112 23310 229678 23338
rect 228640 22296 228692 22302
rect 228640 22238 228692 22244
rect 228364 21480 228416 21486
rect 228364 21422 228416 21428
rect 228376 16046 228404 21422
rect 228364 16040 228416 16046
rect 228364 15982 228416 15988
rect 229112 13326 229140 23310
rect 230676 21622 230704 23324
rect 230860 23310 231702 23338
rect 231964 23310 232714 23338
rect 233252 23310 233726 23338
rect 230664 21616 230716 21622
rect 230664 21558 230716 21564
rect 230480 17604 230532 17610
rect 230480 17546 230532 17552
rect 229100 13320 229152 13326
rect 229100 13262 229152 13268
rect 228272 13116 228324 13122
rect 228272 13058 228324 13064
rect 227536 12028 227588 12034
rect 227536 11970 227588 11976
rect 226890 10296 226946 10305
rect 226890 10231 226946 10240
rect 227548 480 227576 11970
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 13058
rect 230492 6914 230520 17546
rect 230860 13258 230888 23310
rect 231860 14544 231912 14550
rect 231860 14486 231912 14492
rect 230848 13252 230900 13258
rect 230848 13194 230900 13200
rect 230492 6886 231072 6914
rect 231044 480 231072 6886
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 231872 354 231900 14486
rect 231964 13190 231992 23310
rect 231952 13184 232004 13190
rect 231952 13126 232004 13132
rect 233252 13122 233280 23310
rect 234724 20874 234752 23324
rect 234908 23310 235750 23338
rect 236012 23310 236762 23338
rect 237484 23310 237774 23338
rect 238786 23310 238892 23338
rect 234712 20868 234764 20874
rect 234712 20810 234764 20816
rect 234620 15972 234672 15978
rect 234620 15914 234672 15920
rect 233240 13116 233292 13122
rect 233240 13058 233292 13064
rect 234632 3398 234660 15914
rect 234908 7750 234936 23310
rect 236012 14686 236040 23310
rect 237380 20324 237432 20330
rect 237380 20266 237432 20272
rect 236000 14680 236052 14686
rect 236000 14622 236052 14628
rect 234896 7744 234948 7750
rect 234896 7686 234948 7692
rect 237392 6914 237420 20266
rect 237484 14618 237512 23310
rect 237472 14612 237524 14618
rect 237472 14554 237524 14560
rect 238864 14550 238892 23310
rect 238956 23310 239798 23338
rect 240152 23310 240810 23338
rect 238852 14544 238904 14550
rect 238852 14486 238904 14492
rect 238956 14482 238984 23310
rect 240152 14521 240180 23310
rect 241808 22234 241836 23324
rect 241992 23310 242834 23338
rect 244292 23310 244858 23338
rect 241796 22228 241848 22234
rect 241796 22170 241848 22176
rect 240784 20868 240836 20874
rect 240784 20810 240836 20816
rect 240138 14512 240194 14521
rect 238944 14476 238996 14482
rect 240138 14447 240194 14456
rect 238944 14418 238996 14424
rect 239312 14408 239364 14414
rect 239312 14350 239364 14356
rect 237392 6886 237696 6914
rect 234712 3732 234764 3738
rect 234712 3674 234764 3680
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 234724 1850 234752 3674
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 234632 1822 234752 1850
rect 234632 480 234660 1822
rect 235828 480 235856 3334
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 6886
rect 239324 480 239352 14350
rect 240796 4962 240824 20810
rect 241992 11665 242020 23310
rect 242164 21480 242216 21486
rect 242164 21422 242216 21428
rect 242176 11966 242204 21422
rect 242900 17332 242952 17338
rect 242900 17274 242952 17280
rect 242164 11960 242216 11966
rect 242164 11902 242216 11908
rect 241978 11656 242034 11665
rect 241978 11591 242034 11600
rect 241704 10532 241756 10538
rect 241704 10474 241756 10480
rect 240784 4956 240836 4962
rect 240784 4898 240836 4904
rect 241716 480 241744 10474
rect 242912 480 242940 17274
rect 244292 16114 244320 23310
rect 245752 19984 245804 19990
rect 245752 19926 245804 19932
rect 244280 16108 244332 16114
rect 244280 16050 244332 16056
rect 245764 15978 245792 19926
rect 245856 16046 245884 23324
rect 246592 23310 246882 23338
rect 247052 23310 247894 23338
rect 248432 23310 248906 23338
rect 249812 23310 249918 23338
rect 246304 21684 246356 21690
rect 246304 21626 246356 21632
rect 245844 16040 245896 16046
rect 245844 15982 245896 15988
rect 245752 15972 245804 15978
rect 245752 15914 245804 15920
rect 244924 15904 244976 15910
rect 244924 15846 244976 15852
rect 245936 15904 245988 15910
rect 245936 15846 245988 15852
rect 244936 3058 244964 15846
rect 245200 6520 245252 6526
rect 245200 6462 245252 6468
rect 244924 3052 244976 3058
rect 244924 2994 244976 3000
rect 245212 480 245240 6462
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 15846
rect 246316 11966 246344 21626
rect 246592 19990 246620 23310
rect 246580 19984 246632 19990
rect 246580 19926 246632 19932
rect 247052 15910 247080 23310
rect 247682 21448 247738 21457
rect 247682 21383 247738 21392
rect 247696 16250 247724 21383
rect 247684 16244 247736 16250
rect 247684 16186 247736 16192
rect 247040 15904 247092 15910
rect 247040 15846 247092 15852
rect 246304 11960 246356 11966
rect 246304 11902 246356 11908
rect 248432 9081 248460 23310
rect 248788 9376 248840 9382
rect 248788 9318 248840 9324
rect 248418 9072 248474 9081
rect 248418 9007 248474 9016
rect 248800 480 248828 9318
rect 249812 2242 249840 23310
rect 250916 21758 250944 23324
rect 250904 21752 250956 21758
rect 250904 21694 250956 21700
rect 249984 21548 250036 21554
rect 249984 21490 250036 21496
rect 249996 20398 250024 21490
rect 249984 20392 250036 20398
rect 249984 20334 250036 20340
rect 251928 17406 251956 23324
rect 251916 17400 251968 17406
rect 251916 17342 251968 17348
rect 252940 17338 252968 23324
rect 252928 17332 252980 17338
rect 252928 17274 252980 17280
rect 253952 17270 253980 23324
rect 254032 21684 254084 21690
rect 254032 21626 254084 21632
rect 254044 17542 254072 21626
rect 254032 17536 254084 17542
rect 254032 17478 254084 17484
rect 252560 17264 252612 17270
rect 252560 17206 252612 17212
rect 253940 17264 253992 17270
rect 254964 17241 254992 23324
rect 255332 23310 255990 23338
rect 256804 23310 257002 23338
rect 253940 17206 253992 17212
rect 254950 17232 255006 17241
rect 252572 16574 252600 17206
rect 254950 17167 255006 17176
rect 252572 16546 253520 16574
rect 252468 7880 252520 7886
rect 252468 7822 252520 7828
rect 252480 3738 252508 7822
rect 252468 3732 252520 3738
rect 252468 3674 252520 3680
rect 252376 3664 252428 3670
rect 252376 3606 252428 3612
rect 249984 3052 250036 3058
rect 249984 2994 250036 3000
rect 249800 2236 249852 2242
rect 249800 2178 249852 2184
rect 249996 480 250024 2994
rect 252388 480 252416 3606
rect 253492 480 253520 16546
rect 255332 6361 255360 23310
rect 256700 18692 256752 18698
rect 256700 18634 256752 18640
rect 255318 6352 255374 6361
rect 255318 6287 255374 6296
rect 255872 2916 255924 2922
rect 255872 2858 255924 2864
rect 255884 480 255912 2858
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 18634
rect 256804 15881 256832 23310
rect 258000 18834 258028 23324
rect 257988 18828 258040 18834
rect 257988 18770 258040 18776
rect 259012 18766 259040 23324
rect 259000 18760 259052 18766
rect 259000 18702 259052 18708
rect 260024 18698 260052 23324
rect 260012 18692 260064 18698
rect 260012 18634 260064 18640
rect 261036 18630 261064 23324
rect 259460 18624 259512 18630
rect 259460 18566 259512 18572
rect 261024 18624 261076 18630
rect 262048 18601 262076 23324
rect 262864 21616 262916 21622
rect 262864 21558 262916 21564
rect 261024 18566 261076 18572
rect 262034 18592 262090 18601
rect 256790 15872 256846 15881
rect 256790 15807 256846 15816
rect 259472 3398 259500 18566
rect 262034 18527 262090 18536
rect 260104 14816 260156 14822
rect 260104 14758 260156 14764
rect 259552 3732 259604 3738
rect 259552 3674 259604 3680
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259564 1850 259592 3674
rect 260116 2922 260144 14758
rect 262876 13462 262904 21558
rect 263060 21554 263088 23324
rect 263612 23310 264086 23338
rect 263048 21548 263100 21554
rect 263048 21490 263100 21496
rect 262864 13456 262916 13462
rect 262864 13398 262916 13404
rect 262496 10600 262548 10606
rect 262496 10542 262548 10548
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 259472 1822 259592 1850
rect 259472 480 259500 1822
rect 260668 480 260696 3334
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 10542
rect 263612 2174 263640 23310
rect 265084 19961 265112 23324
rect 267936 23310 268134 23338
rect 269224 23310 270158 23338
rect 270512 23310 271170 23338
rect 271984 23310 272182 23338
rect 272904 23310 273194 23338
rect 273272 23310 274206 23338
rect 265070 19952 265126 19961
rect 265070 19887 265126 19896
rect 264152 4888 264204 4894
rect 264152 4830 264204 4836
rect 263600 2168 263652 2174
rect 263600 2110 263652 2116
rect 264164 480 264192 4830
rect 267740 4820 267792 4826
rect 267740 4762 267792 4768
rect 266544 3800 266596 3806
rect 266544 3742 266596 3748
rect 266556 480 266584 3742
rect 267752 480 267780 4762
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 267936 202 267964 23310
rect 269224 16574 269252 23310
rect 269132 16546 269252 16574
rect 269132 4894 269160 16546
rect 269210 7712 269266 7721
rect 269210 7647 269266 7656
rect 269120 4888 269172 4894
rect 269120 4830 269172 4836
rect 269224 3466 269252 7647
rect 270040 6588 270092 6594
rect 270040 6530 270092 6536
rect 269212 3460 269264 3466
rect 269212 3402 269264 3408
rect 270052 480 270080 6530
rect 270512 4826 270540 23310
rect 271880 19984 271932 19990
rect 271880 19926 271932 19932
rect 271236 6248 271288 6254
rect 271236 6190 271288 6196
rect 270500 4820 270552 4826
rect 270500 4762 270552 4768
rect 271248 480 271276 6190
rect 267924 196 267976 202
rect 267924 138 267976 144
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 271892 134 271920 19926
rect 271984 5001 272012 23310
rect 272904 19990 272932 23310
rect 272892 19984 272944 19990
rect 272892 19926 272944 19932
rect 271970 4992 272026 5001
rect 271970 4927 272026 4936
rect 273272 1358 273300 23310
rect 275204 22166 275232 23324
rect 275192 22160 275244 22166
rect 275192 22102 275244 22108
rect 276020 21752 276072 21758
rect 276020 21694 276072 21700
rect 276032 17542 276060 21694
rect 276216 21321 276244 23324
rect 277412 23310 278254 23338
rect 278792 23310 279266 23338
rect 280172 23310 280278 23338
rect 276202 21312 276258 21321
rect 276202 21247 276258 21256
rect 276020 17536 276072 17542
rect 276020 17478 276072 17484
rect 273904 16244 273956 16250
rect 273904 16186 273956 16192
rect 273916 3602 273944 16186
rect 276664 12096 276716 12102
rect 276664 12038 276716 12044
rect 274824 7948 274876 7954
rect 274824 7890 274876 7896
rect 273904 3596 273956 3602
rect 273904 3538 273956 3544
rect 273628 3460 273680 3466
rect 273628 3402 273680 3408
rect 273260 1352 273312 1358
rect 273260 1294 273312 1300
rect 273640 480 273668 3402
rect 274836 480 274864 7890
rect 271880 128 271932 134
rect 271880 70 271932 76
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 12038
rect 277412 6322 277440 23310
rect 278688 21752 278740 21758
rect 278688 21694 278740 21700
rect 278136 21548 278188 21554
rect 278136 21490 278188 21496
rect 278148 19990 278176 21490
rect 278700 20058 278728 21694
rect 278688 20052 278740 20058
rect 278688 19994 278740 20000
rect 278136 19984 278188 19990
rect 278136 19926 278188 19932
rect 277492 7948 277544 7954
rect 277492 7890 277544 7896
rect 277400 6316 277452 6322
rect 277400 6258 277452 6264
rect 277504 3534 277532 7890
rect 278320 7676 278372 7682
rect 278320 7618 278372 7624
rect 277492 3528 277544 3534
rect 277492 3470 277544 3476
rect 278332 480 278360 7618
rect 278792 6254 278820 23310
rect 279424 21548 279476 21554
rect 279424 21490 279476 21496
rect 279436 6594 279464 21490
rect 279424 6588 279476 6594
rect 279424 6530 279476 6536
rect 278780 6248 278832 6254
rect 278780 6190 278832 6196
rect 280068 6180 280120 6186
rect 280068 6122 280120 6128
rect 280080 3505 280108 6122
rect 280066 3496 280122 3505
rect 280066 3431 280122 3440
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280172 66 280200 23310
rect 281276 22137 281304 23324
rect 281552 23310 282302 23338
rect 282932 23310 283314 23338
rect 281262 22128 281318 22137
rect 281262 22063 281318 22072
rect 280712 10668 280764 10674
rect 280712 10610 280764 10616
rect 280724 480 280752 10610
rect 281552 2106 281580 23310
rect 281908 7608 281960 7614
rect 281908 7550 281960 7556
rect 281540 2100 281592 2106
rect 281540 2042 281592 2048
rect 281920 480 281948 7550
rect 282932 4865 282960 23310
rect 284312 6186 284340 23324
rect 284404 23310 285338 23338
rect 285692 23310 286350 23338
rect 287164 23310 287362 23338
rect 287992 23310 288374 23338
rect 284404 16574 284432 23310
rect 284404 16546 284524 16574
rect 284392 8968 284444 8974
rect 284392 8910 284444 8916
rect 284300 6180 284352 6186
rect 284300 6122 284352 6128
rect 282918 4856 282974 4865
rect 282918 4791 282974 4800
rect 284404 3482 284432 8910
rect 284496 7682 284524 16546
rect 284484 7676 284536 7682
rect 284484 7618 284536 7624
rect 285692 7614 285720 23310
rect 287060 19916 287112 19922
rect 287060 19858 287112 19864
rect 285680 7608 285732 7614
rect 285680 7550 285732 7556
rect 285404 5160 285456 5166
rect 285404 5102 285456 5108
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 285416 480 285444 5102
rect 287072 2009 287100 19858
rect 287164 7585 287192 23310
rect 287992 19922 288020 23310
rect 288440 20392 288492 20398
rect 288440 20334 288492 20340
rect 287980 19916 288032 19922
rect 287980 19858 288032 19864
rect 288452 16574 288480 20334
rect 289372 17377 289400 23324
rect 289832 23310 290398 23338
rect 291304 23310 291410 23338
rect 291488 23310 292422 23338
rect 292592 23310 293434 23338
rect 293972 23310 294446 23338
rect 289358 17368 289414 17377
rect 289358 17303 289414 17312
rect 288452 16546 289032 16574
rect 287150 7576 287206 7585
rect 287150 7511 287206 7520
rect 287796 3528 287848 3534
rect 287796 3470 287848 3476
rect 287058 2000 287114 2009
rect 287058 1935 287114 1944
rect 287808 480 287836 3470
rect 289004 480 289032 16546
rect 289832 6225 289860 23310
rect 291200 20052 291252 20058
rect 291200 19994 291252 20000
rect 291212 6914 291240 19994
rect 291304 9042 291332 23310
rect 291292 9036 291344 9042
rect 291292 8978 291344 8984
rect 291488 8945 291516 23310
rect 291844 21820 291896 21826
rect 291844 21762 291896 21768
rect 291856 8974 291884 21762
rect 292592 16574 292620 23310
rect 292592 16546 292712 16574
rect 292580 9308 292632 9314
rect 292580 9250 292632 9256
rect 291844 8968 291896 8974
rect 291474 8936 291530 8945
rect 291844 8910 291896 8916
rect 291474 8871 291530 8880
rect 291212 6886 291424 6914
rect 289818 6216 289874 6225
rect 289818 6151 289874 6160
rect 291396 480 291424 6886
rect 292592 480 292620 9250
rect 292684 8974 292712 16546
rect 292672 8968 292724 8974
rect 292672 8910 292724 8916
rect 293972 7721 294000 23310
rect 295444 17474 295472 23324
rect 296456 18902 296484 23324
rect 297364 21888 297416 21894
rect 297364 21830 297416 21836
rect 296444 18896 296496 18902
rect 296444 18838 296496 18844
rect 295432 17468 295484 17474
rect 295432 17410 295484 17416
rect 297376 9178 297404 21830
rect 297468 21758 297496 23324
rect 297456 21752 297508 21758
rect 297456 21694 297508 21700
rect 298480 21622 298508 23324
rect 298468 21616 298520 21622
rect 298468 21558 298520 21564
rect 299492 21457 299520 23324
rect 299478 21448 299534 21457
rect 299478 21383 299534 21392
rect 298744 20732 298796 20738
rect 298744 20674 298796 20680
rect 298100 18896 298152 18902
rect 298100 18838 298152 18844
rect 297364 9172 297416 9178
rect 297364 9114 297416 9120
rect 293958 7712 294014 7721
rect 293958 7647 294014 7656
rect 294880 3596 294932 3602
rect 294880 3538 294932 3544
rect 294892 480 294920 3538
rect 296074 3496 296130 3505
rect 296074 3431 296130 3440
rect 296088 480 296116 3431
rect 280160 60 280212 66
rect 280160 2 280212 8
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 18838
rect 298756 13025 298784 20674
rect 298742 13016 298798 13025
rect 298742 12951 298798 12960
rect 299584 7954 299612 23854
rect 299664 23792 299716 23798
rect 299664 23734 299716 23740
rect 299572 7948 299624 7954
rect 299572 7890 299624 7896
rect 299676 480 299704 23734
rect 336004 23724 336056 23730
rect 336004 23666 336056 23672
rect 301412 22500 301464 22506
rect 301412 22442 301464 22448
rect 300952 21140 301004 21146
rect 300952 21082 301004 21088
rect 300964 20126 300992 21082
rect 300952 20120 301004 20126
rect 300952 20062 301004 20068
rect 301424 16574 301452 22442
rect 301516 21486 301544 23324
rect 302344 23310 302542 23338
rect 301504 21480 301556 21486
rect 301504 21422 301556 21428
rect 301596 20392 301648 20398
rect 301596 20334 301648 20340
rect 301424 16546 301544 16574
rect 300492 8220 300544 8226
rect 300492 8162 300544 8168
rect 300504 3369 300532 8162
rect 301516 3505 301544 16546
rect 301608 3738 301636 20334
rect 302344 8226 302372 23310
rect 303540 21418 303568 23324
rect 304264 21480 304316 21486
rect 304264 21422 304316 21428
rect 303528 21412 303580 21418
rect 303528 21354 303580 21360
rect 302884 21344 302936 21350
rect 302884 21286 302936 21292
rect 302332 8220 302384 8226
rect 302332 8162 302384 8168
rect 302896 6390 302924 21286
rect 302884 6384 302936 6390
rect 302884 6326 302936 6332
rect 304276 5030 304304 21422
rect 304552 20738 304580 23324
rect 305012 23310 305578 23338
rect 304540 20732 304592 20738
rect 304540 20674 304592 20680
rect 305012 16250 305040 23310
rect 306576 21146 306604 23324
rect 307588 21758 307616 23324
rect 307576 21752 307628 21758
rect 307576 21694 307628 21700
rect 306564 21140 306616 21146
rect 306564 21082 306616 21088
rect 308600 21010 308628 23324
rect 309232 22432 309284 22438
rect 309232 22374 309284 22380
rect 306564 21004 306616 21010
rect 306564 20946 306616 20952
rect 308588 21004 308640 21010
rect 308588 20946 308640 20952
rect 306576 20194 306604 20946
rect 307116 20732 307168 20738
rect 307116 20674 307168 20680
rect 306564 20188 306616 20194
rect 306564 20130 306616 20136
rect 305000 16244 305052 16250
rect 305000 16186 305052 16192
rect 307024 16244 307076 16250
rect 307024 16186 307076 16192
rect 305644 10464 305696 10470
rect 305644 10406 305696 10412
rect 305552 7948 305604 7954
rect 305552 7890 305604 7896
rect 304264 5024 304316 5030
rect 304264 4966 304316 4972
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 301596 3732 301648 3738
rect 301596 3674 301648 3680
rect 301502 3496 301558 3505
rect 301502 3431 301558 3440
rect 300490 3360 300546 3369
rect 300490 3295 300546 3304
rect 301976 480 302004 3810
rect 303158 3496 303214 3505
rect 303158 3431 303214 3440
rect 303172 480 303200 3431
rect 305564 480 305592 7890
rect 305656 3369 305684 10406
rect 307036 3670 307064 16186
rect 307128 9110 307156 20674
rect 307116 9104 307168 9110
rect 307116 9046 307168 9052
rect 307760 9104 307812 9110
rect 307760 9046 307812 9052
rect 307772 3806 307800 9046
rect 309244 6914 309272 22374
rect 309612 20738 309640 23324
rect 309784 21208 309836 21214
rect 309784 21150 309836 21156
rect 309600 20732 309652 20738
rect 309600 20674 309652 20680
rect 309796 14754 309824 21150
rect 310624 18970 310652 23324
rect 311636 21418 311664 23324
rect 312648 21486 312676 23324
rect 313292 23310 313674 23338
rect 312636 21480 312688 21486
rect 312636 21422 312688 21428
rect 311624 21412 311676 21418
rect 311624 21354 311676 21360
rect 311164 21344 311216 21350
rect 311164 21286 311216 21292
rect 310612 18964 310664 18970
rect 310612 18906 310664 18912
rect 309784 14748 309836 14754
rect 309784 14690 309836 14696
rect 311176 7818 311204 21286
rect 312544 21276 312596 21282
rect 312544 21218 312596 21224
rect 311256 20732 311308 20738
rect 311256 20674 311308 20680
rect 311268 16182 311296 20674
rect 311256 16176 311308 16182
rect 311256 16118 311308 16124
rect 311164 7812 311216 7818
rect 311164 7754 311216 7760
rect 309244 6886 309824 6914
rect 307760 3800 307812 3806
rect 307760 3742 307812 3748
rect 307024 3664 307076 3670
rect 307024 3606 307076 3612
rect 309048 3664 309100 3670
rect 309048 3606 309100 3612
rect 305642 3360 305698 3369
rect 305642 3295 305698 3304
rect 306748 2440 306800 2446
rect 306748 2382 306800 2388
rect 306760 480 306788 2382
rect 309060 480 309088 3606
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 312556 6458 312584 21218
rect 313292 9246 313320 23310
rect 314672 20738 314700 23324
rect 315304 21752 315356 21758
rect 315304 21694 315356 21700
rect 314660 20732 314712 20738
rect 314660 20674 314712 20680
rect 315316 12034 315344 21694
rect 315684 20262 315712 23324
rect 316696 21350 316724 23324
rect 317524 23310 317722 23338
rect 316684 21344 316736 21350
rect 316684 21286 316736 21292
rect 317052 20800 317104 20806
rect 317052 20742 317104 20748
rect 315672 20256 315724 20262
rect 315672 20198 315724 20204
rect 317064 17610 317092 20742
rect 317052 17604 317104 17610
rect 317052 17546 317104 17552
rect 315304 12028 315356 12034
rect 315304 11970 315356 11976
rect 316040 10396 316092 10402
rect 316040 10338 316092 10344
rect 316684 10396 316736 10402
rect 316684 10338 316736 10344
rect 313280 9240 313332 9246
rect 313280 9182 313332 9188
rect 312544 6452 312596 6458
rect 312544 6394 312596 6400
rect 312636 3732 312688 3738
rect 312636 3674 312688 3680
rect 312648 480 312676 3674
rect 316052 3398 316080 10338
rect 316224 3800 316276 3806
rect 316224 3742 316276 3748
rect 316040 3392 316092 3398
rect 313830 3360 313886 3369
rect 316040 3334 316092 3340
rect 313830 3295 313886 3304
rect 313844 480 313872 3295
rect 316236 480 316264 3742
rect 316696 3466 316724 10338
rect 317524 10334 317552 23310
rect 318720 21214 318748 23324
rect 319732 21282 319760 23324
rect 320272 22364 320324 22370
rect 320272 22306 320324 22312
rect 319720 21276 319772 21282
rect 319720 21218 319772 21224
rect 318708 21208 318760 21214
rect 318708 21150 318760 21156
rect 318064 20732 318116 20738
rect 318064 20674 318116 20680
rect 318076 13394 318104 20674
rect 319444 20120 319496 20126
rect 319444 20062 319496 20068
rect 318064 13388 318116 13394
rect 318064 13330 318116 13336
rect 317512 10328 317564 10334
rect 317512 10270 317564 10276
rect 319456 3534 319484 20062
rect 320284 16574 320312 22306
rect 320744 20738 320772 23324
rect 321664 23310 321770 23338
rect 320824 21548 320876 21554
rect 320824 21490 320876 21496
rect 320732 20732 320784 20738
rect 320732 20674 320784 20680
rect 320284 16546 320496 16574
rect 319720 3936 319772 3942
rect 319720 3878 319772 3884
rect 319444 3528 319496 3534
rect 319444 3470 319496 3476
rect 316684 3460 316736 3466
rect 316684 3402 316736 3408
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 319732 480 319760 3878
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320836 7954 320864 21490
rect 320824 7948 320876 7954
rect 320824 7890 320876 7896
rect 321664 5098 321692 23310
rect 322768 21758 322796 23324
rect 322756 21752 322808 21758
rect 322756 21694 322808 21700
rect 323584 21684 323636 21690
rect 323584 21626 323636 21632
rect 322756 21208 322808 21214
rect 322756 21150 322808 21156
rect 322768 20330 322796 21150
rect 322756 20324 322808 20330
rect 322756 20266 322808 20272
rect 323596 18902 323624 21626
rect 323780 20806 323808 23324
rect 324332 23310 324806 23338
rect 323768 20800 323820 20806
rect 323768 20742 323820 20748
rect 323584 18896 323636 18902
rect 323584 18838 323636 18844
rect 324332 7886 324360 23310
rect 325700 21344 325752 21350
rect 325700 21286 325752 21292
rect 324320 7880 324372 7886
rect 324320 7822 324372 7828
rect 323584 7812 323636 7818
rect 323584 7754 323636 7760
rect 321652 5092 321704 5098
rect 321652 5034 321704 5040
rect 323596 3602 323624 7754
rect 325712 6914 325740 21286
rect 325804 21214 325832 23324
rect 325896 23310 326830 23338
rect 327092 23310 327842 23338
rect 328472 23310 328854 23338
rect 329866 23310 329972 23338
rect 325792 21208 325844 21214
rect 325792 21150 325844 21156
rect 325896 10538 325924 23310
rect 325884 10532 325936 10538
rect 325884 10474 325936 10480
rect 325712 6886 326384 6914
rect 323584 3596 323636 3602
rect 323584 3538 323636 3544
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 323320 480 323348 3470
rect 324412 2372 324464 2378
rect 324412 2314 324464 2320
rect 324424 480 324452 2314
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 327092 6526 327120 23310
rect 328472 9382 328500 23310
rect 329102 17368 329158 17377
rect 329102 17303 329158 17312
rect 328460 9376 328512 9382
rect 328460 9318 328512 9324
rect 327080 6520 327132 6526
rect 327080 6462 327132 6468
rect 329116 3466 329144 17303
rect 329944 16250 329972 23310
rect 330496 23310 330878 23338
rect 330496 22094 330524 23310
rect 330404 22066 330524 22094
rect 329932 16244 329984 16250
rect 329932 16186 329984 16192
rect 330404 14822 330432 22066
rect 331876 20398 331904 23324
rect 332704 23310 332902 23338
rect 333624 23310 333914 23338
rect 331864 20392 331916 20398
rect 331864 20334 331916 20340
rect 330484 20188 330536 20194
rect 330484 20130 330536 20136
rect 330392 14816 330444 14822
rect 330392 14758 330444 14764
rect 329656 9172 329708 9178
rect 329656 9114 329708 9120
rect 329668 3874 329696 9114
rect 329656 3868 329708 3874
rect 329656 3810 329708 3816
rect 330496 3738 330524 20130
rect 332600 19916 332652 19922
rect 332600 19858 332652 19864
rect 331220 11892 331272 11898
rect 331220 11834 331272 11840
rect 330576 10464 330628 10470
rect 330576 10406 330628 10412
rect 330484 3732 330536 3738
rect 330484 3674 330536 3680
rect 330588 3670 330616 10406
rect 330576 3664 330628 3670
rect 330576 3606 330628 3612
rect 330392 3596 330444 3602
rect 330392 3538 330444 3544
rect 329104 3460 329156 3466
rect 329104 3402 329156 3408
rect 328000 2304 328052 2310
rect 328000 2246 328052 2252
rect 328012 480 328040 2246
rect 330404 480 330432 3538
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 11834
rect 332612 9110 332640 19858
rect 332704 10606 332732 23310
rect 333624 19922 333652 23310
rect 333980 21548 334032 21554
rect 333980 21490 334032 21496
rect 333992 20058 334020 21490
rect 334912 21418 334940 23324
rect 335372 23310 335938 23338
rect 334900 21412 334952 21418
rect 334900 21354 334952 21360
rect 334624 20256 334676 20262
rect 334624 20198 334676 20204
rect 333980 20052 334032 20058
rect 333980 19994 334032 20000
rect 333612 19916 333664 19922
rect 333612 19858 333664 19864
rect 334636 16574 334664 20198
rect 334636 16546 334756 16574
rect 334624 11824 334676 11830
rect 334624 11766 334676 11772
rect 332692 10600 332744 10606
rect 332692 10542 332744 10548
rect 332600 9104 332652 9110
rect 332600 9046 332652 9052
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 333900 480 333928 3946
rect 333980 2848 334032 2854
rect 333980 2790 334032 2796
rect 333992 1358 334020 2790
rect 333980 1352 334032 1358
rect 333980 1294 334032 1300
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 11766
rect 334728 3534 334756 16546
rect 335372 10402 335400 23310
rect 335360 10396 335412 10402
rect 335360 10338 335412 10344
rect 336016 3738 336044 23666
rect 480260 23656 480312 23662
rect 480260 23598 480312 23604
rect 336844 23310 336950 23338
rect 337672 23310 337962 23338
rect 336740 19916 336792 19922
rect 336740 19858 336792 19864
rect 336752 10674 336780 19858
rect 336844 12102 336872 23310
rect 337672 19922 337700 23310
rect 338960 21622 338988 23324
rect 338948 21616 339000 21622
rect 338948 21558 339000 21564
rect 339972 20126 340000 23324
rect 340984 21554 341012 23324
rect 341076 23310 342010 23338
rect 340972 21548 341024 21554
rect 340972 21490 341024 21496
rect 339960 20120 340012 20126
rect 339960 20062 340012 20068
rect 337660 19916 337712 19922
rect 337660 19858 337712 19864
rect 337384 13320 337436 13326
rect 337384 13262 337436 13268
rect 336832 12096 336884 12102
rect 336832 12038 336884 12044
rect 336740 10668 336792 10674
rect 336740 10610 336792 10616
rect 336096 10328 336148 10334
rect 336096 10270 336148 10276
rect 336108 3806 336136 10270
rect 336096 3800 336148 3806
rect 336096 3742 336148 3748
rect 336004 3732 336056 3738
rect 336004 3674 336056 3680
rect 337396 3670 337424 13262
rect 340972 11960 341024 11966
rect 340972 11902 341024 11908
rect 337476 11824 337528 11830
rect 337476 11766 337528 11772
rect 337488 4010 337516 11766
rect 338672 11756 338724 11762
rect 338672 11698 338724 11704
rect 338764 11756 338816 11762
rect 338764 11698 338816 11704
rect 337568 10396 337620 10402
rect 337568 10338 337620 10344
rect 337476 4004 337528 4010
rect 337476 3946 337528 3952
rect 337580 3942 337608 10338
rect 337568 3936 337620 3942
rect 337568 3878 337620 3884
rect 337384 3664 337436 3670
rect 337384 3606 337436 3612
rect 334716 3528 334768 3534
rect 334716 3470 334768 3476
rect 337476 3052 337528 3058
rect 337476 2994 337528 3000
rect 337488 480 337516 2994
rect 338684 480 338712 11698
rect 338776 3602 338804 11698
rect 338764 3596 338816 3602
rect 338764 3538 338816 3544
rect 340984 3534 341012 11902
rect 341076 7818 341104 23310
rect 343008 21690 343036 23324
rect 343744 23310 344034 23338
rect 342996 21684 343048 21690
rect 342996 21626 343048 21632
rect 342904 21616 342956 21622
rect 342904 21558 342956 21564
rect 341064 7812 341116 7818
rect 341064 7754 341116 7760
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 340972 2984 341024 2990
rect 340972 2926 341024 2932
rect 340984 480 341012 2926
rect 342180 480 342208 3470
rect 342916 3058 342944 21558
rect 343640 21548 343692 21554
rect 343640 21490 343692 21496
rect 343652 6914 343680 21490
rect 343744 9178 343772 23310
rect 345032 21486 345060 23324
rect 345124 23310 346058 23338
rect 345020 21480 345072 21486
rect 345020 21422 345072 21428
rect 345124 10470 345152 23310
rect 347056 20194 347084 23324
rect 347884 23310 348082 23338
rect 348344 23310 349094 23338
rect 347780 21004 347832 21010
rect 347780 20946 347832 20952
rect 347044 20188 347096 20194
rect 347044 20130 347096 20136
rect 347044 14680 347096 14686
rect 347044 14622 347096 14628
rect 345112 10464 345164 10470
rect 345112 10406 345164 10412
rect 345664 10464 345716 10470
rect 345664 10406 345716 10412
rect 345294 10296 345350 10305
rect 345294 10231 345350 10240
rect 343732 9172 343784 9178
rect 343732 9114 343784 9120
rect 343652 6886 344600 6914
rect 342904 3052 342956 3058
rect 342904 2994 342956 3000
rect 344572 480 344600 6886
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 10231
rect 345676 2990 345704 10406
rect 347056 3534 347084 14622
rect 347792 6914 347820 20946
rect 347884 10334 347912 23310
rect 348344 10402 348372 23310
rect 349252 22296 349304 22302
rect 349252 22238 349304 22244
rect 348332 10396 348384 10402
rect 348332 10338 348384 10344
rect 347872 10328 347924 10334
rect 347872 10270 347924 10276
rect 348516 7744 348568 7750
rect 348516 7686 348568 7692
rect 347792 6886 348096 6914
rect 347044 3528 347096 3534
rect 347044 3470 347096 3476
rect 345664 2984 345716 2990
rect 345664 2926 345716 2932
rect 348068 480 348096 6886
rect 348528 3602 348556 7686
rect 348516 3596 348568 3602
rect 348516 3538 348568 3544
rect 349264 480 349292 22238
rect 350092 20262 350120 23324
rect 350632 21752 350684 21758
rect 350632 21694 350684 21700
rect 350080 20256 350132 20262
rect 350080 20198 350132 20204
rect 350644 16574 350672 21694
rect 351104 21418 351132 23324
rect 351932 23310 352130 23338
rect 352208 23310 353142 23338
rect 351092 21412 351144 21418
rect 351092 21354 351144 21360
rect 350644 16546 351224 16574
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 351932 11762 351960 23310
rect 352208 11830 352236 23310
rect 354140 21622 354168 23324
rect 354692 23310 355166 23338
rect 354128 21616 354180 21622
rect 354128 21558 354180 21564
rect 352196 11824 352248 11830
rect 352196 11766 352248 11772
rect 351920 11756 351972 11762
rect 351920 11698 351972 11704
rect 354692 10470 354720 23310
rect 356164 21554 356192 23324
rect 356152 21548 356204 21554
rect 356152 21490 356204 21496
rect 357176 21010 357204 23324
rect 358188 21758 358216 23324
rect 358176 21752 358228 21758
rect 358176 21694 358228 21700
rect 357164 21004 357216 21010
rect 357164 20946 357216 20952
rect 359200 20738 359228 23324
rect 360212 20738 360240 23324
rect 361238 23310 361528 23338
rect 361500 20754 361528 23310
rect 356704 20732 356756 20738
rect 356704 20674 356756 20680
rect 359188 20732 359240 20738
rect 359188 20674 359240 20680
rect 359464 20732 359516 20738
rect 359464 20674 359516 20680
rect 360200 20732 360252 20738
rect 361500 20726 361620 20754
rect 362236 20738 362264 23324
rect 363248 21010 363276 23324
rect 363524 23310 364274 23338
rect 363236 21004 363288 21010
rect 363236 20946 363288 20952
rect 360200 20674 360252 20680
rect 356336 13456 356388 13462
rect 356336 13398 356388 13404
rect 354680 10464 354732 10470
rect 354680 10406 354732 10412
rect 352840 3664 352892 3670
rect 352840 3606 352892 3612
rect 352852 480 352880 3606
rect 355232 3392 355284 3398
rect 355232 3334 355284 3340
rect 355244 480 355272 3334
rect 356348 480 356376 13398
rect 356716 3398 356744 20674
rect 359372 13252 359424 13258
rect 359372 13194 359424 13200
rect 356704 3392 356756 3398
rect 356704 3334 356756 3340
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359384 354 359412 13194
rect 359476 3398 359504 20674
rect 361592 16574 361620 20726
rect 362224 20732 362276 20738
rect 362224 20674 362276 20680
rect 361592 16546 361896 16574
rect 359464 3392 359516 3398
rect 359464 3334 359516 3340
rect 359894 354 360006 480
rect 359384 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363420 13184 363472 13190
rect 363420 13126 363472 13132
rect 363432 6914 363460 13126
rect 363524 11762 363552 23310
rect 365272 20738 365300 23324
rect 366284 20806 366312 23324
rect 366364 21004 366416 21010
rect 366364 20946 366416 20952
rect 366272 20800 366324 20806
rect 366272 20742 366324 20748
rect 363604 20732 363656 20738
rect 363604 20674 363656 20680
rect 365260 20732 365312 20738
rect 365260 20674 365312 20680
rect 363512 11756 363564 11762
rect 363512 11698 363564 11704
rect 363432 6886 363552 6914
rect 363524 480 363552 6886
rect 363616 3194 363644 20674
rect 365812 13116 365864 13122
rect 365812 13058 365864 13064
rect 365824 3398 365852 13058
rect 365812 3392 365864 3398
rect 365812 3334 365864 3340
rect 363604 3188 363656 3194
rect 363604 3130 363656 3136
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 365824 480 365852 3130
rect 366376 3126 366404 20946
rect 366456 20732 366508 20738
rect 366456 20674 366508 20680
rect 366468 13122 366496 20674
rect 367296 20058 367324 23324
rect 368308 21418 368336 23324
rect 369320 21690 369348 23324
rect 369872 23310 370346 23338
rect 369308 21684 369360 21690
rect 369308 21626 369360 21632
rect 368296 21412 368348 21418
rect 368296 21354 368348 21360
rect 367744 20800 367796 20806
rect 367744 20742 367796 20748
rect 367284 20052 367336 20058
rect 367284 19994 367336 20000
rect 366456 13116 366508 13122
rect 366456 13058 366508 13064
rect 367756 10470 367784 20742
rect 369872 13190 369900 23310
rect 371148 21684 371200 21690
rect 371148 21626 371200 21632
rect 371160 20126 371188 21626
rect 371344 21554 371372 23324
rect 371528 23310 372370 23338
rect 372724 23310 373382 23338
rect 374012 23310 374394 23338
rect 371332 21548 371384 21554
rect 371332 21490 371384 21496
rect 371148 20120 371200 20126
rect 371148 20062 371200 20068
rect 370504 14612 370556 14618
rect 370504 14554 370556 14560
rect 369860 13184 369912 13190
rect 369860 13126 369912 13132
rect 367744 10464 367796 10470
rect 367744 10406 367796 10412
rect 370516 3670 370544 14554
rect 371528 10334 371556 23310
rect 372724 11830 372752 23310
rect 372712 11824 372764 11830
rect 372712 11766 372764 11772
rect 374012 11762 374040 23310
rect 375392 21078 375420 23324
rect 375484 23310 376418 23338
rect 376772 23310 377430 23338
rect 375380 21072 375432 21078
rect 375380 21014 375432 21020
rect 375484 13258 375512 23310
rect 376772 14618 376800 23310
rect 377496 21548 377548 21554
rect 377496 21490 377548 21496
rect 376760 14612 376812 14618
rect 376760 14554 376812 14560
rect 377404 14544 377456 14550
rect 377404 14486 377456 14492
rect 375472 13252 375524 13258
rect 375472 13194 375524 13200
rect 376024 13116 376076 13122
rect 376024 13058 376076 13064
rect 372896 11756 372948 11762
rect 372896 11698 372948 11704
rect 374000 11756 374052 11762
rect 374000 11698 374052 11704
rect 371516 10328 371568 10334
rect 371516 10270 371568 10276
rect 370596 4956 370648 4962
rect 370596 4898 370648 4904
rect 370504 3664 370556 3670
rect 370504 3606 370556 3612
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 366364 3120 366416 3126
rect 366364 3062 366416 3068
rect 367020 480 367048 3334
rect 369400 3120 369452 3126
rect 369400 3062 369452 3068
rect 369412 480 369440 3062
rect 370608 480 370636 4898
rect 372908 480 372936 11698
rect 374092 3596 374144 3602
rect 374092 3538 374144 3544
rect 374104 480 374132 3538
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 13058
rect 377416 3398 377444 14486
rect 377508 10402 377536 21490
rect 378428 20738 378456 23324
rect 378704 23310 379454 23338
rect 378416 20732 378468 20738
rect 378416 20674 378468 20680
rect 378704 13394 378732 23310
rect 378784 21412 378836 21418
rect 378784 21354 378836 21360
rect 378796 20194 378824 21354
rect 380452 20874 380480 23324
rect 381464 21554 381492 23324
rect 382384 23310 382490 23338
rect 381452 21548 381504 21554
rect 381452 21490 381504 21496
rect 381726 21312 381782 21321
rect 381726 21247 381782 21256
rect 380440 20868 380492 20874
rect 380440 20810 380492 20816
rect 380164 20732 380216 20738
rect 380164 20674 380216 20680
rect 378784 20188 378836 20194
rect 378784 20130 378836 20136
rect 380176 14822 380204 20674
rect 380164 14816 380216 14822
rect 380164 14758 380216 14764
rect 381544 14476 381596 14482
rect 381544 14418 381596 14424
rect 378692 13388 378744 13394
rect 378692 13330 378744 13336
rect 379520 10464 379572 10470
rect 379520 10406 379572 10412
rect 377496 10396 377548 10402
rect 377496 10338 377548 10344
rect 377680 3528 377732 3534
rect 377680 3470 377732 3476
rect 377404 3392 377456 3398
rect 377404 3334 377456 3340
rect 377692 480 377720 3470
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 10406
rect 381556 3670 381584 14418
rect 381740 13326 381768 21247
rect 382280 20052 382332 20058
rect 382280 19994 382332 20000
rect 381728 13320 381780 13326
rect 381728 13262 381780 13268
rect 381636 13184 381688 13190
rect 381636 13126 381688 13132
rect 381176 3664 381228 3670
rect 381176 3606 381228 3612
rect 381544 3664 381596 3670
rect 381544 3606 381596 3612
rect 381188 480 381216 3606
rect 381648 3602 381676 13126
rect 381636 3596 381688 3602
rect 381636 3538 381688 3544
rect 382292 3534 382320 19994
rect 382384 10606 382412 23310
rect 383488 21826 383516 23324
rect 383476 21820 383528 21826
rect 383476 21762 383528 21768
rect 382924 21072 382976 21078
rect 382924 21014 382976 21020
rect 382936 20058 382964 21014
rect 384396 20868 384448 20874
rect 384396 20810 384448 20816
rect 382924 20052 382976 20058
rect 382924 19994 382976 20000
rect 384408 14754 384436 20810
rect 384500 20738 384528 23324
rect 385512 21758 385540 23324
rect 385500 21752 385552 21758
rect 385500 21694 385552 21700
rect 386524 21690 386552 23324
rect 386708 23310 387550 23338
rect 386512 21684 386564 21690
rect 386512 21626 386564 21632
rect 384488 20732 384540 20738
rect 384488 20674 384540 20680
rect 386420 20188 386472 20194
rect 386420 20130 386472 20136
rect 384396 14748 384448 14754
rect 384396 14690 384448 14696
rect 384302 14512 384358 14521
rect 384302 14447 384358 14456
rect 382372 10600 382424 10606
rect 382372 10542 382424 10548
rect 384316 3534 384344 14447
rect 386432 6914 386460 20130
rect 386708 13190 386736 23310
rect 388444 21820 388496 21826
rect 388444 21762 388496 21768
rect 387064 21548 387116 21554
rect 387064 21490 387116 21496
rect 386696 13184 386748 13190
rect 386696 13126 386748 13132
rect 387076 12034 387104 21490
rect 388456 14686 388484 21762
rect 388548 21622 388576 23324
rect 388536 21616 388588 21622
rect 388536 21558 388588 21564
rect 389560 19582 389588 23324
rect 390572 21486 390600 23324
rect 390664 23310 391598 23338
rect 390560 21480 390612 21486
rect 390560 21422 390612 21428
rect 389548 19576 389600 19582
rect 389548 19518 389600 19524
rect 390664 16574 390692 23310
rect 392596 21554 392624 23324
rect 393332 23310 393622 23338
rect 394528 23310 394634 23338
rect 394804 23310 395646 23338
rect 392584 21548 392636 21554
rect 392584 21490 392636 21496
rect 392584 20732 392636 20738
rect 392584 20674 392636 20680
rect 390744 20120 390796 20126
rect 390744 20062 390796 20068
rect 390572 16546 390692 16574
rect 388444 14680 388496 14686
rect 388444 14622 388496 14628
rect 387064 12028 387116 12034
rect 387064 11970 387116 11976
rect 386432 6886 386736 6914
rect 382280 3528 382332 3534
rect 382280 3470 382332 3476
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 384304 3528 384356 3534
rect 384304 3470 384356 3476
rect 383580 480 383608 3470
rect 384764 3392 384816 3398
rect 384764 3334 384816 3340
rect 384776 480 384804 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 6886
rect 390572 3670 390600 16546
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 390560 3664 390612 3670
rect 390560 3606 390612 3612
rect 388272 480 388300 3606
rect 390284 3596 390336 3602
rect 390284 3538 390336 3544
rect 390296 3398 390324 3538
rect 390284 3392 390336 3398
rect 390284 3334 390336 3340
rect 390756 2774 390784 20062
rect 392596 7818 392624 20674
rect 393332 11014 393360 23310
rect 394528 21418 394556 23310
rect 394700 22228 394752 22234
rect 394700 22170 394752 22176
rect 394608 21752 394660 21758
rect 394608 21694 394660 21700
rect 394516 21412 394568 21418
rect 394516 21354 394568 21360
rect 394620 20262 394648 21694
rect 394608 20256 394660 20262
rect 394608 20198 394660 20204
rect 393964 19576 394016 19582
rect 393964 19518 394016 19524
rect 393320 11008 393372 11014
rect 393320 10950 393372 10956
rect 392584 7812 392636 7818
rect 392584 7754 392636 7760
rect 393976 3670 394004 19518
rect 393964 3664 394016 3670
rect 393964 3606 394016 3612
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390664 2746 390784 2774
rect 390664 480 390692 2746
rect 391860 480 391888 3470
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 394252 480 394280 3334
rect 394712 2774 394740 22170
rect 394804 9178 394832 23310
rect 396644 20194 396672 23324
rect 396632 20188 396684 20194
rect 396632 20130 396684 20136
rect 397656 20126 397684 23324
rect 398668 21758 398696 23324
rect 398852 23310 399694 23338
rect 400232 23310 400706 23338
rect 398656 21752 398708 21758
rect 398656 21694 398708 21700
rect 397644 20120 397696 20126
rect 397644 20062 397696 20068
rect 398852 10538 398880 23310
rect 398930 11656 398986 11665
rect 398930 11591 398986 11600
rect 398840 10532 398892 10538
rect 398840 10474 398892 10480
rect 397736 10396 397788 10402
rect 397736 10338 397788 10344
rect 394792 9172 394844 9178
rect 394792 9114 394844 9120
rect 394712 2746 395384 2774
rect 395356 480 395384 2746
rect 397748 480 397776 10338
rect 398944 480 398972 11591
rect 399484 11008 399536 11014
rect 399484 10950 399536 10956
rect 399496 3602 399524 10950
rect 400232 10470 400260 23310
rect 401600 19916 401652 19922
rect 401600 19858 401652 19864
rect 400220 10464 400272 10470
rect 400220 10406 400272 10412
rect 401612 10402 401640 19858
rect 401704 16250 401732 23324
rect 402440 23310 402730 23338
rect 402992 23310 403742 23338
rect 404372 23310 404754 23338
rect 405766 23310 405872 23338
rect 402440 19922 402468 23310
rect 402428 19916 402480 19922
rect 402428 19858 402480 19864
rect 401692 16244 401744 16250
rect 401692 16186 401744 16192
rect 402992 16182 403020 23310
rect 402980 16176 403032 16182
rect 402980 16118 403032 16124
rect 401600 10396 401652 10402
rect 401600 10338 401652 10344
rect 400864 10328 400916 10334
rect 400864 10270 400916 10276
rect 399484 3596 399536 3602
rect 399484 3538 399536 3544
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 10270
rect 404372 9110 404400 23310
rect 405844 11966 405872 23310
rect 405936 23310 406778 23338
rect 407224 23310 407790 23338
rect 408696 23310 408802 23338
rect 409432 23310 409814 23338
rect 409892 23310 410826 23338
rect 405832 11960 405884 11966
rect 405832 11902 405884 11908
rect 405936 11898 405964 23310
rect 406016 16108 406068 16114
rect 406016 16050 406068 16056
rect 405924 11892 405976 11898
rect 405924 11834 405976 11840
rect 404452 11824 404504 11830
rect 404452 11766 404504 11772
rect 404360 9104 404412 9110
rect 404360 9046 404412 9052
rect 402520 3732 402572 3738
rect 402520 3674 402572 3680
rect 402532 480 402560 3674
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404464 354 404492 11766
rect 406028 480 406056 16050
rect 407224 11830 407252 23310
rect 408592 19916 408644 19922
rect 408592 19858 408644 19864
rect 407212 11824 407264 11830
rect 407212 11766 407264 11772
rect 408604 11762 408632 19858
rect 408696 16046 408724 23310
rect 409432 19922 409460 23310
rect 409420 19916 409472 19922
rect 409420 19858 409472 19864
rect 409144 16108 409196 16114
rect 409144 16050 409196 16056
rect 408684 16040 408736 16046
rect 408684 15982 408736 15988
rect 407120 11756 407172 11762
rect 407120 11698 407172 11704
rect 408592 11756 408644 11762
rect 408592 11698 408644 11704
rect 407132 3398 407160 11698
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404464 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16050
rect 409892 10334 409920 23310
rect 411824 20058 411852 23324
rect 411260 20052 411312 20058
rect 411260 19994 411312 20000
rect 411812 20052 411864 20058
rect 411812 19994 411864 20000
rect 411272 16574 411300 19994
rect 412732 19916 412784 19922
rect 412732 19858 412784 19864
rect 411272 16546 411944 16574
rect 409880 10328 409932 10334
rect 409880 10270 409932 10276
rect 411916 480 411944 16546
rect 412640 15972 412692 15978
rect 412640 15914 412692 15920
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 15914
rect 412744 13258 412772 19858
rect 412836 15978 412864 23324
rect 413480 23310 413862 23338
rect 414032 23310 414874 23338
rect 415596 23310 415886 23338
rect 413480 19922 413508 23310
rect 413468 19916 413520 19922
rect 413468 19858 413520 19864
rect 412824 15972 412876 15978
rect 412824 15914 412876 15920
rect 412732 13252 412784 13258
rect 412732 13194 412784 13200
rect 414032 13190 414060 23310
rect 415400 15904 415452 15910
rect 415400 15846 415452 15852
rect 413284 13184 413336 13190
rect 413284 13126 413336 13132
rect 414020 13184 414072 13190
rect 414020 13126 414072 13132
rect 413296 3738 413324 13126
rect 413284 3732 413336 3738
rect 413284 3674 413336 3680
rect 415412 2786 415440 15846
rect 415596 13122 415624 23310
rect 416884 17474 416912 23324
rect 417068 23310 417910 23338
rect 418172 23310 418922 23338
rect 419552 23310 419934 23338
rect 420946 23310 421052 23338
rect 416872 17468 416924 17474
rect 416872 17410 416924 17416
rect 415492 13116 415544 13122
rect 415492 13058 415544 13064
rect 415584 13116 415636 13122
rect 415584 13058 415636 13064
rect 415400 2780 415452 2786
rect 415400 2722 415452 2728
rect 415504 480 415532 13058
rect 417068 7750 417096 23310
rect 417056 7744 417108 7750
rect 417056 7686 417108 7692
rect 418172 4962 418200 23310
rect 419552 14618 419580 23310
rect 420920 18964 420972 18970
rect 420920 18906 420972 18912
rect 418528 14612 418580 14618
rect 418528 14554 418580 14560
rect 419540 14612 419592 14618
rect 419540 14554 419592 14560
rect 418160 4956 418212 4962
rect 418160 4898 418212 4904
rect 416688 2780 416740 2786
rect 416688 2722 416740 2728
rect 416700 480 416728 2722
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 354 418568 14554
rect 420932 14482 420960 18906
rect 421024 14550 421052 23310
rect 421576 23310 421958 23338
rect 422312 23310 422970 23338
rect 421576 18970 421604 23310
rect 421564 18964 421616 18970
rect 421564 18906 421616 18912
rect 421012 14544 421064 14550
rect 421012 14486 421064 14492
rect 420920 14476 420972 14482
rect 420920 14418 420972 14424
rect 420182 9072 420238 9081
rect 420182 9007 420238 9016
rect 420196 480 420224 9007
rect 422312 6390 422340 23310
rect 437572 21752 437624 21758
rect 437572 21694 437624 21700
rect 426808 21684 426860 21690
rect 426808 21626 426860 21632
rect 426820 17542 426848 21626
rect 426440 17536 426492 17542
rect 426440 17478 426492 17484
rect 426808 17536 426860 17542
rect 426808 17478 426860 17484
rect 426452 16574 426480 17478
rect 430580 17400 430632 17406
rect 430580 17342 430632 17348
rect 430592 16574 430620 17342
rect 433340 17332 433392 17338
rect 433340 17274 433392 17280
rect 433352 16574 433380 17274
rect 437584 17270 437612 21694
rect 440240 21616 440292 21622
rect 440240 21558 440292 21564
rect 440252 17338 440280 21558
rect 456892 21548 456944 21554
rect 456892 21490 456944 21496
rect 447140 20256 447192 20262
rect 447140 20198 447192 20204
rect 440240 17332 440292 17338
rect 440240 17274 440292 17280
rect 437480 17264 437532 17270
rect 437480 17206 437532 17212
rect 437572 17264 437624 17270
rect 437572 17206 437624 17212
rect 440238 17232 440294 17241
rect 426452 16546 426848 16574
rect 430592 16546 430896 16574
rect 433352 16546 434024 16574
rect 422576 14816 422628 14822
rect 422576 14758 422628 14764
rect 422300 6384 422352 6390
rect 422300 6326 422352 6332
rect 422588 480 422616 14758
rect 425704 13388 425756 13394
rect 425704 13330 425756 13336
rect 423772 2236 423824 2242
rect 423772 2178 423824 2184
rect 423784 480 423812 2178
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 13330
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 429200 14748 429252 14754
rect 429200 14690 429252 14696
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 14690
rect 430868 480 430896 16546
rect 431960 12028 432012 12034
rect 431960 11970 432012 11976
rect 431972 3398 432000 11970
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 436744 10600 436796 10606
rect 436744 10542 436796 10548
rect 436756 480 436784 10542
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 17206
rect 440238 17167 440294 17176
rect 440252 1970 440280 17167
rect 447152 16574 447180 20198
rect 451280 18828 451332 18834
rect 451280 18770 451332 18776
rect 449900 17536 449952 17542
rect 449900 17478 449952 17484
rect 449912 16574 449940 17478
rect 451292 16574 451320 18770
rect 455420 18760 455472 18766
rect 455420 18702 455472 18708
rect 455432 16574 455460 18702
rect 456904 17338 456932 21490
rect 465080 21480 465132 21486
rect 465080 21422 465132 21428
rect 458180 18692 458232 18698
rect 458180 18634 458232 18640
rect 456800 17332 456852 17338
rect 456800 17274 456852 17280
rect 456892 17332 456944 17338
rect 456892 17274 456944 17280
rect 447152 16546 447456 16574
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 455432 16546 455736 16574
rect 440332 14680 440384 14686
rect 440332 14622 440384 14628
rect 440240 1964 440292 1970
rect 440240 1906 440292 1912
rect 440344 480 440372 14622
rect 443828 7812 443880 7818
rect 443828 7754 443880 7760
rect 441528 1964 441580 1970
rect 441528 1906 441580 1912
rect 441540 480 441568 1906
rect 443840 480 443868 7754
rect 445022 6352 445078 6361
rect 445022 6287 445078 6296
rect 445036 480 445064 6287
rect 447428 480 447456 16546
rect 448610 15872 448666 15881
rect 448610 15807 448666 15816
rect 448624 480 448652 15807
rect 450924 480 450952 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 454500 3732 454552 3738
rect 454500 3674 454552 3680
rect 454512 480 454540 3674
rect 455708 480 455736 16546
rect 456812 3398 456840 17274
rect 458192 16574 458220 18634
rect 462320 18624 462372 18630
rect 462320 18566 462372 18572
rect 458192 16546 459232 16574
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 461584 3664 461636 3670
rect 461584 3606 461636 3612
rect 461596 480 461624 3606
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 18566
rect 465092 6914 465120 21422
rect 478880 21412 478932 21418
rect 478880 21354 478932 21360
rect 469220 19984 469272 19990
rect 469220 19926 469272 19932
rect 476118 19952 476174 19961
rect 465170 18592 465226 18601
rect 465170 18527 465226 18536
rect 465184 16574 465212 18527
rect 469232 16574 469260 19926
rect 476118 19887 476174 19896
rect 471980 17332 472032 17338
rect 471980 17274 472032 17280
rect 471992 16574 472020 17274
rect 476132 16574 476160 19887
rect 465184 16546 465856 16574
rect 469232 16546 469904 16574
rect 471992 16546 472296 16574
rect 476132 16546 476528 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 468760 6384 468812 6390
rect 468760 6326 468812 6332
rect 468772 3534 468800 6326
rect 468668 3528 468720 3534
rect 468668 3470 468720 3476
rect 468760 3528 468812 3534
rect 468760 3470 468812 3476
rect 468680 480 468708 3470
rect 469876 480 469904 16546
rect 472268 480 472296 16546
rect 475752 3596 475804 3602
rect 475752 3538 475804 3544
rect 473452 2168 473504 2174
rect 473452 2110 473504 2116
rect 473464 480 473492 2110
rect 475764 480 475792 3538
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 21354
rect 480272 16574 480300 23598
rect 483020 23588 483072 23594
rect 483020 23530 483072 23536
rect 483032 16574 483060 23530
rect 489920 23520 489972 23526
rect 489920 23462 489972 23468
rect 518898 23488 518954 23497
rect 485780 20188 485832 20194
rect 485780 20130 485832 20136
rect 485792 16574 485820 20130
rect 480272 16546 480576 16574
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 480258 7576 480314 7585
rect 480258 7511 480314 7520
rect 480272 3602 480300 7511
rect 480260 3596 480312 3602
rect 480260 3538 480312 3544
rect 480548 480 480576 16546
rect 482836 9172 482888 9178
rect 482836 9114 482888 9120
rect 482848 480 482876 9114
rect 484044 480 484072 16546
rect 486436 480 486464 16546
rect 487160 4888 487212 4894
rect 487160 4830 487212 4836
rect 487172 3670 487200 4830
rect 487160 3664 487212 3670
rect 487160 3606 487212 3612
rect 489932 3398 489960 23462
rect 518898 23423 518954 23432
rect 512000 22160 512052 22166
rect 512000 22102 512052 22108
rect 490012 20120 490064 20126
rect 490012 20062 490064 20068
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 3210 490052 20062
rect 492680 17264 492732 17270
rect 492680 17206 492732 17212
rect 492692 16574 492720 17206
rect 492692 16546 493088 16574
rect 490748 3392 490800 3398
rect 490748 3334 490800 3340
rect 489932 3182 490052 3210
rect 489932 480 489960 3182
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 218 487702 480
rect 487264 202 487702 218
rect 487252 196 487702 202
rect 487304 190 487702 196
rect 487252 138 487304 144
rect 487590 -960 487702 190
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3334
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 503720 16244 503772 16250
rect 503720 16186 503772 16192
rect 494796 11960 494848 11966
rect 494796 11902 494848 11908
rect 494808 3670 494836 11902
rect 497096 10532 497148 10538
rect 497096 10474 497148 10480
rect 494704 3664 494756 3670
rect 494704 3606 494756 3612
rect 494796 3664 494848 3670
rect 494796 3606 494848 3612
rect 494716 480 494744 3606
rect 497108 480 497136 10474
rect 500592 10464 500644 10470
rect 500592 10406 500644 10412
rect 498200 4820 498252 4826
rect 498200 4762 498252 4768
rect 498212 480 498240 4762
rect 500604 480 500632 10406
rect 501786 4992 501842 5001
rect 501786 4927 501842 4936
rect 501800 480 501828 4927
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 16186
rect 511264 16176 511316 16182
rect 511264 16118 511316 16124
rect 507216 10396 507268 10402
rect 507216 10338 507268 10344
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505560 128 505612 134
rect 505346 76 505560 82
rect 505346 70 505612 76
rect 505346 54 505600 70
rect 505346 -960 505458 54
rect 506450 -960 506562 480
rect 507228 354 507256 10338
rect 508872 2848 508924 2854
rect 508872 2790 508924 2796
rect 508884 480 508912 2790
rect 511276 480 511304 16118
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 22102
rect 518912 16574 518940 23423
rect 532698 22128 532754 22137
rect 532698 22063 532754 22072
rect 532712 16574 532740 22063
rect 539600 20052 539652 20058
rect 539600 19994 539652 20000
rect 518912 16546 519584 16574
rect 532712 16546 533752 16574
rect 515496 13320 515548 13326
rect 515496 13262 515548 13268
rect 514760 9104 514812 9110
rect 514760 9046 514812 9052
rect 514772 480 514800 9046
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515508 354 515536 13262
rect 518348 3664 518400 3670
rect 518348 3606 518400 3612
rect 518360 480 518388 3606
rect 519556 480 519584 16546
rect 528560 16040 528612 16046
rect 528560 15982 528612 15988
rect 521660 11892 521712 11898
rect 521660 11834 521712 11840
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521672 354 521700 11834
rect 525432 11824 525484 11830
rect 525432 11766 525484 11772
rect 523040 6316 523092 6322
rect 523040 6258 523092 6264
rect 523052 480 523080 6258
rect 525444 480 525472 11766
rect 526628 6248 526680 6254
rect 526628 6190 526680 6196
rect 526640 480 526668 6190
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 15982
rect 532056 11756 532108 11762
rect 532056 11698 532108 11704
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 82 530206 480
rect 529952 66 530206 82
rect 529940 60 530206 66
rect 529992 54 530206 60
rect 529940 2 529992 8
rect 530094 -960 530206 54
rect 531290 -960 531402 480
rect 532068 354 532096 11698
rect 533724 480 533752 16546
rect 536104 10328 536156 10334
rect 536104 10270 536156 10276
rect 536116 480 536144 10270
rect 537208 2100 537260 2106
rect 537208 2042 537260 2048
rect 537220 480 537248 2042
rect 539612 480 539640 19994
rect 556160 17468 556212 17474
rect 556160 17410 556212 17416
rect 556172 16574 556200 17410
rect 556172 16546 556936 16574
rect 542728 15972 542780 15978
rect 542728 15914 542780 15920
rect 540794 4856 540850 4865
rect 540794 4791 540850 4800
rect 540808 480 540836 4791
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 15914
rect 546500 13252 546552 13258
rect 546500 13194 546552 13200
rect 544384 6180 544436 6186
rect 544384 6122 544436 6128
rect 544396 480 544424 6122
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 13194
rect 550272 13184 550324 13190
rect 550272 13126 550324 13132
rect 547880 7676 547932 7682
rect 547880 7618 547932 7624
rect 547892 480 547920 7618
rect 550284 480 550312 13126
rect 553768 13116 553820 13122
rect 553768 13058 553820 13064
rect 551468 7608 551520 7614
rect 551468 7550 551520 7556
rect 551480 480 551508 7550
rect 553780 480 553808 13058
rect 555424 9036 555476 9042
rect 555424 8978 555476 8984
rect 555436 3602 555464 8978
rect 554964 3596 555016 3602
rect 554964 3538 555016 3544
rect 555424 3596 555476 3602
rect 555424 3538 555476 3544
rect 554976 480 555004 3538
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 560852 7744 560904 7750
rect 560852 7686 560904 7692
rect 558550 2000 558606 2009
rect 558550 1935 558606 1944
rect 558564 480 558592 1935
rect 560864 480 560892 7686
rect 564440 4956 564492 4962
rect 564440 4898 564492 4904
rect 562048 3460 562100 3466
rect 562048 3402 562100 3408
rect 562060 480 562088 3402
rect 564452 480 564480 4898
rect 565096 3466 565124 37266
rect 567568 14612 567620 14618
rect 567568 14554 567620 14560
rect 565634 6216 565690 6225
rect 565634 6151 565690 6160
rect 565084 3460 565136 3466
rect 565084 3402 565136 3408
rect 565648 480 565676 6151
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 14554
rect 571340 14544 571392 14550
rect 571340 14486 571392 14492
rect 569132 3596 569184 3602
rect 569132 3538 569184 3544
rect 569144 480 569172 3538
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 14486
rect 575112 14476 575164 14482
rect 575112 14418 575164 14424
rect 572718 8936 572774 8945
rect 572718 8871 572774 8880
rect 572732 480 572760 8871
rect 575124 480 575152 14418
rect 576308 8968 576360 8974
rect 576308 8910 576360 8916
rect 576320 480 576348 8910
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 19246 699760 19302 699816
rect 3514 671200 3570 671256
rect 2778 658144 2834 658200
rect 2778 606056 2834 606112
rect 3422 566888 3478 566944
rect 2778 553832 2834 553888
rect 2870 514820 2926 514856
rect 2870 514800 2872 514820
rect 2872 514800 2924 514820
rect 2924 514800 2926 514820
rect 2778 501744 2834 501800
rect 3330 462576 3386 462632
rect 2778 449520 2834 449576
rect 3146 410488 3202 410544
rect 2778 397432 2834 397488
rect 2962 358400 3018 358456
rect 3330 345364 3386 345400
rect 3330 345344 3332 345364
rect 3332 345344 3384 345364
rect 3384 345344 3386 345364
rect 3330 319232 3386 319288
rect 3330 267144 3386 267200
rect 2778 241032 2834 241088
rect 3330 214920 3386 214976
rect 3606 619112 3662 619168
rect 3514 332424 3570 332480
rect 3514 293120 3570 293176
rect 3422 204040 3478 204096
rect 2778 188808 2834 188864
rect 2962 149776 3018 149832
rect 2778 136740 2834 136776
rect 2778 136720 2780 136740
rect 2780 136720 2832 136740
rect 2832 136720 2834 136740
rect 3422 110608 3478 110664
rect 2778 84632 2834 84688
rect 3422 71576 3478 71632
rect 3514 45464 3570 45520
rect 3606 32408 3662 32464
rect 16394 460128 16450 460184
rect 17130 199144 17186 199200
rect 18786 458804 18788 458824
rect 18788 458804 18840 458824
rect 18840 458804 18842 458824
rect 18786 458768 18842 458804
rect 17406 185952 17462 186008
rect 17590 74432 17646 74488
rect 20350 571920 20406 571976
rect 20350 204176 20406 204232
rect 19338 203904 19394 203960
rect 397458 700304 397514 700360
rect 23202 585792 23258 585848
rect 22926 458904 22982 458960
rect 21638 331744 21694 331800
rect 20626 202816 20682 202872
rect 63590 585792 63646 585848
rect 83830 585656 83886 585712
rect 149978 585792 150034 585848
rect 134430 582936 134486 582992
rect 175186 580216 175242 580272
rect 109038 571920 109094 571976
rect 226154 585656 226210 585712
rect 210974 582936 211030 582992
rect 527270 699760 527326 699816
rect 527178 697448 527234 697504
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 287518 585656 287574 585712
rect 286414 585112 286470 585168
rect 276018 572056 276074 572112
rect 204258 571920 204314 571976
rect 39302 570560 39358 570616
rect 286230 461896 286286 461952
rect 24858 460264 24914 460320
rect 34518 458940 34520 458960
rect 34520 458940 34572 458960
rect 34572 458940 34574 458960
rect 34518 458904 34574 458940
rect 93950 458768 94006 458824
rect 124310 460264 124366 460320
rect 134430 460128 134486 460184
rect 83830 458088 83886 458144
rect 160006 460808 160062 460864
rect 24950 444216 25006 444272
rect 175186 460128 175242 460184
rect 211158 458088 211214 458144
rect 285310 460128 285366 460184
rect 281446 459448 281502 459504
rect 276754 459040 276810 459096
rect 285402 458224 285458 458280
rect 285402 443808 285458 443864
rect 204258 443672 204314 443728
rect 286322 460708 286324 460728
rect 286324 460708 286376 460728
rect 286376 460708 286378 460728
rect 286322 460672 286378 460708
rect 286874 458904 286930 458960
rect 287610 459584 287666 459640
rect 287702 459448 287758 459504
rect 288714 460264 288770 460320
rect 288714 459720 288770 459776
rect 286230 456864 286286 456920
rect 285770 333784 285826 333840
rect 286966 333784 287022 333840
rect 22650 331744 22706 331800
rect 28170 332424 28226 332480
rect 22006 315868 22008 315888
rect 22008 315868 22060 315888
rect 22060 315868 22062 315888
rect 22006 315832 22062 315868
rect 22006 204196 22062 204232
rect 22006 204176 22008 204196
rect 22008 204176 22060 204196
rect 22060 204176 22062 204196
rect 22190 204176 22246 204232
rect 22190 203904 22246 203960
rect 22742 202816 22798 202872
rect 23386 330964 23388 330984
rect 23388 330964 23440 330984
rect 23440 330964 23442 330984
rect 23386 330928 23442 330964
rect 68650 331744 68706 331800
rect 149610 331744 149666 331800
rect 160098 330384 160154 330440
rect 171782 315288 171838 315344
rect 241334 332424 241390 332480
rect 204258 315288 204314 315344
rect 285402 316648 285458 316704
rect 285678 332188 285680 332208
rect 285680 332188 285732 332208
rect 285732 332188 285734 332208
rect 285678 332152 285734 332188
rect 286874 333648 286930 333704
rect 286690 331200 286746 331256
rect 287610 457952 287666 458008
rect 286966 315424 287022 315480
rect 23846 205808 23902 205864
rect 23018 203904 23074 203960
rect 23202 203904 23258 203960
rect 22926 202716 22928 202736
rect 22928 202716 22980 202736
rect 22980 202716 22982 202736
rect 22926 202680 22982 202716
rect 23754 205672 23810 205728
rect 284942 205672 284998 205728
rect 28170 204040 28226 204096
rect 43350 203904 43406 203960
rect 94042 204176 94098 204232
rect 68650 202816 68706 202872
rect 24858 202136 24914 202192
rect 96618 202136 96674 202192
rect 24858 186360 24914 186416
rect 124218 185952 124274 186008
rect 271694 203496 271750 203552
rect 204258 188264 204314 188320
rect 285770 205808 285826 205864
rect 285678 203632 285734 203688
rect 286966 204856 287022 204912
rect 284942 185952 284998 186008
rect 286966 186088 287022 186144
rect 285126 185816 285182 185872
rect 25594 77832 25650 77888
rect 52458 77016 52514 77072
rect 53792 77016 53848 77072
rect 52458 75928 52514 75984
rect 84106 75656 84162 75712
rect 79414 75520 79470 75576
rect 98642 75792 98698 75848
rect 104162 74432 104218 74488
rect 129002 71712 129058 71768
rect 151726 76472 151782 76528
rect 151634 53080 151690 53136
rect 150438 50496 150494 50552
rect 150438 49544 150494 49600
rect 150438 48220 150440 48240
rect 150440 48220 150492 48240
rect 150492 48220 150494 48240
rect 150438 48184 150494 48220
rect 150530 47640 150586 47696
rect 150438 46688 150494 46744
rect 151082 45464 151138 45520
rect 150438 44784 150494 44840
rect 150438 43832 150494 43888
rect 150438 42472 150494 42528
rect 150438 41248 150494 41304
rect 151542 39888 151598 39944
rect 150438 35844 150440 35864
rect 150440 35844 150492 35864
rect 150492 35844 150494 35864
rect 150438 35808 150494 35844
rect 150438 34312 150494 34368
rect 150438 32408 150494 32464
rect 150438 31456 150494 31512
rect 150438 30096 150494 30152
rect 150438 28908 150440 28928
rect 150440 28908 150492 28928
rect 150492 28908 150494 28928
rect 150438 28872 150494 28908
rect 153014 40364 153070 40420
rect 194598 77832 194654 77888
rect 195794 77832 195850 77888
rect 198830 68176 198886 68232
rect 204350 73752 204406 73808
rect 202878 54440 202934 54496
rect 217230 59880 217286 59936
rect 215758 57432 215814 57488
rect 213918 57296 213974 57352
rect 224958 76608 225014 76664
rect 233238 75112 233294 75168
rect 284298 77696 284354 77752
rect 282182 76744 282238 76800
rect 276478 54576 276534 54632
rect 280158 54712 280214 54768
rect 282274 73888 282330 73944
rect 282182 54440 282238 54496
rect 283838 54440 283894 54496
rect 285770 53896 285826 53952
rect 287610 54848 287666 54904
rect 288622 334192 288678 334248
rect 290094 433880 290150 433936
rect 290094 334056 290150 334112
rect 291382 459720 291438 459776
rect 288622 177928 288678 177984
rect 289910 332424 289966 332480
rect 291474 305632 291530 305688
rect 291474 205944 291530 206000
rect 290002 203632 290058 203688
rect 298006 582936 298062 582992
rect 293222 331880 293278 331936
rect 294050 205672 294106 205728
rect 291474 185816 291530 185872
rect 291474 77696 291530 77752
rect 291474 76336 291530 76392
rect 295338 185952 295394 186008
rect 295338 77832 295394 77888
rect 297178 443944 297234 444000
rect 297914 442856 297970 442912
rect 297178 76880 297234 76936
rect 297914 204992 297970 205048
rect 299110 329704 299166 329760
rect 300490 458224 300546 458280
rect 300122 331744 300178 331800
rect 299202 201184 299258 201240
rect 301870 459468 301926 459504
rect 301870 459448 301872 459468
rect 301872 459448 301924 459468
rect 301924 459448 301926 459468
rect 303158 459040 303214 459096
rect 301502 203496 301558 203552
rect 369214 582936 369270 582992
rect 389454 580216 389510 580272
rect 404358 571920 404414 571976
rect 440054 580216 440110 580272
rect 450174 580352 450230 580408
rect 485594 585792 485650 585848
rect 480534 585656 480590 585712
rect 490654 582936 490710 582992
rect 505834 583072 505890 583128
rect 556434 585792 556490 585848
rect 551374 585656 551430 585712
rect 566554 585112 566610 585168
rect 434718 571920 434774 571976
rect 424322 570560 424378 570616
rect 303526 461896 303582 461952
rect 305090 461760 305146 461816
rect 302882 313928 302938 313984
rect 303066 307672 303122 307728
rect 313278 459040 313334 459096
rect 414018 443672 414074 443728
rect 455234 460128 455290 460184
rect 485594 458904 485650 458960
rect 480534 458768 480590 458824
rect 490654 458088 490710 458144
rect 556158 459584 556214 459640
rect 565726 460944 565782 461000
rect 564898 460264 564954 460320
rect 561494 459448 561550 459504
rect 564438 459040 564494 459096
rect 551374 458768 551430 458824
rect 424322 443536 424378 443592
rect 565910 458108 565966 458144
rect 565910 458088 565912 458108
rect 565912 458088 565964 458108
rect 565964 458088 565966 458108
rect 304998 442856 305054 442912
rect 565818 442856 565874 442912
rect 304262 333784 304318 333840
rect 565726 333784 565782 333840
rect 303434 332424 303490 332480
rect 303618 330540 303674 330576
rect 303618 330520 303620 330540
rect 303620 330520 303672 330540
rect 303672 330520 303674 330540
rect 485594 331744 485650 331800
rect 480534 329024 480590 329080
rect 495438 315968 495494 316024
rect 551374 331744 551430 331800
rect 567750 458632 567806 458688
rect 567658 433336 567714 433392
rect 566554 331336 566610 331392
rect 566462 331200 566518 331256
rect 566370 315832 566426 315888
rect 305182 313928 305238 313984
rect 566462 313928 566518 313984
rect 303526 205536 303582 205592
rect 303802 205808 303858 205864
rect 565726 205808 565782 205864
rect 303710 205672 303766 205728
rect 564438 205536 564494 205592
rect 305182 204992 305238 205048
rect 308494 204176 308550 204232
rect 305182 187584 305238 187640
rect 305734 187620 305736 187640
rect 305736 187620 305788 187640
rect 305788 187620 305790 187640
rect 305734 187584 305790 187620
rect 450174 204312 450230 204368
rect 485594 203496 485650 203552
rect 480534 200640 480590 200696
rect 536194 204040 536250 204096
rect 568670 459584 568726 459640
rect 564346 187584 564402 187640
rect 303618 185816 303674 185872
rect 303526 77832 303582 77888
rect 308494 75792 308550 75848
rect 336738 77832 336794 77888
rect 454038 77832 454094 77888
rect 455326 77832 455382 77888
rect 386418 76608 386474 76664
rect 381358 57296 381414 57352
rect 387798 76472 387854 76528
rect 398838 76744 398894 76800
rect 403070 73752 403126 73808
rect 401598 59880 401654 59936
rect 407118 73888 407174 73944
rect 420182 68856 420238 68912
rect 419998 57160 420054 57216
rect 421838 54576 421894 54632
rect 423678 54440 423734 54496
rect 425518 54440 425574 54496
rect 439502 62736 439558 62792
rect 465722 71712 465778 71768
rect 505834 75112 505890 75168
rect 558182 69672 558238 69728
rect 568026 204312 568082 204368
rect 568854 459584 568910 459640
rect 568762 459448 568818 459504
rect 571338 585792 571394 585848
rect 568854 314608 568910 314664
rect 568854 205536 568910 205592
rect 568578 204040 568634 204096
rect 569958 73888 570014 73944
rect 570326 201320 570382 201376
rect 570234 79328 570290 79384
rect 571430 459584 571486 459640
rect 571430 76064 571486 76120
rect 579618 524476 579674 524512
rect 579618 524456 579620 524476
rect 579620 524456 579672 524476
rect 579672 524456 579674 524476
rect 572994 315968 573050 316024
rect 572994 314744 573050 314800
rect 572902 205808 572958 205864
rect 571338 73752 571394 73808
rect 574098 314744 574154 314800
rect 574190 76472 574246 76528
rect 575570 457408 575626 457464
rect 580906 644000 580962 644056
rect 580354 630808 580410 630864
rect 580262 378392 580318 378448
rect 577686 318008 577742 318064
rect 577594 75792 577650 75848
rect 580906 590960 580962 591016
rect 580538 577632 580594 577688
rect 580446 471416 580502 471472
rect 580354 332424 580410 332480
rect 580906 537784 580962 537840
rect 580630 484628 580686 484664
rect 580630 484608 580632 484628
rect 580632 484608 580684 484628
rect 580684 484608 580686 484628
rect 580906 484608 580962 484664
rect 580906 431568 580962 431624
rect 580906 378392 580962 378448
rect 580630 365064 580686 365120
rect 580446 204176 580502 204232
rect 153106 38664 153162 38720
rect 151726 38120 151782 38176
rect 437386 37576 437442 37632
rect 151634 37168 151690 37224
rect 151174 33088 151230 33144
rect 151082 28464 151138 28520
rect 151082 26424 151138 26480
rect 150438 26188 150440 26208
rect 150440 26188 150492 26208
rect 150492 26188 150494 26208
rect 150438 26152 150494 26188
rect 3422 6432 3478 6488
rect 277306 23432 277362 23488
rect 163686 12960 163742 13016
rect 156602 3304 156658 3360
rect 226890 10240 226946 10296
rect 240138 14456 240194 14512
rect 241978 11600 242034 11656
rect 247682 21392 247738 21448
rect 248418 9016 248474 9072
rect 254950 17176 255006 17232
rect 255318 6296 255374 6352
rect 256790 15816 256846 15872
rect 262034 18536 262090 18592
rect 265070 19896 265126 19952
rect 269210 7656 269266 7712
rect 271970 4936 272026 4992
rect 276202 21256 276258 21312
rect 280066 3440 280122 3496
rect 281262 22072 281318 22128
rect 282918 4800 282974 4856
rect 289358 17312 289414 17368
rect 287150 7520 287206 7576
rect 287058 1944 287114 2000
rect 291474 8880 291530 8936
rect 289818 6160 289874 6216
rect 299478 21392 299534 21448
rect 293958 7656 294014 7712
rect 296074 3440 296130 3496
rect 298742 12960 298798 13016
rect 301502 3440 301558 3496
rect 300490 3304 300546 3360
rect 303158 3440 303214 3496
rect 305642 3304 305698 3360
rect 313830 3304 313886 3360
rect 329102 17312 329158 17368
rect 345294 10240 345350 10296
rect 381726 21256 381782 21312
rect 384302 14456 384358 14512
rect 398930 11600 398986 11656
rect 420182 9016 420238 9072
rect 440238 17176 440294 17232
rect 445022 6296 445078 6352
rect 448610 15816 448666 15872
rect 465170 18536 465226 18592
rect 476118 19896 476174 19952
rect 480258 7520 480314 7576
rect 518898 23432 518954 23488
rect 501786 4936 501842 4992
rect 532698 22072 532754 22128
rect 540794 4800 540850 4856
rect 558550 1944 558606 2000
rect 565634 6160 565690 6216
rect 572718 8880 572774 8936
<< metal3 >>
rect 288934 700300 288940 700364
rect 289004 700362 289010 700364
rect 397453 700362 397519 700365
rect 289004 700360 397519 700362
rect 289004 700304 397458 700360
rect 397514 700304 397519 700360
rect 289004 700302 397519 700304
rect 289004 700300 289010 700302
rect 397453 700299 397519 700302
rect 19241 699820 19307 699821
rect 19190 699818 19196 699820
rect 19150 699758 19196 699818
rect 19260 699816 19307 699820
rect 19302 699760 19307 699816
rect 19190 699756 19196 699758
rect 19260 699756 19307 699760
rect 287646 699756 287652 699820
rect 287716 699818 287722 699820
rect 527265 699818 527331 699821
rect 287716 699816 527331 699818
rect 287716 699760 527270 699816
rect 527326 699760 527331 699816
rect 287716 699758 527331 699760
rect 287716 699756 287722 699758
rect 19241 699755 19307 699756
rect 527265 699755 527331 699758
rect -960 697220 480 697460
rect 303470 697444 303476 697508
rect 303540 697506 303546 697508
rect 527173 697506 527239 697509
rect 303540 697504 527239 697506
rect 303540 697448 527178 697504
rect 527234 697448 527239 697504
rect 303540 697446 527239 697448
rect 303540 697444 303546 697446
rect 527173 697443 527239 697446
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 583520 617388 584960 617628
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 575238 590956 575244 591020
rect 575308 591018 575314 591020
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 575308 591016 584960 591018
rect 575308 590960 580906 591016
rect 580962 590960 584960 591016
rect 575308 590958 584960 590960
rect 575308 590956 575314 590958
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect 23197 585850 23263 585853
rect 63585 585850 63651 585853
rect 23197 585848 63651 585850
rect 23197 585792 23202 585848
rect 23258 585792 63590 585848
rect 63646 585792 63651 585848
rect 23197 585790 63651 585792
rect 23197 585787 23263 585790
rect 63585 585787 63651 585790
rect 149973 585850 150039 585853
rect 292614 585850 292620 585852
rect 149973 585848 292620 585850
rect 149973 585792 149978 585848
rect 150034 585792 292620 585848
rect 149973 585790 292620 585792
rect 149973 585787 150039 585790
rect 292614 585788 292620 585790
rect 292684 585788 292690 585852
rect 297950 585788 297956 585852
rect 298020 585850 298026 585852
rect 485589 585850 485655 585853
rect 298020 585848 485655 585850
rect 298020 585792 485594 585848
rect 485650 585792 485655 585848
rect 298020 585790 485655 585792
rect 298020 585788 298026 585790
rect 485589 585787 485655 585790
rect 556429 585850 556495 585853
rect 571333 585850 571399 585853
rect 556429 585848 571399 585850
rect 556429 585792 556434 585848
rect 556490 585792 571338 585848
rect 571394 585792 571399 585848
rect 556429 585790 571399 585792
rect 556429 585787 556495 585790
rect 571333 585787 571399 585790
rect 23238 585652 23244 585716
rect 23308 585714 23314 585716
rect 83825 585714 83891 585717
rect 23308 585712 83891 585714
rect 23308 585656 83830 585712
rect 83886 585656 83891 585712
rect 23308 585654 83891 585656
rect 23308 585652 23314 585654
rect 83825 585651 83891 585654
rect 226149 585714 226215 585717
rect 287513 585714 287579 585717
rect 226149 585712 287579 585714
rect 226149 585656 226154 585712
rect 226210 585656 287518 585712
rect 287574 585656 287579 585712
rect 226149 585654 287579 585656
rect 226149 585651 226215 585654
rect 287513 585651 287579 585654
rect 292430 585652 292436 585716
rect 292500 585714 292506 585716
rect 480529 585714 480595 585717
rect 292500 585712 480595 585714
rect 292500 585656 480534 585712
rect 480590 585656 480595 585712
rect 292500 585654 480595 585656
rect 292500 585652 292506 585654
rect 480529 585651 480595 585654
rect 551369 585714 551435 585717
rect 571374 585714 571380 585716
rect 551369 585712 571380 585714
rect 551369 585656 551374 585712
rect 551430 585656 571380 585712
rect 551369 585654 571380 585656
rect 551369 585651 551435 585654
rect 571374 585652 571380 585654
rect 571444 585652 571450 585716
rect 286174 585108 286180 585172
rect 286244 585170 286250 585172
rect 286409 585170 286475 585173
rect 286244 585168 286475 585170
rect 286244 585112 286414 585168
rect 286470 585112 286475 585168
rect 286244 585110 286475 585112
rect 286244 585108 286250 585110
rect 286409 585107 286475 585110
rect 566549 585170 566615 585173
rect 566958 585170 566964 585172
rect 566549 585168 566964 585170
rect 566549 585112 566554 585168
rect 566610 585112 566964 585168
rect 566549 585110 566964 585112
rect 566549 585107 566615 585110
rect 566958 585108 566964 585110
rect 567028 585108 567034 585172
rect 505829 583130 505895 583133
rect 565854 583130 565860 583132
rect 505829 583128 565860 583130
rect 505829 583072 505834 583128
rect 505890 583072 565860 583128
rect 505829 583070 565860 583072
rect 505829 583067 505895 583070
rect 565854 583068 565860 583070
rect 565924 583068 565930 583132
rect 17718 582932 17724 582996
rect 17788 582994 17794 582996
rect 134425 582994 134491 582997
rect 17788 582992 134491 582994
rect 17788 582936 134430 582992
rect 134486 582936 134491 582992
rect 17788 582934 134491 582936
rect 17788 582932 17794 582934
rect 134425 582931 134491 582934
rect 210969 582994 211035 582997
rect 285622 582994 285628 582996
rect 210969 582992 285628 582994
rect 210969 582936 210974 582992
rect 211030 582936 285628 582992
rect 210969 582934 285628 582936
rect 210969 582931 211035 582934
rect 285622 582932 285628 582934
rect 285692 582932 285698 582996
rect 298001 582994 298067 582997
rect 369209 582994 369275 582997
rect 298001 582992 369275 582994
rect 298001 582936 298006 582992
rect 298062 582936 369214 582992
rect 369270 582936 369275 582992
rect 298001 582934 369275 582936
rect 298001 582931 298067 582934
rect 369209 582931 369275 582934
rect 490649 582994 490715 582997
rect 566038 582994 566044 582996
rect 490649 582992 566044 582994
rect 490649 582936 490654 582992
rect 490710 582936 566044 582992
rect 490649 582934 566044 582936
rect 490649 582931 490715 582934
rect 566038 582932 566044 582934
rect 566108 582932 566114 582996
rect 450169 580410 450235 580413
rect 567326 580410 567332 580412
rect 450169 580408 567332 580410
rect 450169 580352 450174 580408
rect 450230 580352 567332 580408
rect 450169 580350 567332 580352
rect 450169 580347 450235 580350
rect 567326 580348 567332 580350
rect 567396 580348 567402 580412
rect 175181 580274 175247 580277
rect 290038 580274 290044 580276
rect 175181 580272 290044 580274
rect 175181 580216 175186 580272
rect 175242 580216 290044 580272
rect 175181 580214 290044 580216
rect 175181 580211 175247 580214
rect 290038 580212 290044 580214
rect 290108 580212 290114 580276
rect 301630 580212 301636 580276
rect 301700 580274 301706 580276
rect 389449 580274 389515 580277
rect 301700 580272 389515 580274
rect 301700 580216 389454 580272
rect 389510 580216 389515 580272
rect 301700 580214 389515 580216
rect 301700 580212 301706 580214
rect 389449 580211 389515 580214
rect 440049 580274 440115 580277
rect 570086 580274 570092 580276
rect 440049 580272 570092 580274
rect 440049 580216 440054 580272
rect 440110 580216 570092 580272
rect 440049 580214 570092 580216
rect 440049 580211 440115 580214
rect 570086 580212 570092 580214
rect 570156 580212 570162 580276
rect -960 579852 480 580092
rect 580533 577690 580599 577693
rect 583520 577690 584960 577780
rect 580533 577688 584960 577690
rect 580533 577632 580538 577688
rect 580594 577632 584960 577688
rect 580533 577630 584960 577632
rect 580533 577627 580599 577630
rect 583520 577540 584960 577630
rect 276013 572114 276079 572117
rect 295926 572114 295932 572116
rect 276013 572112 295932 572114
rect 276013 572056 276018 572112
rect 276074 572056 295932 572112
rect 276013 572054 295932 572056
rect 276013 572051 276079 572054
rect 295926 572052 295932 572054
rect 295996 572052 296002 572116
rect 20345 571978 20411 571981
rect 109033 571978 109099 571981
rect 20345 571976 109099 571978
rect 20345 571920 20350 571976
rect 20406 571920 109038 571976
rect 109094 571920 109099 571976
rect 20345 571918 109099 571920
rect 20345 571915 20411 571918
rect 109033 571915 109099 571918
rect 204253 571978 204319 571981
rect 292798 571978 292804 571980
rect 204253 571976 292804 571978
rect 204253 571920 204258 571976
rect 204314 571920 292804 571976
rect 204253 571918 292804 571920
rect 204253 571915 204319 571918
rect 292798 571916 292804 571918
rect 292868 571916 292874 571980
rect 302182 571916 302188 571980
rect 302252 571978 302258 571980
rect 404353 571978 404419 571981
rect 302252 571976 404419 571978
rect 302252 571920 404358 571976
rect 404414 571920 404419 571976
rect 302252 571918 404419 571920
rect 302252 571916 302258 571918
rect 404353 571915 404419 571918
rect 434713 571978 434779 571981
rect 568614 571978 568620 571980
rect 434713 571976 568620 571978
rect 434713 571920 434718 571976
rect 434774 571920 568620 571976
rect 434713 571918 568620 571920
rect 434713 571915 434779 571918
rect 568614 571916 568620 571918
rect 568684 571916 568690 571980
rect 21950 570556 21956 570620
rect 22020 570618 22026 570620
rect 39297 570618 39363 570621
rect 22020 570616 39363 570618
rect 22020 570560 39302 570616
rect 39358 570560 39363 570616
rect 22020 570558 39363 570560
rect 22020 570556 22026 570558
rect 39297 570555 39363 570558
rect 288198 570556 288204 570620
rect 288268 570618 288274 570620
rect 424317 570618 424383 570621
rect 288268 570616 424383 570618
rect 288268 570560 424322 570616
rect 424378 570560 424383 570616
rect 288268 570558 424383 570560
rect 288268 570556 288274 570558
rect 424317 570555 424383 570558
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 579613 524514 579679 524517
rect 583520 524514 584960 524604
rect 579613 524512 584960 524514
rect 579613 524456 579618 524512
rect 579674 524456 584960 524512
rect 579613 524454 584960 524456
rect 579613 524451 579679 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2865 514858 2931 514861
rect -960 514856 2931 514858
rect -960 514800 2870 514856
rect 2926 514800 2931 514856
rect -960 514798 2931 514800
rect -960 514708 480 514798
rect 2865 514795 2931 514798
rect 583520 511172 584960 511412
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580625 484666 580691 484669
rect 580901 484666 580967 484669
rect 583520 484666 584960 484756
rect 580625 484664 584960 484666
rect 580625 484608 580630 484664
rect 580686 484608 580906 484664
rect 580962 484608 584960 484664
rect 580625 484606 584960 484608
rect 580625 484603 580691 484606
rect 580901 484603 580967 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 580441 471474 580507 471477
rect 583520 471474 584960 471564
rect 580441 471472 584960 471474
rect 580441 471416 580446 471472
rect 580502 471416 584960 471472
rect 580441 471414 584960 471416
rect 580441 471411 580507 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 286225 461956 286291 461957
rect 303521 461956 303587 461957
rect 286174 461954 286180 461956
rect 286134 461894 286180 461954
rect 286244 461952 286291 461956
rect 286286 461896 286291 461952
rect 286174 461892 286180 461894
rect 286244 461892 286291 461896
rect 303470 461892 303476 461956
rect 303540 461954 303587 461956
rect 303540 461952 303632 461954
rect 303582 461896 303632 461952
rect 303540 461894 303632 461896
rect 303540 461892 303587 461894
rect 286225 461891 286291 461892
rect 303521 461891 303587 461892
rect 301998 461756 302004 461820
rect 302068 461818 302074 461820
rect 305085 461818 305151 461821
rect 302068 461816 305151 461818
rect 302068 461760 305090 461816
rect 305146 461760 305151 461816
rect 302068 461758 305151 461760
rect 302068 461756 302074 461758
rect 305085 461755 305151 461758
rect 565721 461002 565787 461005
rect 568614 461002 568620 461004
rect 565721 461000 568620 461002
rect 565721 460944 565726 461000
rect 565782 460944 568620 461000
rect 565721 460942 568620 460944
rect 565721 460939 565787 460942
rect 568614 460940 568620 460942
rect 568684 460940 568690 461004
rect 160001 460866 160067 460869
rect 160001 460864 277410 460866
rect 160001 460808 160006 460864
rect 160062 460808 277410 460864
rect 160001 460806 277410 460808
rect 160001 460803 160067 460806
rect 21950 460260 21956 460324
rect 22020 460322 22026 460324
rect 24853 460322 24919 460325
rect 124305 460322 124371 460325
rect 22020 460320 124371 460322
rect 22020 460264 24858 460320
rect 24914 460264 124310 460320
rect 124366 460264 124371 460320
rect 22020 460262 124371 460264
rect 277350 460322 277410 460806
rect 286174 460668 286180 460732
rect 286244 460730 286250 460732
rect 286317 460730 286383 460733
rect 286244 460728 286383 460730
rect 286244 460672 286322 460728
rect 286378 460672 286383 460728
rect 286244 460670 286383 460672
rect 286244 460668 286250 460670
rect 286317 460667 286383 460670
rect 288709 460322 288775 460325
rect 277350 460320 288775 460322
rect 277350 460264 288714 460320
rect 288770 460264 288775 460320
rect 277350 460262 288775 460264
rect 22020 460260 22026 460262
rect 24853 460259 24919 460262
rect 124305 460259 124371 460262
rect 288709 460259 288775 460262
rect 564893 460322 564959 460325
rect 570086 460322 570092 460324
rect 564893 460320 570092 460322
rect 564893 460264 564898 460320
rect 564954 460264 570092 460320
rect 564893 460262 570092 460264
rect 564893 460259 564959 460262
rect 570086 460260 570092 460262
rect 570156 460260 570162 460324
rect 16389 460186 16455 460189
rect 17718 460186 17724 460188
rect 16389 460184 17724 460186
rect 16389 460128 16394 460184
rect 16450 460128 17724 460184
rect 16389 460126 17724 460128
rect 16389 460123 16455 460126
rect 17718 460124 17724 460126
rect 17788 460186 17794 460188
rect 134425 460186 134491 460189
rect 17788 460184 134491 460186
rect 17788 460128 134430 460184
rect 134486 460128 134491 460184
rect 17788 460126 134491 460128
rect 17788 460124 17794 460126
rect 134425 460123 134491 460126
rect 175181 460186 175247 460189
rect 285305 460186 285371 460189
rect 290038 460186 290044 460188
rect 175181 460184 290044 460186
rect 175181 460128 175186 460184
rect 175242 460128 285310 460184
rect 285366 460128 290044 460184
rect 175181 460126 290044 460128
rect 175181 460123 175247 460126
rect 285305 460123 285371 460126
rect 290038 460124 290044 460126
rect 290108 460124 290114 460188
rect 455229 460186 455295 460189
rect 570086 460186 570092 460188
rect 455229 460184 570092 460186
rect 455229 460128 455234 460184
rect 455290 460128 570092 460184
rect 455229 460126 570092 460128
rect 455229 460123 455295 460126
rect 570086 460124 570092 460126
rect 570156 460124 570162 460188
rect 288709 459778 288775 459781
rect 291377 459778 291443 459781
rect 288709 459776 291443 459778
rect 288709 459720 288714 459776
rect 288770 459720 291382 459776
rect 291438 459720 291443 459776
rect 288709 459718 291443 459720
rect 288709 459715 288775 459718
rect 291377 459715 291443 459718
rect 287605 459642 287671 459645
rect 289854 459642 289860 459644
rect 287605 459640 289860 459642
rect 287605 459584 287610 459640
rect 287666 459584 289860 459640
rect 287605 459582 289860 459584
rect 287605 459579 287671 459582
rect 289854 459580 289860 459582
rect 289924 459580 289930 459644
rect 556153 459642 556219 459645
rect 568665 459642 568731 459645
rect 568849 459642 568915 459645
rect 556153 459640 568915 459642
rect 556153 459584 556158 459640
rect 556214 459584 568670 459640
rect 568726 459584 568854 459640
rect 568910 459584 568915 459640
rect 556153 459582 568915 459584
rect 556153 459579 556219 459582
rect 568665 459579 568731 459582
rect 568849 459579 568915 459582
rect 570086 459580 570092 459644
rect 570156 459642 570162 459644
rect 571425 459642 571491 459645
rect 570156 459640 571491 459642
rect 570156 459584 571430 459640
rect 571486 459584 571491 459640
rect 570156 459582 571491 459584
rect 570156 459580 570162 459582
rect 571425 459579 571491 459582
rect 281441 459506 281507 459509
rect 287697 459506 287763 459509
rect 281441 459504 287763 459506
rect 281441 459448 281446 459504
rect 281502 459448 287702 459504
rect 287758 459448 287763 459504
rect 281441 459446 287763 459448
rect 281441 459443 281507 459446
rect 287697 459443 287763 459446
rect 301630 459444 301636 459508
rect 301700 459506 301706 459508
rect 301865 459506 301931 459509
rect 301700 459504 301931 459506
rect 301700 459448 301870 459504
rect 301926 459448 301931 459504
rect 301700 459446 301931 459448
rect 301700 459444 301706 459446
rect 301865 459443 301931 459446
rect 561489 459506 561555 459509
rect 568757 459506 568823 459509
rect 561489 459504 568823 459506
rect 561489 459448 561494 459504
rect 561550 459448 568762 459504
rect 568818 459448 568823 459504
rect 561489 459446 568823 459448
rect 561489 459443 561555 459446
rect 568757 459443 568823 459446
rect 276749 459098 276815 459101
rect 302734 459098 302740 459100
rect 276749 459096 302740 459098
rect 276749 459040 276754 459096
rect 276810 459040 302740 459096
rect 276749 459038 302740 459040
rect 276749 459035 276815 459038
rect 302734 459036 302740 459038
rect 302804 459036 302810 459100
rect 303153 459098 303219 459101
rect 313273 459098 313339 459101
rect 303153 459096 313339 459098
rect 303153 459040 303158 459096
rect 303214 459040 313278 459096
rect 313334 459040 313339 459096
rect 303153 459038 313339 459040
rect 303153 459035 303219 459038
rect 313273 459035 313339 459038
rect 564433 459098 564499 459101
rect 565670 459098 565676 459100
rect 564433 459096 565676 459098
rect 564433 459040 564438 459096
rect 564494 459040 565676 459096
rect 564433 459038 565676 459040
rect 564433 459035 564499 459038
rect 565670 459036 565676 459038
rect 565740 459098 565746 459100
rect 567326 459098 567332 459100
rect 565740 459038 567332 459098
rect 565740 459036 565746 459038
rect 567326 459036 567332 459038
rect 567396 459036 567402 459100
rect 22921 458962 22987 458965
rect 34513 458962 34579 458965
rect 22921 458960 34579 458962
rect 22921 458904 22926 458960
rect 22982 458904 34518 458960
rect 34574 458904 34579 458960
rect 22921 458902 34579 458904
rect 22921 458899 22987 458902
rect 34513 458899 34579 458902
rect 286869 458962 286935 458965
rect 299974 458962 299980 458964
rect 286869 458960 299980 458962
rect 286869 458904 286874 458960
rect 286930 458904 299980 458960
rect 286869 458902 299980 458904
rect 286869 458899 286935 458902
rect 299974 458900 299980 458902
rect 300044 458900 300050 458964
rect 301446 458900 301452 458964
rect 301516 458962 301522 458964
rect 485589 458962 485655 458965
rect 301516 458960 485655 458962
rect 301516 458904 485594 458960
rect 485650 458904 485655 458960
rect 301516 458902 485655 458904
rect 301516 458900 301522 458902
rect 485589 458899 485655 458902
rect 18781 458826 18847 458829
rect 93945 458826 94011 458829
rect 18781 458824 94011 458826
rect 18781 458768 18786 458824
rect 18842 458768 93950 458824
rect 94006 458768 94011 458824
rect 18781 458766 94011 458768
rect 18781 458763 18847 458766
rect 93945 458763 94011 458766
rect 295006 458764 295012 458828
rect 295076 458826 295082 458828
rect 480529 458826 480595 458829
rect 295076 458824 480595 458826
rect 295076 458768 480534 458824
rect 480590 458768 480595 458824
rect 295076 458766 480595 458768
rect 295076 458764 295082 458766
rect 480529 458763 480595 458766
rect 551369 458826 551435 458829
rect 567326 458826 567332 458828
rect 551369 458824 567332 458826
rect 551369 458768 551374 458824
rect 551430 458768 567332 458824
rect 551369 458766 567332 458768
rect 551369 458763 551435 458766
rect 567326 458764 567332 458766
rect 567396 458764 567402 458828
rect 567745 458690 567811 458693
rect 568614 458690 568620 458692
rect 567745 458688 568620 458690
rect 567745 458632 567750 458688
rect 567806 458632 568620 458688
rect 567745 458630 568620 458632
rect 567745 458627 567811 458630
rect 568614 458628 568620 458630
rect 568684 458628 568690 458692
rect 285397 458284 285463 458285
rect 285397 458280 285444 458284
rect 285508 458282 285514 458284
rect 300485 458282 300551 458285
rect 301630 458282 301636 458284
rect 285397 458224 285402 458280
rect 285397 458220 285444 458224
rect 285508 458222 285554 458282
rect 300485 458280 301636 458282
rect 300485 458224 300490 458280
rect 300546 458224 301636 458280
rect 300485 458222 301636 458224
rect 285508 458220 285514 458222
rect 285397 458219 285463 458220
rect 300485 458219 300551 458222
rect 301630 458220 301636 458222
rect 301700 458220 301706 458284
rect 23238 458084 23244 458148
rect 23308 458146 23314 458148
rect 83825 458146 83891 458149
rect 23308 458144 83891 458146
rect 23308 458088 83830 458144
rect 83886 458088 83891 458144
rect 23308 458086 83891 458088
rect 23308 458084 23314 458086
rect 83825 458083 83891 458086
rect 211153 458146 211219 458149
rect 285622 458146 285628 458148
rect 211153 458144 285628 458146
rect 211153 458088 211158 458144
rect 211214 458088 285628 458144
rect 211153 458086 285628 458088
rect 211153 458083 211219 458086
rect 285622 458084 285628 458086
rect 285692 458146 285698 458148
rect 490649 458146 490715 458149
rect 565905 458148 565971 458149
rect 285692 458086 287070 458146
rect 285692 458084 285698 458086
rect 287010 458010 287070 458086
rect 490649 458144 547890 458146
rect 490649 458088 490654 458144
rect 490710 458088 547890 458144
rect 490649 458086 547890 458088
rect 490649 458083 490715 458086
rect 287605 458010 287671 458013
rect 287010 458008 287671 458010
rect 287010 457952 287610 458008
rect 287666 457952 287671 458008
rect 287010 457950 287671 457952
rect 287605 457947 287671 457950
rect 547830 457466 547890 458086
rect 565854 458084 565860 458148
rect 565924 458146 565971 458148
rect 565924 458144 566016 458146
rect 565966 458088 566016 458144
rect 565924 458086 566016 458088
rect 565924 458084 565971 458086
rect 565905 458083 565971 458084
rect 583520 457996 584960 458236
rect 566038 457466 566044 457468
rect 547830 457406 566044 457466
rect 566038 457404 566044 457406
rect 566108 457466 566114 457468
rect 575565 457466 575631 457469
rect 566108 457464 575631 457466
rect 566108 457408 575570 457464
rect 575626 457408 575631 457464
rect 566108 457406 575631 457408
rect 566108 457404 566114 457406
rect 575565 457403 575631 457406
rect 21950 456860 21956 456924
rect 22020 456922 22026 456924
rect 23238 456922 23244 456924
rect 22020 456862 23244 456922
rect 22020 456860 22026 456862
rect 23238 456860 23244 456862
rect 23308 456860 23314 456924
rect 286225 456922 286291 456925
rect 286358 456922 286364 456924
rect 286225 456920 286364 456922
rect 286225 456864 286230 456920
rect 286286 456864 286364 456920
rect 286225 456862 286364 456864
rect 286225 456859 286291 456862
rect 286358 456860 286364 456862
rect 286428 456860 286434 456924
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 583520 444668 584960 444908
rect 23238 444212 23244 444276
rect 23308 444274 23314 444276
rect 24945 444274 25011 444277
rect 23308 444272 25011 444274
rect 23308 444216 24950 444272
rect 25006 444216 25011 444272
rect 23308 444214 25011 444216
rect 23308 444212 23314 444214
rect 24945 444211 25011 444214
rect 297173 444002 297239 444005
rect 297766 444002 297772 444004
rect 297173 444000 297772 444002
rect 297173 443944 297178 444000
rect 297234 443944 297772 444000
rect 297173 443942 297772 443944
rect 297173 443939 297239 443942
rect 297766 443940 297772 443942
rect 297836 443940 297842 444004
rect 285397 443866 285463 443869
rect 290038 443866 290044 443868
rect 285397 443864 290044 443866
rect 285397 443808 285402 443864
rect 285458 443808 290044 443864
rect 285397 443806 290044 443808
rect 285397 443803 285463 443806
rect 290038 443804 290044 443806
rect 290108 443804 290114 443868
rect 204253 443730 204319 443733
rect 291142 443730 291148 443732
rect 204253 443728 291148 443730
rect 204253 443672 204258 443728
rect 204314 443672 291148 443728
rect 204253 443670 291148 443672
rect 204253 443667 204319 443670
rect 291142 443668 291148 443670
rect 291212 443668 291218 443732
rect 298686 443668 298692 443732
rect 298756 443730 298762 443732
rect 414013 443730 414079 443733
rect 298756 443728 414079 443730
rect 298756 443672 414018 443728
rect 414074 443672 414079 443728
rect 298756 443670 414079 443672
rect 298756 443668 298762 443670
rect 414013 443667 414079 443670
rect 289118 443532 289124 443596
rect 289188 443594 289194 443596
rect 424317 443594 424383 443597
rect 289188 443592 424383 443594
rect 289188 443536 424322 443592
rect 424378 443536 424383 443592
rect 289188 443534 424383 443536
rect 289188 443532 289194 443534
rect 424317 443531 424383 443534
rect 297909 442914 297975 442917
rect 298686 442914 298692 442916
rect 297909 442912 298692 442914
rect 297909 442856 297914 442912
rect 297970 442856 298692 442912
rect 297909 442854 298692 442856
rect 297909 442851 297975 442854
rect 298686 442852 298692 442854
rect 298756 442852 298762 442916
rect 301998 442852 302004 442916
rect 302068 442914 302074 442916
rect 304993 442914 305059 442917
rect 302068 442912 305059 442914
rect 302068 442856 304998 442912
rect 305054 442856 305059 442912
rect 302068 442854 305059 442856
rect 302068 442852 302074 442854
rect 304993 442851 305059 442854
rect 565813 442914 565879 442917
rect 566590 442914 566596 442916
rect 565813 442912 566596 442914
rect 565813 442856 565818 442912
rect 565874 442856 566596 442912
rect 565813 442854 566596 442856
rect 565813 442851 565879 442854
rect 566590 442852 566596 442854
rect 566660 442852 566666 442916
rect -960 436508 480 436748
rect 285438 433876 285444 433940
rect 285508 433938 285514 433940
rect 290089 433938 290155 433941
rect 285508 433936 290155 433938
rect 285508 433880 290094 433936
rect 290150 433880 290155 433936
rect 285508 433878 290155 433880
rect 285508 433876 285514 433878
rect 290089 433875 290155 433878
rect 565670 433332 565676 433396
rect 565740 433394 565746 433396
rect 567653 433394 567719 433397
rect 565740 433392 567719 433394
rect 565740 433336 567658 433392
rect 567714 433336 567719 433392
rect 565740 433334 567719 433336
rect 565740 433332 565746 433334
rect 567653 433331 567719 433334
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 569166 418236 569172 418300
rect 569236 418298 569242 418300
rect 583520 418298 584960 418388
rect 569236 418238 584960 418298
rect 569236 418236 569242 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580257 378450 580323 378453
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 580906 378448
rect 580962 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 580625 365122 580691 365125
rect 583520 365122 584960 365212
rect 580625 365120 584960 365122
rect 580625 365064 580630 365120
rect 580686 365064 584960 365120
rect 580625 365062 584960 365064
rect 580625 365059 580691 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2957 358458 3023 358461
rect -960 358456 3023 358458
rect -960 358400 2962 358456
rect 3018 358400 3023 358456
rect -960 358398 3023 358400
rect -960 358308 480 358398
rect 2957 358395 3023 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect 570086 334658 570092 334660
rect 565678 334598 570092 334658
rect 288617 334250 288683 334253
rect 285814 334248 288683 334250
rect 285814 334192 288622 334248
rect 288678 334192 288683 334248
rect 285814 334190 288683 334192
rect 285814 333845 285874 334190
rect 288617 334187 288683 334190
rect 286358 334052 286364 334116
rect 286428 334114 286434 334116
rect 290089 334114 290155 334117
rect 286428 334054 286978 334114
rect 286428 334052 286434 334054
rect 285765 333840 285874 333845
rect 285765 333784 285770 333840
rect 285826 333784 285874 333840
rect 285765 333782 285874 333784
rect 286918 333845 286978 334054
rect 287102 334112 290155 334114
rect 287102 334056 290094 334112
rect 290150 334056 290155 334112
rect 287102 334054 290155 334056
rect 286918 333840 287027 333845
rect 286918 333784 286966 333840
rect 287022 333784 287027 333840
rect 286918 333782 287027 333784
rect 285765 333779 285831 333782
rect 286961 333779 287027 333782
rect 286869 333706 286935 333709
rect 287102 333706 287162 334054
rect 290089 334051 290155 334054
rect 301998 334052 302004 334116
rect 302068 334114 302074 334116
rect 302068 334054 303722 334114
rect 302068 334052 302074 334054
rect 303662 333842 303722 334054
rect 565678 333845 565738 334598
rect 570086 334596 570092 334598
rect 570156 334596 570162 334660
rect 304257 333842 304323 333845
rect 303662 333840 304323 333842
rect 303662 333784 304262 333840
rect 304318 333784 304323 333840
rect 303662 333782 304323 333784
rect 565678 333840 565787 333845
rect 565678 333784 565726 333840
rect 565782 333784 565787 333840
rect 565678 333782 565787 333784
rect 304257 333779 304323 333782
rect 565721 333779 565787 333782
rect 286869 333704 287162 333706
rect 286869 333648 286874 333704
rect 286930 333648 287162 333704
rect 286869 333646 287162 333648
rect 286869 333643 286935 333646
rect 3509 332482 3575 332485
rect 28165 332482 28231 332485
rect 3509 332480 28231 332482
rect -960 332196 480 332436
rect 3509 332424 3514 332480
rect 3570 332424 28170 332480
rect 28226 332424 28231 332480
rect 3509 332422 28231 332424
rect 3509 332419 3575 332422
rect 28165 332419 28231 332422
rect 241329 332482 241395 332485
rect 289905 332484 289971 332485
rect 289854 332482 289860 332484
rect 241329 332480 289860 332482
rect 289924 332480 289971 332484
rect 241329 332424 241334 332480
rect 241390 332424 289860 332480
rect 289966 332424 289971 332480
rect 241329 332422 289860 332424
rect 241329 332419 241395 332422
rect 289854 332420 289860 332422
rect 289924 332420 289971 332424
rect 289905 332419 289971 332420
rect 303429 332482 303495 332485
rect 580349 332482 580415 332485
rect 303429 332480 580415 332482
rect 303429 332424 303434 332480
rect 303490 332424 580354 332480
rect 580410 332424 580415 332480
rect 303429 332422 580415 332424
rect 303429 332419 303495 332422
rect 580349 332419 580415 332422
rect 285673 332210 285739 332213
rect 286174 332210 286180 332212
rect 285673 332208 286180 332210
rect 285673 332152 285678 332208
rect 285734 332152 286180 332208
rect 285673 332150 286180 332152
rect 285673 332147 285739 332150
rect 286174 332148 286180 332150
rect 286244 332148 286250 332212
rect 293217 331938 293283 331941
rect 301630 331938 301636 331940
rect 293217 331936 301636 331938
rect 293217 331880 293222 331936
rect 293278 331880 301636 331936
rect 293217 331878 301636 331880
rect 293217 331875 293283 331878
rect 301630 331876 301636 331878
rect 301700 331876 301706 331940
rect 21633 331802 21699 331805
rect 22645 331802 22711 331805
rect 68645 331802 68711 331805
rect 21633 331800 68711 331802
rect 21633 331744 21638 331800
rect 21694 331744 22650 331800
rect 22706 331744 68650 331800
rect 68706 331744 68711 331800
rect 21633 331742 68711 331744
rect 21633 331739 21699 331742
rect 22645 331739 22711 331742
rect 68645 331739 68711 331742
rect 149605 331802 149671 331805
rect 289854 331802 289860 331804
rect 149605 331800 289860 331802
rect 149605 331744 149610 331800
rect 149666 331744 289860 331800
rect 149605 331742 289860 331744
rect 149605 331739 149671 331742
rect 289854 331740 289860 331742
rect 289924 331740 289930 331804
rect 300117 331802 300183 331805
rect 485589 331802 485655 331805
rect 300117 331800 485655 331802
rect 300117 331744 300122 331800
rect 300178 331744 485594 331800
rect 485650 331744 485655 331800
rect 300117 331742 485655 331744
rect 300117 331739 300183 331742
rect 485589 331739 485655 331742
rect 551369 331802 551435 331805
rect 570086 331802 570092 331804
rect 551369 331800 570092 331802
rect 551369 331744 551374 331800
rect 551430 331744 570092 331800
rect 551369 331742 570092 331744
rect 551369 331739 551435 331742
rect 570086 331740 570092 331742
rect 570156 331740 570162 331804
rect 565854 331332 565860 331396
rect 565924 331394 565930 331396
rect 566549 331394 566615 331397
rect 565924 331392 566615 331394
rect 565924 331336 566554 331392
rect 566610 331336 566615 331392
rect 565924 331334 566615 331336
rect 565924 331332 565930 331334
rect 566549 331331 566615 331334
rect 286685 331258 286751 331261
rect 286910 331258 286916 331260
rect 286685 331256 286916 331258
rect 286685 331200 286690 331256
rect 286746 331200 286916 331256
rect 286685 331198 286916 331200
rect 286685 331195 286751 331198
rect 286910 331196 286916 331198
rect 286980 331196 286986 331260
rect 566457 331258 566523 331261
rect 566590 331258 566596 331260
rect 566457 331256 566596 331258
rect 566457 331200 566462 331256
rect 566518 331200 566596 331256
rect 566457 331198 566596 331200
rect 566457 331195 566523 331198
rect 566590 331196 566596 331198
rect 566660 331196 566666 331260
rect 23238 330924 23244 330988
rect 23308 330986 23314 330988
rect 23381 330986 23447 330989
rect 23308 330984 23447 330986
rect 23308 330928 23386 330984
rect 23442 330928 23447 330984
rect 23308 330926 23447 330928
rect 23308 330924 23314 330926
rect 23381 330923 23447 330926
rect 298686 330516 298692 330580
rect 298756 330578 298762 330580
rect 303613 330578 303679 330581
rect 298756 330576 303679 330578
rect 298756 330520 303618 330576
rect 303674 330520 303679 330576
rect 298756 330518 303679 330520
rect 298756 330516 298762 330518
rect 303613 330515 303679 330518
rect 21766 330380 21772 330444
rect 21836 330442 21842 330444
rect 160093 330442 160159 330445
rect 21836 330440 160159 330442
rect 21836 330384 160098 330440
rect 160154 330384 160159 330440
rect 21836 330382 160159 330384
rect 21836 330380 21842 330382
rect 160093 330379 160159 330382
rect 298686 329700 298692 329764
rect 298756 329762 298762 329764
rect 299105 329762 299171 329765
rect 298756 329760 299171 329762
rect 298756 329704 299110 329760
rect 299166 329704 299171 329760
rect 298756 329702 299171 329704
rect 298756 329700 298762 329702
rect 299105 329699 299171 329702
rect 296110 329020 296116 329084
rect 296180 329082 296186 329084
rect 480529 329082 480595 329085
rect 296180 329080 480595 329082
rect 296180 329024 480534 329080
rect 480590 329024 480595 329080
rect 296180 329022 480595 329024
rect 296180 329020 296186 329022
rect 480529 329019 480595 329022
rect 583520 325124 584960 325364
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 303470 318004 303476 318068
rect 303540 318066 303546 318068
rect 577681 318066 577747 318069
rect 303540 318064 577747 318066
rect 303540 318008 577686 318064
rect 577742 318008 577747 318064
rect 303540 318006 577747 318008
rect 303540 318004 303546 318006
rect 577681 318003 577747 318006
rect 285397 316708 285463 316709
rect 285397 316704 285444 316708
rect 285508 316706 285514 316708
rect 290038 316706 290044 316708
rect 285397 316648 285402 316704
rect 285397 316644 285444 316648
rect 285508 316646 290044 316706
rect 285508 316644 285514 316646
rect 290038 316644 290044 316646
rect 290108 316644 290114 316708
rect 285397 316643 285463 316644
rect 495433 316026 495499 316029
rect 572989 316026 573055 316029
rect 495433 316024 573055 316026
rect 495433 315968 495438 316024
rect 495494 315968 572994 316024
rect 573050 315968 573055 316024
rect 495433 315966 573055 315968
rect 495433 315963 495499 315966
rect 572989 315963 573055 315966
rect 22001 315892 22067 315893
rect 21950 315828 21956 315892
rect 22020 315890 22067 315892
rect 566365 315892 566431 315893
rect 22020 315888 22112 315890
rect 22062 315832 22112 315888
rect 22020 315830 22112 315832
rect 566365 315888 566412 315892
rect 566476 315890 566482 315892
rect 566365 315832 566370 315888
rect 22020 315828 22067 315830
rect 22001 315827 22067 315828
rect 566365 315828 566412 315832
rect 566476 315830 566522 315890
rect 566476 315828 566482 315830
rect 566365 315827 566431 315828
rect 286961 315482 287027 315485
rect 300158 315482 300164 315484
rect 286961 315480 300164 315482
rect 286961 315424 286966 315480
rect 287022 315424 300164 315480
rect 286961 315422 300164 315424
rect 286961 315419 287027 315422
rect 300158 315420 300164 315422
rect 300228 315420 300234 315484
rect 20478 315284 20484 315348
rect 20548 315346 20554 315348
rect 171777 315346 171843 315349
rect 20548 315344 171843 315346
rect 20548 315288 171782 315344
rect 171838 315288 171843 315344
rect 20548 315286 171843 315288
rect 20548 315284 20554 315286
rect 171777 315283 171843 315286
rect 204253 315346 204319 315349
rect 290038 315346 290044 315348
rect 204253 315344 290044 315346
rect 204253 315288 204258 315344
rect 204314 315288 290044 315344
rect 204253 315286 290044 315288
rect 204253 315283 204319 315286
rect 290038 315284 290044 315286
rect 290108 315284 290114 315348
rect 21214 314740 21220 314804
rect 21284 314802 21290 314804
rect 21950 314802 21956 314804
rect 21284 314742 21956 314802
rect 21284 314740 21290 314742
rect 21950 314740 21956 314742
rect 22020 314740 22026 314804
rect 572989 314802 573055 314805
rect 574093 314802 574159 314805
rect 572989 314800 574159 314802
rect 572989 314744 572994 314800
rect 573050 314744 574098 314800
rect 574154 314744 574159 314800
rect 572989 314742 574159 314744
rect 572989 314739 573055 314742
rect 574093 314739 574159 314742
rect 568614 314604 568620 314668
rect 568684 314666 568690 314668
rect 568849 314666 568915 314669
rect 568684 314664 568915 314666
rect 568684 314608 568854 314664
rect 568910 314608 568915 314664
rect 568684 314606 568915 314608
rect 568684 314604 568690 314606
rect 568849 314603 568915 314606
rect 302877 313986 302943 313989
rect 305177 313986 305243 313989
rect 302877 313984 305243 313986
rect 302877 313928 302882 313984
rect 302938 313928 305182 313984
rect 305238 313928 305243 313984
rect 302877 313926 305243 313928
rect 302877 313923 302943 313926
rect 305177 313923 305243 313926
rect 566038 313924 566044 313988
rect 566108 313986 566114 313988
rect 566457 313986 566523 313989
rect 566108 313984 566523 313986
rect 566108 313928 566462 313984
rect 566518 313928 566523 313984
rect 566108 313926 566523 313928
rect 566108 313924 566114 313926
rect 566457 313923 566523 313926
rect 583520 311932 584960 312172
rect 299238 307668 299244 307732
rect 299308 307730 299314 307732
rect 303061 307730 303127 307733
rect 299308 307728 303127 307730
rect 299308 307672 303066 307728
rect 303122 307672 303127 307728
rect 299308 307670 303127 307672
rect 299308 307668 299314 307670
rect 303061 307667 303127 307670
rect -960 306084 480 306324
rect 285438 305628 285444 305692
rect 285508 305690 285514 305692
rect 291469 305690 291535 305693
rect 285508 305688 291535 305690
rect 285508 305632 291474 305688
rect 291530 305632 291535 305688
rect 285508 305630 291535 305632
rect 285508 305628 285514 305630
rect 291469 305627 291535 305630
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 291469 206002 291535 206005
rect 287010 206000 291535 206002
rect 287010 205944 291474 206000
rect 291530 205944 291535 206000
rect 287010 205942 291535 205944
rect 20478 205804 20484 205868
rect 20548 205866 20554 205868
rect 23841 205866 23907 205869
rect 20548 205864 23907 205866
rect 20548 205808 23846 205864
rect 23902 205808 23907 205864
rect 20548 205806 23907 205808
rect 20548 205804 20554 205806
rect 23841 205803 23907 205806
rect 285765 205866 285831 205869
rect 287010 205866 287070 205942
rect 291469 205939 291535 205942
rect 299238 205940 299244 206004
rect 299308 206002 299314 206004
rect 299308 205942 303722 206002
rect 299308 205940 299314 205942
rect 285765 205864 287070 205866
rect 285765 205808 285770 205864
rect 285826 205808 287070 205864
rect 285765 205806 287070 205808
rect 303662 205866 303722 205942
rect 303797 205866 303863 205869
rect 303662 205864 303863 205866
rect 303662 205808 303802 205864
rect 303858 205808 303863 205864
rect 303662 205806 303863 205808
rect 285765 205803 285831 205806
rect 303797 205803 303863 205806
rect 565721 205866 565787 205869
rect 572897 205866 572963 205869
rect 565721 205864 572963 205866
rect 565721 205808 565726 205864
rect 565782 205808 572902 205864
rect 572958 205808 572963 205864
rect 565721 205806 572963 205808
rect 565721 205803 565787 205806
rect 572897 205803 572963 205806
rect 21766 205668 21772 205732
rect 21836 205730 21842 205732
rect 23749 205730 23815 205733
rect 21836 205728 23815 205730
rect 21836 205672 23754 205728
rect 23810 205672 23815 205728
rect 21836 205670 23815 205672
rect 21836 205668 21842 205670
rect 23749 205667 23815 205670
rect 284937 205730 285003 205733
rect 294045 205730 294111 205733
rect 284937 205728 294111 205730
rect 284937 205672 284942 205728
rect 284998 205672 294050 205728
rect 294106 205672 294111 205728
rect 284937 205670 294111 205672
rect 284937 205667 285003 205670
rect 294045 205667 294111 205670
rect 301630 205668 301636 205732
rect 301700 205730 301706 205732
rect 303705 205730 303771 205733
rect 301700 205728 303771 205730
rect 301700 205672 303710 205728
rect 303766 205672 303771 205728
rect 301700 205670 303771 205672
rect 301700 205668 301706 205670
rect 303705 205667 303771 205670
rect 303521 205596 303587 205597
rect 303470 205532 303476 205596
rect 303540 205594 303587 205596
rect 564433 205594 564499 205597
rect 568849 205594 568915 205597
rect 303540 205592 303632 205594
rect 303582 205536 303632 205592
rect 303540 205534 303632 205536
rect 564433 205592 568915 205594
rect 564433 205536 564438 205592
rect 564494 205536 568854 205592
rect 568910 205536 568915 205592
rect 583520 205580 584960 205820
rect 564433 205534 568915 205536
rect 303540 205532 303587 205534
rect 303521 205531 303587 205532
rect 564433 205531 564499 205534
rect 568849 205531 568915 205534
rect 297909 205050 297975 205053
rect 305177 205050 305243 205053
rect 297909 205048 305243 205050
rect 297909 204992 297914 205048
rect 297970 204992 305182 205048
rect 305238 204992 305243 205048
rect 297909 204990 305243 204992
rect 297909 204987 297975 204990
rect 305177 204987 305243 204990
rect 286961 204914 287027 204917
rect 301446 204914 301452 204916
rect 286961 204912 301452 204914
rect 286961 204856 286966 204912
rect 287022 204856 301452 204912
rect 286961 204854 301452 204856
rect 286961 204851 287027 204854
rect 301446 204852 301452 204854
rect 301516 204852 301522 204916
rect 450169 204370 450235 204373
rect 568021 204370 568087 204373
rect 450169 204368 568087 204370
rect 450169 204312 450174 204368
rect 450230 204312 568026 204368
rect 568082 204312 568087 204368
rect 450169 204310 568087 204312
rect 450169 204307 450235 204310
rect 568021 204307 568087 204310
rect 19558 204172 19564 204236
rect 19628 204234 19634 204236
rect 20345 204234 20411 204237
rect 19628 204232 20411 204234
rect 19628 204176 20350 204232
rect 20406 204176 20411 204232
rect 19628 204174 20411 204176
rect 19628 204172 19634 204174
rect 20345 204171 20411 204174
rect 21214 204172 21220 204236
rect 21284 204234 21290 204236
rect 22001 204234 22067 204237
rect 21284 204232 22067 204234
rect 21284 204176 22006 204232
rect 22062 204176 22067 204232
rect 21284 204174 22067 204176
rect 21284 204172 21290 204174
rect 22001 204171 22067 204174
rect 22185 204234 22251 204237
rect 94037 204234 94103 204237
rect 22185 204232 94103 204234
rect 22185 204176 22190 204232
rect 22246 204176 94042 204232
rect 94098 204176 94103 204232
rect 22185 204174 94103 204176
rect 22185 204171 22251 204174
rect 94037 204171 94103 204174
rect 308489 204234 308555 204237
rect 580441 204234 580507 204237
rect 308489 204232 580507 204234
rect 308489 204176 308494 204232
rect 308550 204176 580446 204232
rect 580502 204176 580507 204232
rect 308489 204174 580507 204176
rect 308489 204171 308555 204174
rect 580441 204171 580507 204174
rect 3417 204098 3483 204101
rect 28165 204098 28231 204101
rect 3417 204096 28231 204098
rect 3417 204040 3422 204096
rect 3478 204040 28170 204096
rect 28226 204040 28231 204096
rect 3417 204038 28231 204040
rect 3417 204035 3483 204038
rect 28165 204035 28231 204038
rect 536189 204098 536255 204101
rect 568573 204098 568639 204101
rect 536189 204096 568639 204098
rect 536189 204040 536194 204096
rect 536250 204040 568578 204096
rect 568634 204040 568639 204096
rect 536189 204038 568639 204040
rect 536189 204035 536255 204038
rect 568573 204035 568639 204038
rect 19333 203962 19399 203965
rect 22185 203962 22251 203965
rect 19333 203960 22251 203962
rect 19333 203904 19338 203960
rect 19394 203904 22190 203960
rect 22246 203904 22251 203960
rect 19333 203902 22251 203904
rect 19333 203899 19399 203902
rect 22185 203899 22251 203902
rect 23013 203962 23079 203965
rect 23197 203962 23263 203965
rect 43345 203962 43411 203965
rect 23013 203960 43411 203962
rect 23013 203904 23018 203960
rect 23074 203904 23202 203960
rect 23258 203904 43350 203960
rect 43406 203904 43411 203960
rect 23013 203902 43411 203904
rect 23013 203899 23079 203902
rect 23197 203899 23263 203902
rect 43345 203899 43411 203902
rect 285673 203690 285739 203693
rect 286726 203690 286732 203692
rect 285673 203688 286732 203690
rect 285673 203632 285678 203688
rect 285734 203632 286732 203688
rect 285673 203630 286732 203632
rect 285673 203627 285739 203630
rect 286726 203628 286732 203630
rect 286796 203690 286802 203692
rect 289997 203690 290063 203693
rect 286796 203688 290063 203690
rect 286796 203632 290002 203688
rect 290058 203632 290063 203688
rect 286796 203630 290063 203632
rect 286796 203628 286802 203630
rect 289997 203627 290063 203630
rect 271689 203554 271755 203557
rect 301497 203554 301563 203557
rect 271689 203552 301563 203554
rect 271689 203496 271694 203552
rect 271750 203496 301502 203552
rect 301558 203496 301563 203552
rect 271689 203494 301563 203496
rect 271689 203491 271755 203494
rect 301497 203491 301563 203494
rect 301630 203492 301636 203556
rect 301700 203554 301706 203556
rect 485589 203554 485655 203557
rect 301700 203552 485655 203554
rect 301700 203496 485594 203552
rect 485650 203496 485655 203552
rect 301700 203494 485655 203496
rect 301700 203492 301706 203494
rect 485589 203491 485655 203494
rect 20621 202874 20687 202877
rect 22737 202874 22803 202877
rect 68645 202874 68711 202877
rect 20621 202872 68711 202874
rect 20621 202816 20626 202872
rect 20682 202816 22742 202872
rect 22798 202816 68650 202872
rect 68706 202816 68711 202872
rect 20621 202814 68711 202816
rect 20621 202811 20687 202814
rect 22737 202811 22803 202814
rect 68645 202811 68711 202814
rect 22921 202740 22987 202741
rect 22870 202738 22876 202740
rect 22830 202678 22876 202738
rect 22940 202736 22987 202740
rect 22982 202680 22987 202736
rect 22870 202676 22876 202678
rect 22940 202676 22987 202680
rect 22921 202675 22987 202676
rect 23238 202132 23244 202196
rect 23308 202194 23314 202196
rect 24853 202194 24919 202197
rect 96613 202194 96679 202197
rect 23308 202192 96679 202194
rect 23308 202136 24858 202192
rect 24914 202136 96618 202192
rect 96674 202136 96679 202192
rect 23308 202134 96679 202136
rect 23308 202132 23314 202134
rect 24853 202131 24919 202134
rect 96613 202131 96679 202134
rect -960 201772 480 202012
rect 570321 201380 570387 201381
rect 570270 201378 570276 201380
rect 570230 201318 570276 201378
rect 570340 201376 570387 201380
rect 570382 201320 570387 201376
rect 570270 201316 570276 201318
rect 570340 201316 570387 201320
rect 570321 201315 570387 201316
rect 298686 201180 298692 201244
rect 298756 201242 298762 201244
rect 299197 201242 299263 201245
rect 298756 201240 299263 201242
rect 298756 201184 299202 201240
rect 299258 201184 299263 201240
rect 298756 201182 299263 201184
rect 298756 201180 298762 201182
rect 299197 201179 299263 201182
rect 298870 200636 298876 200700
rect 298940 200698 298946 200700
rect 480529 200698 480595 200701
rect 298940 200696 480595 200698
rect 298940 200640 480534 200696
rect 480590 200640 480595 200696
rect 298940 200638 480595 200640
rect 298940 200636 298946 200638
rect 480529 200635 480595 200638
rect 17125 199202 17191 199205
rect 17718 199202 17724 199204
rect 17125 199200 17724 199202
rect 17125 199144 17130 199200
rect 17186 199144 17724 199200
rect 17125 199142 17724 199144
rect 17125 199139 17191 199142
rect 17718 199140 17724 199142
rect 17788 199140 17794 199204
rect 583520 192388 584960 192628
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 204253 188322 204319 188325
rect 285254 188322 285260 188324
rect 204253 188320 285260 188322
rect 204253 188264 204258 188320
rect 204314 188264 285260 188320
rect 204253 188262 285260 188264
rect 204253 188259 204319 188262
rect 285254 188260 285260 188262
rect 285324 188260 285330 188324
rect 303470 188260 303476 188324
rect 303540 188322 303546 188324
rect 569166 188322 569172 188324
rect 303540 188262 569172 188322
rect 303540 188260 303546 188262
rect 569166 188260 569172 188262
rect 569236 188260 569242 188324
rect 301998 187580 302004 187644
rect 302068 187642 302074 187644
rect 305177 187642 305243 187645
rect 305729 187642 305795 187645
rect 302068 187640 305795 187642
rect 302068 187584 305182 187640
rect 305238 187584 305734 187640
rect 305790 187584 305795 187640
rect 302068 187582 305795 187584
rect 302068 187580 302074 187582
rect 305177 187579 305243 187582
rect 305729 187579 305795 187582
rect 564341 187642 564407 187645
rect 568614 187642 568620 187644
rect 564341 187640 568620 187642
rect 564341 187584 564346 187640
rect 564402 187584 568620 187640
rect 564341 187582 568620 187584
rect 564341 187579 564407 187582
rect 568614 187580 568620 187582
rect 568684 187580 568690 187644
rect 23054 186356 23060 186420
rect 23124 186418 23130 186420
rect 24853 186418 24919 186421
rect 23124 186416 24919 186418
rect 23124 186360 24858 186416
rect 24914 186360 24919 186416
rect 23124 186358 24919 186360
rect 23124 186356 23130 186358
rect 24853 186355 24919 186358
rect 286174 186084 286180 186148
rect 286244 186146 286250 186148
rect 286961 186146 287027 186149
rect 286244 186144 287027 186146
rect 286244 186088 286966 186144
rect 287022 186088 287027 186144
rect 286244 186086 287027 186088
rect 286244 186084 286250 186086
rect 286961 186083 287027 186086
rect 17401 186010 17467 186013
rect 21766 186010 21772 186012
rect 17401 186008 21772 186010
rect 17401 185952 17406 186008
rect 17462 185952 21772 186008
rect 17401 185950 21772 185952
rect 17401 185947 17467 185950
rect 21766 185948 21772 185950
rect 21836 186010 21842 186012
rect 124213 186010 124279 186013
rect 21836 186008 124279 186010
rect 21836 185952 124218 186008
rect 124274 185952 124279 186008
rect 21836 185950 124279 185952
rect 21836 185948 21842 185950
rect 124213 185947 124279 185950
rect 284937 186010 285003 186013
rect 295333 186010 295399 186013
rect 284937 186008 295399 186010
rect 284937 185952 284942 186008
rect 284998 185952 295338 186008
rect 295394 185952 295399 186008
rect 284937 185950 295399 185952
rect 284937 185947 285003 185950
rect 295333 185947 295399 185950
rect 285121 185874 285187 185877
rect 291469 185874 291535 185877
rect 285121 185872 291535 185874
rect 285121 185816 285126 185872
rect 285182 185816 291474 185872
rect 291530 185816 291535 185872
rect 285121 185814 291535 185816
rect 285121 185811 285187 185814
rect 291469 185811 291535 185814
rect 298686 185812 298692 185876
rect 298756 185874 298762 185876
rect 303613 185874 303679 185877
rect 298756 185872 303679 185874
rect 298756 185816 303618 185872
rect 303674 185816 303679 185872
rect 298756 185814 303679 185816
rect 298756 185812 298762 185814
rect 303613 185811 303679 185814
rect 583520 179060 584960 179300
rect 285254 177924 285260 177988
rect 285324 177986 285330 177988
rect 288617 177986 288683 177989
rect 285324 177984 288683 177986
rect 285324 177928 288622 177984
rect 288678 177928 288683 177984
rect 285324 177926 288683 177928
rect 285324 177924 285330 177926
rect 288617 177923 288683 177926
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 2957 149834 3023 149837
rect -960 149832 3023 149834
rect -960 149776 2962 149832
rect 3018 149776 3023 149832
rect -960 149774 3023 149776
rect -960 149684 480 149774
rect 2957 149771 3023 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 565302 79324 565308 79388
rect 565372 79386 565378 79388
rect 570229 79386 570295 79389
rect 565372 79384 570295 79386
rect 565372 79328 570234 79384
rect 570290 79328 570295 79384
rect 565372 79326 570295 79328
rect 565372 79324 565378 79326
rect 570229 79323 570295 79326
rect 21766 77828 21772 77892
rect 21836 77890 21842 77892
rect 25589 77890 25655 77893
rect 21836 77888 25655 77890
rect 21836 77832 25594 77888
rect 25650 77832 25655 77888
rect 21836 77830 25655 77832
rect 21836 77828 21842 77830
rect 25589 77827 25655 77830
rect 194593 77890 194659 77893
rect 195789 77890 195855 77893
rect 295333 77890 295399 77893
rect 303521 77892 303587 77893
rect 194593 77888 295399 77890
rect 194593 77832 194598 77888
rect 194654 77832 195794 77888
rect 195850 77832 295338 77888
rect 295394 77832 295399 77888
rect 194593 77830 295399 77832
rect 194593 77827 194659 77830
rect 195789 77827 195855 77830
rect 295333 77827 295399 77830
rect 303470 77828 303476 77892
rect 303540 77890 303587 77892
rect 336733 77890 336799 77893
rect 303540 77888 303632 77890
rect 303582 77832 303632 77888
rect 303540 77830 303632 77832
rect 306330 77888 336799 77890
rect 306330 77832 336738 77888
rect 336794 77832 336799 77888
rect 306330 77830 336799 77832
rect 303540 77828 303587 77830
rect 303521 77827 303587 77828
rect 284293 77754 284359 77757
rect 291469 77754 291535 77757
rect 284293 77752 291535 77754
rect 284293 77696 284298 77752
rect 284354 77696 291474 77752
rect 291530 77696 291535 77752
rect 284293 77694 291535 77696
rect 284293 77691 284359 77694
rect 291469 77691 291535 77694
rect 301998 77692 302004 77756
rect 302068 77754 302074 77756
rect 306330 77754 306390 77830
rect 336733 77827 336799 77830
rect 454033 77890 454099 77893
rect 455321 77890 455387 77893
rect 568614 77890 568620 77892
rect 454033 77888 568620 77890
rect 454033 77832 454038 77888
rect 454094 77832 455326 77888
rect 455382 77832 568620 77888
rect 454033 77830 568620 77832
rect 454033 77827 454099 77830
rect 455321 77827 455387 77830
rect 568614 77828 568620 77830
rect 568684 77828 568690 77892
rect 302068 77694 306390 77754
rect 302068 77692 302074 77694
rect 52453 77074 52519 77077
rect 53787 77074 53853 77077
rect 52453 77072 53853 77074
rect 52453 77016 52458 77072
rect 52514 77016 53792 77072
rect 53848 77016 53853 77072
rect 52453 77014 53853 77016
rect 52453 77011 52519 77014
rect 53787 77011 53853 77014
rect 297173 76938 297239 76941
rect 297950 76938 297956 76940
rect 297173 76936 297956 76938
rect 297173 76880 297178 76936
rect 297234 76880 297956 76936
rect 297173 76878 297956 76880
rect 297173 76875 297239 76878
rect 297950 76876 297956 76878
rect 298020 76876 298026 76940
rect 282177 76802 282243 76805
rect 295006 76802 295012 76804
rect 282177 76800 295012 76802
rect 282177 76744 282182 76800
rect 282238 76744 295012 76800
rect 282177 76742 295012 76744
rect 282177 76739 282243 76742
rect 295006 76740 295012 76742
rect 295076 76740 295082 76804
rect 302734 76740 302740 76804
rect 302804 76802 302810 76804
rect 398833 76802 398899 76805
rect 302804 76800 398899 76802
rect 302804 76744 398838 76800
rect 398894 76744 398899 76800
rect 302804 76742 398899 76744
rect 302804 76740 302810 76742
rect 398833 76739 398899 76742
rect 224953 76666 225019 76669
rect 301630 76666 301636 76668
rect 224953 76664 301636 76666
rect 224953 76608 224958 76664
rect 225014 76608 301636 76664
rect 224953 76606 301636 76608
rect 224953 76603 225019 76606
rect 301630 76604 301636 76606
rect 301700 76604 301706 76668
rect 386413 76666 386479 76669
rect 567326 76666 567332 76668
rect 386413 76664 567332 76666
rect 386413 76608 386418 76664
rect 386474 76608 567332 76664
rect 386413 76606 567332 76608
rect 386413 76603 386479 76606
rect 567326 76604 567332 76606
rect 567396 76604 567402 76668
rect 151721 76530 151787 76533
rect 287646 76530 287652 76532
rect 151721 76528 287652 76530
rect 151721 76472 151726 76528
rect 151782 76472 287652 76528
rect 151721 76470 287652 76472
rect 151721 76467 151787 76470
rect 287646 76468 287652 76470
rect 287716 76468 287722 76532
rect 387793 76530 387859 76533
rect 569902 76530 569908 76532
rect 387793 76528 569908 76530
rect 387793 76472 387798 76528
rect 387854 76472 569908 76528
rect 387793 76470 569908 76472
rect 387793 76467 387859 76470
rect 569902 76468 569908 76470
rect 569972 76468 569978 76532
rect 574185 76530 574251 76533
rect 575238 76530 575244 76532
rect 574185 76528 575244 76530
rect 574185 76472 574190 76528
rect 574246 76472 575244 76528
rect 574185 76470 575244 76472
rect 574185 76467 574251 76470
rect 575238 76468 575244 76470
rect 575308 76468 575314 76532
rect 291469 76394 291535 76397
rect 292430 76394 292436 76396
rect 291469 76392 292436 76394
rect 291469 76336 291474 76392
rect 291530 76336 292436 76392
rect 291469 76334 292436 76336
rect 291469 76331 291535 76334
rect 292430 76332 292436 76334
rect 292500 76332 292506 76396
rect 571425 76124 571491 76125
rect 571374 76060 571380 76124
rect 571444 76122 571491 76124
rect 571444 76120 571536 76122
rect 571486 76064 571536 76120
rect 571444 76062 571536 76064
rect 571444 76060 571491 76062
rect 571425 76059 571491 76060
rect 22870 75924 22876 75988
rect 22940 75986 22946 75988
rect 52453 75986 52519 75989
rect 22940 75984 52519 75986
rect 22940 75928 52458 75984
rect 52514 75928 52519 75984
rect 22940 75926 52519 75928
rect 22940 75924 22946 75926
rect 52453 75923 52519 75926
rect 23054 75788 23060 75852
rect 23124 75850 23130 75852
rect 98637 75850 98703 75853
rect 23124 75848 98703 75850
rect 23124 75792 98642 75848
rect 98698 75792 98703 75848
rect 23124 75790 98703 75792
rect 23124 75788 23130 75790
rect 98637 75787 98703 75790
rect 308489 75850 308555 75853
rect 577589 75850 577655 75853
rect 308489 75848 577655 75850
rect 308489 75792 308494 75848
rect 308550 75792 577594 75848
rect 577650 75792 577655 75848
rect 308489 75790 577655 75792
rect 308489 75787 308555 75790
rect 577589 75787 577655 75790
rect 21950 75652 21956 75716
rect 22020 75714 22026 75716
rect 84101 75714 84167 75717
rect 22020 75712 84167 75714
rect 22020 75656 84106 75712
rect 84162 75656 84167 75712
rect 22020 75654 84167 75656
rect 22020 75652 22026 75654
rect 84101 75651 84167 75654
rect 19558 75516 19564 75580
rect 19628 75578 19634 75580
rect 79409 75578 79475 75581
rect 19628 75576 79475 75578
rect 19628 75520 79414 75576
rect 79470 75520 79475 75576
rect 19628 75518 79475 75520
rect 19628 75516 19634 75518
rect 79409 75515 79475 75518
rect 233233 75170 233299 75173
rect 505829 75170 505895 75173
rect 233233 75168 505895 75170
rect 233233 75112 233238 75168
rect 233294 75112 505834 75168
rect 505890 75112 505895 75168
rect 233233 75110 505895 75112
rect 233233 75107 233299 75110
rect 505829 75107 505895 75110
rect 17585 74490 17651 74493
rect 104157 74490 104223 74493
rect 17585 74488 104223 74490
rect 17585 74432 17590 74488
rect 17646 74432 104162 74488
rect 104218 74432 104223 74488
rect 17585 74430 104223 74432
rect 17585 74427 17651 74430
rect 104157 74427 104223 74430
rect 282269 73946 282335 73949
rect 298870 73946 298876 73948
rect 282269 73944 298876 73946
rect 282269 73888 282274 73944
rect 282330 73888 298876 73944
rect 282269 73886 298876 73888
rect 282269 73883 282335 73886
rect 298870 73884 298876 73886
rect 298940 73884 298946 73948
rect 407113 73946 407179 73949
rect 569953 73946 570019 73949
rect 407113 73944 570019 73946
rect 407113 73888 407118 73944
rect 407174 73888 569958 73944
rect 570014 73888 570019 73944
rect 407113 73886 570019 73888
rect 407113 73883 407179 73886
rect 569953 73883 570019 73886
rect 204345 73810 204411 73813
rect 296110 73810 296116 73812
rect 204345 73808 296116 73810
rect 204345 73752 204350 73808
rect 204406 73752 296116 73808
rect 204345 73750 296116 73752
rect 204345 73747 204411 73750
rect 296110 73748 296116 73750
rect 296180 73748 296186 73812
rect 403065 73810 403131 73813
rect 571333 73810 571399 73813
rect 403065 73808 571399 73810
rect 403065 73752 403070 73808
rect 403126 73752 571338 73808
rect 571394 73752 571399 73808
rect 403065 73750 571399 73752
rect 403065 73747 403131 73750
rect 571333 73747 571399 73750
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 17718 71708 17724 71772
rect 17788 71770 17794 71772
rect 128997 71770 129063 71773
rect 17788 71768 129063 71770
rect 17788 71712 129002 71768
rect 129058 71712 129063 71768
rect 17788 71710 129063 71712
rect 17788 71708 17794 71710
rect 128997 71707 129063 71710
rect 465717 71770 465783 71773
rect 570086 71770 570092 71772
rect 465717 71768 570092 71770
rect 465717 71712 465722 71768
rect 465778 71712 570092 71768
rect 465717 71710 570092 71712
rect 465717 71707 465783 71710
rect 570086 71708 570092 71710
rect 570156 71708 570162 71772
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 558177 69730 558243 69733
rect 566038 69730 566044 69732
rect 558177 69728 566044 69730
rect 558177 69672 558182 69728
rect 558238 69672 566044 69728
rect 558177 69670 566044 69672
rect 558177 69667 558243 69670
rect 566038 69668 566044 69670
rect 566108 69668 566114 69732
rect 420177 68914 420243 68917
rect 565302 68914 565308 68916
rect 420177 68912 565308 68914
rect 420177 68856 420182 68912
rect 420238 68856 565308 68912
rect 420177 68854 565308 68856
rect 420177 68851 420243 68854
rect 565302 68852 565308 68854
rect 565372 68852 565378 68916
rect 198825 68234 198891 68237
rect 298686 68234 298692 68236
rect 198825 68232 298692 68234
rect 198825 68176 198830 68232
rect 198886 68176 298692 68232
rect 198825 68174 298692 68176
rect 198825 68171 198891 68174
rect 298686 68172 298692 68174
rect 298756 68172 298762 68236
rect 439497 62794 439563 62797
rect 565854 62794 565860 62796
rect 439497 62792 565860 62794
rect 439497 62736 439502 62792
rect 439558 62736 565860 62792
rect 439497 62734 565860 62736
rect 439497 62731 439563 62734
rect 565854 62732 565860 62734
rect 565924 62732 565930 62796
rect 217225 59938 217291 59941
rect 292798 59938 292804 59940
rect 217225 59936 292804 59938
rect 217225 59880 217230 59936
rect 217286 59880 292804 59936
rect 217225 59878 292804 59880
rect 217225 59875 217291 59878
rect 292798 59876 292804 59878
rect 292868 59876 292874 59940
rect 295926 59876 295932 59940
rect 295996 59938 296002 59940
rect 401593 59938 401659 59941
rect 295996 59936 401659 59938
rect 295996 59880 401598 59936
rect 401654 59880 401659 59936
rect 295996 59878 401659 59880
rect 295996 59876 296002 59878
rect 401593 59875 401659 59878
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 215753 57490 215819 57493
rect 291142 57490 291148 57492
rect 215753 57488 291148 57490
rect 215753 57432 215758 57488
rect 215814 57432 291148 57488
rect 215753 57430 291148 57432
rect 215753 57427 215819 57430
rect 291142 57428 291148 57430
rect 291212 57428 291218 57492
rect 213913 57354 213979 57357
rect 290038 57354 290044 57356
rect 213913 57352 290044 57354
rect 213913 57296 213918 57352
rect 213974 57296 290044 57352
rect 213913 57294 290044 57296
rect 213913 57291 213979 57294
rect 290038 57292 290044 57294
rect 290108 57292 290114 57356
rect 297766 57292 297772 57356
rect 297836 57354 297842 57356
rect 381353 57354 381419 57357
rect 297836 57352 381419 57354
rect 297836 57296 381358 57352
rect 381414 57296 381419 57352
rect 297836 57294 381419 57296
rect 297836 57292 297842 57294
rect 381353 57291 381419 57294
rect 286910 57156 286916 57220
rect 286980 57218 286986 57220
rect 419993 57218 420059 57221
rect 286980 57216 420059 57218
rect 286980 57160 419998 57216
rect 420054 57160 420059 57216
rect 286980 57158 420059 57160
rect 286980 57156 286986 57158
rect 419993 57155 420059 57158
rect 287605 54906 287671 54909
rect 288198 54906 288204 54908
rect 287605 54904 288204 54906
rect 287605 54848 287610 54904
rect 287666 54848 288204 54904
rect 287605 54846 288204 54848
rect 287605 54843 287671 54846
rect 288198 54844 288204 54846
rect 288268 54844 288274 54908
rect 280153 54770 280219 54773
rect 292614 54770 292620 54772
rect 280153 54768 292620 54770
rect 280153 54712 280158 54768
rect 280214 54712 292620 54768
rect 280153 54710 292620 54712
rect 280153 54707 280219 54710
rect 292614 54708 292620 54710
rect 292684 54708 292690 54772
rect 276473 54634 276539 54637
rect 289854 54634 289860 54636
rect 276473 54632 289860 54634
rect 276473 54576 276478 54632
rect 276534 54576 289860 54632
rect 276473 54574 289860 54576
rect 276473 54571 276539 54574
rect 289854 54572 289860 54574
rect 289924 54572 289930 54636
rect 299974 54572 299980 54636
rect 300044 54634 300050 54636
rect 421833 54634 421899 54637
rect 300044 54632 421899 54634
rect 300044 54576 421838 54632
rect 421894 54576 421899 54632
rect 300044 54574 421899 54576
rect 300044 54572 300050 54574
rect 421833 54571 421899 54574
rect 202873 54498 202939 54501
rect 282177 54498 282243 54501
rect 202873 54496 282243 54498
rect 202873 54440 202878 54496
rect 202934 54440 282182 54496
rect 282238 54440 282243 54496
rect 202873 54438 282243 54440
rect 202873 54435 202939 54438
rect 282177 54435 282243 54438
rect 283833 54498 283899 54501
rect 289118 54498 289124 54500
rect 283833 54496 289124 54498
rect 283833 54440 283838 54496
rect 283894 54440 289124 54496
rect 283833 54438 289124 54440
rect 283833 54435 283899 54438
rect 289118 54436 289124 54438
rect 289188 54436 289194 54500
rect 300158 54436 300164 54500
rect 300228 54498 300234 54500
rect 423673 54498 423739 54501
rect 300228 54496 423739 54498
rect 300228 54440 423678 54496
rect 423734 54440 423739 54496
rect 300228 54438 423739 54440
rect 300228 54436 300234 54438
rect 423673 54435 423739 54438
rect 425513 54498 425579 54501
rect 566958 54498 566964 54500
rect 425513 54496 566964 54498
rect 425513 54440 425518 54496
rect 425574 54440 566964 54496
rect 425513 54438 566964 54440
rect 425513 54435 425579 54438
rect 566958 54436 566964 54438
rect 567028 54436 567034 54500
rect 285765 53954 285831 53957
rect 286174 53954 286180 53956
rect 285765 53952 286180 53954
rect 285765 53896 285770 53952
rect 285826 53896 286180 53952
rect 285765 53894 286180 53896
rect 285765 53891 285831 53894
rect 286174 53892 286180 53894
rect 286244 53892 286250 53956
rect 151629 53138 151695 53141
rect 288934 53138 288940 53140
rect 151629 53136 288940 53138
rect 151629 53080 151634 53136
rect 151690 53080 288940 53136
rect 151629 53078 288940 53080
rect 151629 53075 151695 53078
rect 288934 53076 288940 53078
rect 289004 53076 289010 53140
rect 150433 50554 150499 50557
rect 150433 50552 153394 50554
rect 150433 50496 150438 50552
rect 150494 50496 153394 50552
rect 150433 50494 153394 50496
rect 150433 50491 150499 50494
rect 153334 49912 153394 50494
rect 150433 49602 150499 49605
rect 150433 49600 153394 49602
rect 150433 49544 150438 49600
rect 150494 49544 153394 49600
rect 150433 49542 153394 49544
rect 150433 49539 150499 49542
rect 153334 48960 153394 49542
rect 150433 48242 150499 48245
rect 150433 48240 153394 48242
rect 150433 48184 150438 48240
rect 150494 48184 153394 48240
rect 150433 48182 153394 48184
rect 150433 48179 150499 48182
rect 153334 48008 153394 48182
rect 150525 47698 150591 47701
rect 150525 47696 153394 47698
rect 150525 47640 150530 47696
rect 150586 47640 153394 47696
rect 150525 47638 153394 47640
rect 150525 47635 150591 47638
rect 153334 47056 153394 47638
rect 150433 46746 150499 46749
rect 150433 46744 153394 46746
rect 150433 46688 150438 46744
rect 150494 46688 153394 46744
rect 150433 46686 153394 46688
rect 150433 46683 150499 46686
rect 153334 46104 153394 46686
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 151077 45522 151143 45525
rect 151077 45520 153394 45522
rect 151077 45464 151082 45520
rect 151138 45464 153394 45520
rect 151077 45462 153394 45464
rect 151077 45459 151143 45462
rect 153334 45152 153394 45462
rect 150433 44842 150499 44845
rect 150433 44840 153394 44842
rect 150433 44784 150438 44840
rect 150494 44784 153394 44840
rect 150433 44782 153394 44784
rect 150433 44779 150499 44782
rect 153334 44200 153394 44782
rect 150433 43890 150499 43893
rect 150433 43888 153394 43890
rect 150433 43832 150438 43888
rect 150494 43832 153394 43888
rect 150433 43830 153394 43832
rect 150433 43827 150499 43830
rect 153334 43248 153394 43830
rect 150433 42530 150499 42533
rect 150433 42528 153394 42530
rect 150433 42472 150438 42528
rect 150494 42472 153394 42528
rect 150433 42470 153394 42472
rect 150433 42467 150499 42470
rect 153334 42296 153394 42470
rect 150433 41306 150499 41309
rect 153334 41306 153394 41344
rect 150433 41304 153394 41306
rect 150433 41248 150438 41304
rect 150494 41248 153394 41304
rect 150433 41246 153394 41248
rect 150433 41243 150499 41246
rect 153009 40422 153075 40425
rect 153009 40420 153364 40422
rect 153009 40364 153014 40420
rect 153070 40364 153364 40420
rect 153009 40362 153364 40364
rect 153009 40359 153075 40362
rect 151537 39946 151603 39949
rect 151537 39944 153394 39946
rect 151537 39888 151542 39944
rect 151598 39888 153394 39944
rect 151537 39886 153394 39888
rect 151537 39883 151603 39886
rect 153334 39440 153394 39886
rect 153101 38722 153167 38725
rect 153101 38720 153394 38722
rect 153101 38664 153106 38720
rect 153162 38664 153394 38720
rect 153101 38662 153394 38664
rect 153101 38659 153167 38662
rect 153334 38488 153394 38662
rect 151721 38178 151787 38181
rect 151721 38176 153394 38178
rect 151721 38120 151726 38176
rect 151782 38120 153394 38176
rect 151721 38118 153394 38120
rect 151721 38115 151787 38118
rect 153334 37536 153394 38118
rect 434670 37634 434730 37944
rect 437381 37634 437447 37637
rect 434670 37632 437447 37634
rect 434670 37576 437386 37632
rect 437442 37576 437447 37632
rect 434670 37574 437447 37576
rect 437381 37571 437447 37574
rect 151629 37226 151695 37229
rect 151629 37224 153394 37226
rect 151629 37168 151634 37224
rect 151690 37168 153394 37224
rect 151629 37166 153394 37168
rect 151629 37163 151695 37166
rect 153334 36584 153394 37166
rect 150433 35866 150499 35869
rect 150433 35864 153394 35866
rect 150433 35808 150438 35864
rect 150494 35808 153394 35864
rect 150433 35806 153394 35808
rect 150433 35803 150499 35806
rect 153334 35632 153394 35806
rect 19190 34580 19196 34644
rect 19260 34642 19266 34644
rect 153334 34642 153394 34680
rect 19260 34582 153394 34642
rect 19260 34580 19266 34582
rect 150433 34370 150499 34373
rect 150433 34368 153394 34370
rect 150433 34312 150438 34368
rect 150494 34312 153394 34368
rect 150433 34310 153394 34312
rect 150433 34307 150499 34310
rect 153334 33728 153394 34310
rect 151169 33146 151235 33149
rect 151169 33144 153394 33146
rect 151169 33088 151174 33144
rect 151230 33088 153394 33144
rect 151169 33086 153394 33088
rect 151169 33083 151235 33086
rect 153334 32776 153394 33086
rect 583520 32996 584960 33236
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 150433 32466 150499 32469
rect 150433 32464 153394 32466
rect 150433 32408 150438 32464
rect 150494 32408 153394 32464
rect 150433 32406 153394 32408
rect 150433 32403 150499 32406
rect 153334 31824 153394 32406
rect 150433 31514 150499 31517
rect 150433 31512 153394 31514
rect 150433 31456 150438 31512
rect 150494 31456 153394 31512
rect 150433 31454 153394 31456
rect 150433 31451 150499 31454
rect 153334 30872 153394 31454
rect 150433 30154 150499 30157
rect 150433 30152 153394 30154
rect 150433 30096 150438 30152
rect 150494 30096 153394 30152
rect 150433 30094 153394 30096
rect 150433 30091 150499 30094
rect 153334 29920 153394 30094
rect 150433 28930 150499 28933
rect 153334 28930 153394 28968
rect 150433 28928 153394 28930
rect 150433 28872 150438 28928
rect 150494 28872 153394 28928
rect 150433 28870 153394 28872
rect 150433 28867 150499 28870
rect 151077 28522 151143 28525
rect 151077 28520 153394 28522
rect 151077 28464 151082 28520
rect 151138 28464 153394 28520
rect 151077 28462 153394 28464
rect 151077 28459 151143 28462
rect 153334 28016 153394 28462
rect 151077 26482 151143 26485
rect 153334 26482 153394 27064
rect 151077 26480 153394 26482
rect 151077 26424 151082 26480
rect 151138 26424 153394 26480
rect 151077 26422 153394 26424
rect 151077 26419 151143 26422
rect 150433 26210 150499 26213
rect 150433 26208 153394 26210
rect 150433 26152 150438 26208
rect 150494 26152 153394 26208
rect 150433 26150 153394 26152
rect 150433 26147 150499 26150
rect 153334 26112 153394 26150
rect 277301 23490 277367 23493
rect 518893 23490 518959 23493
rect 277301 23488 518959 23490
rect 277301 23432 277306 23488
rect 277362 23432 518898 23488
rect 518954 23432 518959 23488
rect 277301 23430 518959 23432
rect 277301 23427 277367 23430
rect 518893 23427 518959 23430
rect 281257 22130 281323 22133
rect 532693 22130 532759 22133
rect 281257 22128 532759 22130
rect 281257 22072 281262 22128
rect 281318 22072 532698 22128
rect 532754 22072 532759 22128
rect 281257 22070 532759 22072
rect 281257 22067 281323 22070
rect 532693 22067 532759 22070
rect 247677 21450 247743 21453
rect 299473 21450 299539 21453
rect 247677 21448 299539 21450
rect 247677 21392 247682 21448
rect 247738 21392 299478 21448
rect 299534 21392 299539 21448
rect 247677 21390 299539 21392
rect 247677 21387 247743 21390
rect 299473 21387 299539 21390
rect 276197 21314 276263 21317
rect 381721 21314 381787 21317
rect 276197 21312 381787 21314
rect 276197 21256 276202 21312
rect 276258 21256 381726 21312
rect 381782 21256 381787 21312
rect 276197 21254 381787 21256
rect 276197 21251 276263 21254
rect 381721 21251 381787 21254
rect 265065 19954 265131 19957
rect 476113 19954 476179 19957
rect 265065 19952 476179 19954
rect 265065 19896 265070 19952
rect 265126 19896 476118 19952
rect 476174 19896 476179 19952
rect 265065 19894 476179 19896
rect 265065 19891 265131 19894
rect 476113 19891 476179 19894
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 262029 18594 262095 18597
rect 465165 18594 465231 18597
rect 262029 18592 465231 18594
rect 262029 18536 262034 18592
rect 262090 18536 465170 18592
rect 465226 18536 465231 18592
rect 262029 18534 465231 18536
rect 262029 18531 262095 18534
rect 465165 18531 465231 18534
rect 289353 17370 289419 17373
rect 329097 17370 329163 17373
rect 289353 17368 329163 17370
rect 289353 17312 289358 17368
rect 289414 17312 329102 17368
rect 329158 17312 329163 17368
rect 289353 17310 329163 17312
rect 289353 17307 289419 17310
rect 329097 17307 329163 17310
rect 254945 17234 255011 17237
rect 440233 17234 440299 17237
rect 254945 17232 440299 17234
rect 254945 17176 254950 17232
rect 255006 17176 440238 17232
rect 440294 17176 440299 17232
rect 254945 17174 440299 17176
rect 254945 17171 255011 17174
rect 440233 17171 440299 17174
rect 256785 15874 256851 15877
rect 448605 15874 448671 15877
rect 256785 15872 448671 15874
rect 256785 15816 256790 15872
rect 256846 15816 448610 15872
rect 448666 15816 448671 15872
rect 256785 15814 448671 15816
rect 256785 15811 256851 15814
rect 448605 15811 448671 15814
rect 240133 14514 240199 14517
rect 384297 14514 384363 14517
rect 240133 14512 384363 14514
rect 240133 14456 240138 14512
rect 240194 14456 384302 14512
rect 384358 14456 384363 14512
rect 240133 14454 384363 14456
rect 240133 14451 240199 14454
rect 384297 14451 384363 14454
rect 163681 13018 163747 13021
rect 298737 13018 298803 13021
rect 163681 13016 298803 13018
rect 163681 12960 163686 13016
rect 163742 12960 298742 13016
rect 298798 12960 298803 13016
rect 163681 12958 298803 12960
rect 163681 12955 163747 12958
rect 298737 12955 298803 12958
rect 241973 11658 242039 11661
rect 398925 11658 398991 11661
rect 241973 11656 398991 11658
rect 241973 11600 241978 11656
rect 242034 11600 398930 11656
rect 398986 11600 398991 11656
rect 241973 11598 398991 11600
rect 241973 11595 242039 11598
rect 398925 11595 398991 11598
rect 226885 10298 226951 10301
rect 345289 10298 345355 10301
rect 226885 10296 345355 10298
rect 226885 10240 226890 10296
rect 226946 10240 345294 10296
rect 345350 10240 345355 10296
rect 226885 10238 345355 10240
rect 226885 10235 226951 10238
rect 345289 10235 345355 10238
rect 248413 9074 248479 9077
rect 420177 9074 420243 9077
rect 248413 9072 420243 9074
rect 248413 9016 248418 9072
rect 248474 9016 420182 9072
rect 420238 9016 420243 9072
rect 248413 9014 420243 9016
rect 248413 9011 248479 9014
rect 420177 9011 420243 9014
rect 291469 8938 291535 8941
rect 572713 8938 572779 8941
rect 291469 8936 572779 8938
rect 291469 8880 291474 8936
rect 291530 8880 572718 8936
rect 572774 8880 572779 8936
rect 291469 8878 572779 8880
rect 291469 8875 291535 8878
rect 572713 8875 572779 8878
rect 269205 7714 269271 7717
rect 293953 7714 294019 7717
rect 269205 7712 294019 7714
rect 269205 7656 269210 7712
rect 269266 7656 293958 7712
rect 294014 7656 294019 7712
rect 269205 7654 294019 7656
rect 269205 7651 269271 7654
rect 293953 7651 294019 7654
rect 287145 7578 287211 7581
rect 480253 7578 480319 7581
rect 287145 7576 480319 7578
rect 287145 7520 287150 7576
rect 287206 7520 480258 7576
rect 480314 7520 480319 7576
rect 287145 7518 480319 7520
rect 287145 7515 287211 7518
rect 480253 7515 480319 7518
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 255313 6354 255379 6357
rect 445017 6354 445083 6357
rect 255313 6352 445083 6354
rect 255313 6296 255318 6352
rect 255374 6296 445022 6352
rect 445078 6296 445083 6352
rect 255313 6294 445083 6296
rect 255313 6291 255379 6294
rect 445017 6291 445083 6294
rect 289813 6218 289879 6221
rect 565629 6218 565695 6221
rect 289813 6216 565695 6218
rect 289813 6160 289818 6216
rect 289874 6160 565634 6216
rect 565690 6160 565695 6216
rect 289813 6158 565695 6160
rect 289813 6155 289879 6158
rect 565629 6155 565695 6158
rect 271965 4994 272031 4997
rect 501781 4994 501847 4997
rect 271965 4992 501847 4994
rect 271965 4936 271970 4992
rect 272026 4936 501786 4992
rect 501842 4936 501847 4992
rect 271965 4934 501847 4936
rect 271965 4931 272031 4934
rect 501781 4931 501847 4934
rect 282913 4858 282979 4861
rect 540789 4858 540855 4861
rect 282913 4856 540855 4858
rect 282913 4800 282918 4856
rect 282974 4800 540794 4856
rect 540850 4800 540855 4856
rect 282913 4798 540855 4800
rect 282913 4795 282979 4798
rect 540789 4795 540855 4798
rect 280061 3498 280127 3501
rect 296069 3498 296135 3501
rect 280061 3496 296135 3498
rect 280061 3440 280066 3496
rect 280122 3440 296074 3496
rect 296130 3440 296135 3496
rect 280061 3438 296135 3440
rect 280061 3435 280127 3438
rect 296069 3435 296135 3438
rect 301497 3498 301563 3501
rect 303153 3498 303219 3501
rect 301497 3496 303219 3498
rect 301497 3440 301502 3496
rect 301558 3440 303158 3496
rect 303214 3440 303219 3496
rect 301497 3438 303219 3440
rect 301497 3435 301563 3438
rect 303153 3435 303219 3438
rect 156597 3362 156663 3365
rect 300485 3362 300551 3365
rect 156597 3360 300551 3362
rect 156597 3304 156602 3360
rect 156658 3304 300490 3360
rect 300546 3304 300551 3360
rect 156597 3302 300551 3304
rect 156597 3299 156663 3302
rect 300485 3299 300551 3302
rect 305637 3362 305703 3365
rect 313825 3362 313891 3365
rect 305637 3360 313891 3362
rect 305637 3304 305642 3360
rect 305698 3304 313830 3360
rect 313886 3304 313891 3360
rect 305637 3302 313891 3304
rect 305637 3299 305703 3302
rect 313825 3299 313891 3302
rect 287053 2002 287119 2005
rect 558545 2002 558611 2005
rect 287053 2000 558611 2002
rect 287053 1944 287058 2000
rect 287114 1944 558550 2000
rect 558606 1944 558611 2000
rect 287053 1942 558611 1944
rect 287053 1939 287119 1942
rect 558545 1939 558611 1942
<< via3 >>
rect 288940 700300 289004 700364
rect 19196 699816 19260 699820
rect 19196 699760 19246 699816
rect 19246 699760 19260 699816
rect 19196 699756 19260 699760
rect 287652 699756 287716 699820
rect 303476 697444 303540 697508
rect 575244 590956 575308 591020
rect 292620 585788 292684 585852
rect 297956 585788 298020 585852
rect 23244 585652 23308 585716
rect 292436 585652 292500 585716
rect 571380 585652 571444 585716
rect 286180 585108 286244 585172
rect 566964 585108 567028 585172
rect 565860 583068 565924 583132
rect 17724 582932 17788 582996
rect 285628 582932 285692 582996
rect 566044 582932 566108 582996
rect 567332 580348 567396 580412
rect 290044 580212 290108 580276
rect 301636 580212 301700 580276
rect 570092 580212 570156 580276
rect 295932 572052 295996 572116
rect 292804 571916 292868 571980
rect 302188 571916 302252 571980
rect 568620 571916 568684 571980
rect 21956 570556 22020 570620
rect 288204 570556 288268 570620
rect 286180 461952 286244 461956
rect 286180 461896 286230 461952
rect 286230 461896 286244 461952
rect 286180 461892 286244 461896
rect 303476 461952 303540 461956
rect 303476 461896 303526 461952
rect 303526 461896 303540 461952
rect 303476 461892 303540 461896
rect 302004 461756 302068 461820
rect 568620 460940 568684 461004
rect 21956 460260 22020 460324
rect 286180 460668 286244 460732
rect 570092 460260 570156 460324
rect 17724 460124 17788 460188
rect 290044 460124 290108 460188
rect 570092 460124 570156 460188
rect 289860 459580 289924 459644
rect 570092 459580 570156 459644
rect 301636 459444 301700 459508
rect 302740 459036 302804 459100
rect 565676 459036 565740 459100
rect 567332 459036 567396 459100
rect 299980 458900 300044 458964
rect 301452 458900 301516 458964
rect 295012 458764 295076 458828
rect 567332 458764 567396 458828
rect 568620 458628 568684 458692
rect 285444 458280 285508 458284
rect 285444 458224 285458 458280
rect 285458 458224 285508 458280
rect 285444 458220 285508 458224
rect 301636 458220 301700 458284
rect 23244 458084 23308 458148
rect 285628 458084 285692 458148
rect 565860 458144 565924 458148
rect 565860 458088 565910 458144
rect 565910 458088 565924 458144
rect 565860 458084 565924 458088
rect 566044 457404 566108 457468
rect 21956 456860 22020 456924
rect 23244 456860 23308 456924
rect 286364 456860 286428 456924
rect 23244 444212 23308 444276
rect 297772 443940 297836 444004
rect 290044 443804 290108 443868
rect 291148 443668 291212 443732
rect 298692 443668 298756 443732
rect 289124 443532 289188 443596
rect 298692 442852 298756 442916
rect 302004 442852 302068 442916
rect 566596 442852 566660 442916
rect 285444 433876 285508 433940
rect 565676 433332 565740 433396
rect 569172 418236 569236 418300
rect 286364 334052 286428 334116
rect 302004 334052 302068 334116
rect 570092 334596 570156 334660
rect 289860 332480 289924 332484
rect 289860 332424 289910 332480
rect 289910 332424 289924 332480
rect 289860 332420 289924 332424
rect 286180 332148 286244 332212
rect 301636 331876 301700 331940
rect 289860 331740 289924 331804
rect 570092 331740 570156 331804
rect 565860 331332 565924 331396
rect 286916 331196 286980 331260
rect 566596 331196 566660 331260
rect 23244 330924 23308 330988
rect 298692 330516 298756 330580
rect 21772 330380 21836 330444
rect 298692 329700 298756 329764
rect 296116 329020 296180 329084
rect 303476 318004 303540 318068
rect 285444 316704 285508 316708
rect 285444 316648 285458 316704
rect 285458 316648 285508 316704
rect 285444 316644 285508 316648
rect 290044 316644 290108 316708
rect 21956 315888 22020 315892
rect 21956 315832 22006 315888
rect 22006 315832 22020 315888
rect 21956 315828 22020 315832
rect 566412 315888 566476 315892
rect 566412 315832 566426 315888
rect 566426 315832 566476 315888
rect 566412 315828 566476 315832
rect 300164 315420 300228 315484
rect 20484 315284 20548 315348
rect 290044 315284 290108 315348
rect 21220 314740 21284 314804
rect 21956 314740 22020 314804
rect 568620 314604 568684 314668
rect 566044 313924 566108 313988
rect 299244 307668 299308 307732
rect 285444 305628 285508 305692
rect 20484 205804 20548 205868
rect 299244 205940 299308 206004
rect 21772 205668 21836 205732
rect 301636 205668 301700 205732
rect 303476 205592 303540 205596
rect 303476 205536 303526 205592
rect 303526 205536 303540 205592
rect 303476 205532 303540 205536
rect 301452 204852 301516 204916
rect 19564 204172 19628 204236
rect 21220 204172 21284 204236
rect 286732 203628 286796 203692
rect 301636 203492 301700 203556
rect 22876 202736 22940 202740
rect 22876 202680 22926 202736
rect 22926 202680 22940 202736
rect 22876 202676 22940 202680
rect 23244 202132 23308 202196
rect 570276 201376 570340 201380
rect 570276 201320 570326 201376
rect 570326 201320 570340 201376
rect 570276 201316 570340 201320
rect 298692 201180 298756 201244
rect 298876 200636 298940 200700
rect 17724 199140 17788 199204
rect 285260 188260 285324 188324
rect 303476 188260 303540 188324
rect 569172 188260 569236 188324
rect 302004 187580 302068 187644
rect 568620 187580 568684 187644
rect 23060 186356 23124 186420
rect 286180 186084 286244 186148
rect 21772 185948 21836 186012
rect 298692 185812 298756 185876
rect 285260 177924 285324 177988
rect 565308 79324 565372 79388
rect 21772 77828 21836 77892
rect 303476 77888 303540 77892
rect 303476 77832 303526 77888
rect 303526 77832 303540 77888
rect 303476 77828 303540 77832
rect 302004 77692 302068 77756
rect 568620 77828 568684 77892
rect 297956 76876 298020 76940
rect 295012 76740 295076 76804
rect 302740 76740 302804 76804
rect 301636 76604 301700 76668
rect 567332 76604 567396 76668
rect 287652 76468 287716 76532
rect 569908 76468 569972 76532
rect 575244 76468 575308 76532
rect 292436 76332 292500 76396
rect 571380 76120 571444 76124
rect 571380 76064 571430 76120
rect 571430 76064 571444 76120
rect 571380 76060 571444 76064
rect 22876 75924 22940 75988
rect 23060 75788 23124 75852
rect 21956 75652 22020 75716
rect 19564 75516 19628 75580
rect 298876 73884 298940 73948
rect 296116 73748 296180 73812
rect 17724 71708 17788 71772
rect 570092 71708 570156 71772
rect 566044 69668 566108 69732
rect 565308 68852 565372 68916
rect 298692 68172 298756 68236
rect 565860 62732 565924 62796
rect 292804 59876 292868 59940
rect 295932 59876 295996 59940
rect 291148 57428 291212 57492
rect 290044 57292 290108 57356
rect 297772 57292 297836 57356
rect 286916 57156 286980 57220
rect 288204 54844 288268 54908
rect 292620 54708 292684 54772
rect 289860 54572 289924 54636
rect 299980 54572 300044 54636
rect 289124 54436 289188 54500
rect 300164 54436 300228 54500
rect 566964 54436 567028 54500
rect 286180 53892 286244 53956
rect 288940 53076 289004 53140
rect 19196 34580 19260 34644
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 700000 51914 700398
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 700000 87914 700398
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 700000 123914 700398
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 700000 159914 700398
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 700000 195914 700398
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 700000 231914 700398
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 700000 267914 700398
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 288939 700364 289005 700365
rect 288939 700300 288940 700364
rect 289004 700300 289005 700364
rect 288939 700299 289005 700300
rect 19195 699820 19261 699821
rect 19195 699756 19196 699820
rect 19260 699756 19261 699820
rect 19195 699755 19261 699756
rect 287651 699820 287717 699821
rect 287651 699756 287652 699820
rect 287716 699756 287717 699820
rect 287651 699755 287717 699756
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 17723 582996 17789 582997
rect 17723 582932 17724 582996
rect 17788 582932 17789 582996
rect 17723 582931 17789 582932
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 17726 460189 17786 582931
rect 17723 460188 17789 460189
rect 17723 460124 17724 460188
rect 17788 460124 17789 460188
rect 17723 460123 17789 460124
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 17723 199204 17789 199205
rect 17723 199140 17724 199204
rect 17788 199140 17789 199204
rect 17723 199139 17789 199140
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 17726 71773 17786 199139
rect 17723 71772 17789 71773
rect 17723 71708 17724 71772
rect 17788 71708 17789 71772
rect 17723 71707 17789 71708
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 19198 34645 19258 699755
rect 33868 691954 34868 691986
rect 33868 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 34868 691954
rect 33868 691634 34868 691718
rect 33868 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 34868 691634
rect 33868 691366 34868 691398
rect 53868 691954 54868 691986
rect 53868 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 54868 691954
rect 53868 691634 54868 691718
rect 53868 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 54868 691634
rect 53868 691366 54868 691398
rect 73868 691954 74868 691986
rect 73868 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 74868 691954
rect 73868 691634 74868 691718
rect 73868 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 74868 691634
rect 73868 691366 74868 691398
rect 93868 691954 94868 691986
rect 93868 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 94868 691954
rect 93868 691634 94868 691718
rect 93868 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 94868 691634
rect 93868 691366 94868 691398
rect 113868 691954 114868 691986
rect 113868 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 114868 691954
rect 113868 691634 114868 691718
rect 113868 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 114868 691634
rect 113868 691366 114868 691398
rect 133868 691954 134868 691986
rect 133868 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 134868 691954
rect 133868 691634 134868 691718
rect 133868 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 134868 691634
rect 133868 691366 134868 691398
rect 153868 691954 154868 691986
rect 153868 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 154868 691954
rect 153868 691634 154868 691718
rect 153868 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 154868 691634
rect 153868 691366 154868 691398
rect 173868 691954 174868 691986
rect 173868 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 174868 691954
rect 173868 691634 174868 691718
rect 173868 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 174868 691634
rect 173868 691366 174868 691398
rect 193868 691954 194868 691986
rect 193868 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 194868 691954
rect 193868 691634 194868 691718
rect 193868 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 194868 691634
rect 193868 691366 194868 691398
rect 213868 691954 214868 691986
rect 213868 691718 213930 691954
rect 214166 691718 214250 691954
rect 214486 691718 214570 691954
rect 214806 691718 214868 691954
rect 213868 691634 214868 691718
rect 213868 691398 213930 691634
rect 214166 691398 214250 691634
rect 214486 691398 214570 691634
rect 214806 691398 214868 691634
rect 213868 691366 214868 691398
rect 233868 691954 234868 691986
rect 233868 691718 233930 691954
rect 234166 691718 234250 691954
rect 234486 691718 234570 691954
rect 234806 691718 234868 691954
rect 233868 691634 234868 691718
rect 233868 691398 233930 691634
rect 234166 691398 234250 691634
rect 234486 691398 234570 691634
rect 234806 691398 234868 691634
rect 233868 691366 234868 691398
rect 253868 691954 254868 691986
rect 253868 691718 253930 691954
rect 254166 691718 254250 691954
rect 254486 691718 254570 691954
rect 254806 691718 254868 691954
rect 253868 691634 254868 691718
rect 253868 691398 253930 691634
rect 254166 691398 254250 691634
rect 254486 691398 254570 691634
rect 254806 691398 254868 691634
rect 253868 691366 254868 691398
rect 273868 691954 274868 691986
rect 273868 691718 273930 691954
rect 274166 691718 274250 691954
rect 274486 691718 274570 691954
rect 274806 691718 274868 691954
rect 273868 691634 274868 691718
rect 273868 691398 273930 691634
rect 274166 691398 274250 691634
rect 274486 691398 274570 691634
rect 274806 691398 274868 691634
rect 273868 691366 274868 691398
rect 23868 687454 24868 687486
rect 23868 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 24868 687454
rect 23868 687134 24868 687218
rect 23868 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 24868 687134
rect 23868 686866 24868 686898
rect 43868 687454 44868 687486
rect 43868 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 44868 687454
rect 43868 687134 44868 687218
rect 43868 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 44868 687134
rect 43868 686866 44868 686898
rect 63868 687454 64868 687486
rect 63868 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 64868 687454
rect 63868 687134 64868 687218
rect 63868 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 64868 687134
rect 63868 686866 64868 686898
rect 83868 687454 84868 687486
rect 83868 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 84868 687454
rect 83868 687134 84868 687218
rect 83868 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 84868 687134
rect 83868 686866 84868 686898
rect 103868 687454 104868 687486
rect 103868 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 104868 687454
rect 103868 687134 104868 687218
rect 103868 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 104868 687134
rect 103868 686866 104868 686898
rect 123868 687454 124868 687486
rect 123868 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 124868 687454
rect 123868 687134 124868 687218
rect 123868 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 124868 687134
rect 123868 686866 124868 686898
rect 143868 687454 144868 687486
rect 143868 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 144868 687454
rect 143868 687134 144868 687218
rect 143868 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 144868 687134
rect 143868 686866 144868 686898
rect 163868 687454 164868 687486
rect 163868 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 164868 687454
rect 163868 687134 164868 687218
rect 163868 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 164868 687134
rect 163868 686866 164868 686898
rect 183868 687454 184868 687486
rect 183868 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 184868 687454
rect 183868 687134 184868 687218
rect 183868 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 184868 687134
rect 183868 686866 184868 686898
rect 203868 687454 204868 687486
rect 203868 687218 203930 687454
rect 204166 687218 204250 687454
rect 204486 687218 204570 687454
rect 204806 687218 204868 687454
rect 203868 687134 204868 687218
rect 203868 686898 203930 687134
rect 204166 686898 204250 687134
rect 204486 686898 204570 687134
rect 204806 686898 204868 687134
rect 203868 686866 204868 686898
rect 223868 687454 224868 687486
rect 223868 687218 223930 687454
rect 224166 687218 224250 687454
rect 224486 687218 224570 687454
rect 224806 687218 224868 687454
rect 223868 687134 224868 687218
rect 223868 686898 223930 687134
rect 224166 686898 224250 687134
rect 224486 686898 224570 687134
rect 224806 686898 224868 687134
rect 223868 686866 224868 686898
rect 243868 687454 244868 687486
rect 243868 687218 243930 687454
rect 244166 687218 244250 687454
rect 244486 687218 244570 687454
rect 244806 687218 244868 687454
rect 243868 687134 244868 687218
rect 243868 686898 243930 687134
rect 244166 686898 244250 687134
rect 244486 686898 244570 687134
rect 244806 686898 244868 687134
rect 243868 686866 244868 686898
rect 263868 687454 264868 687486
rect 263868 687218 263930 687454
rect 264166 687218 264250 687454
rect 264486 687218 264570 687454
rect 264806 687218 264868 687454
rect 263868 687134 264868 687218
rect 263868 686898 263930 687134
rect 264166 686898 264250 687134
rect 264486 686898 264570 687134
rect 264806 686898 264868 687134
rect 263868 686866 264868 686898
rect 283868 687454 284868 687486
rect 283868 687218 283930 687454
rect 284166 687218 284250 687454
rect 284486 687218 284570 687454
rect 284806 687218 284868 687454
rect 283868 687134 284868 687218
rect 283868 686898 283930 687134
rect 284166 686898 284250 687134
rect 284486 686898 284570 687134
rect 284806 686898 284868 687134
rect 283868 686866 284868 686898
rect 33868 655954 34868 655986
rect 33868 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 34868 655954
rect 33868 655634 34868 655718
rect 33868 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 34868 655634
rect 33868 655366 34868 655398
rect 53868 655954 54868 655986
rect 53868 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 54868 655954
rect 53868 655634 54868 655718
rect 53868 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 54868 655634
rect 53868 655366 54868 655398
rect 73868 655954 74868 655986
rect 73868 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 74868 655954
rect 73868 655634 74868 655718
rect 73868 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 74868 655634
rect 73868 655366 74868 655398
rect 93868 655954 94868 655986
rect 93868 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 94868 655954
rect 93868 655634 94868 655718
rect 93868 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 94868 655634
rect 93868 655366 94868 655398
rect 113868 655954 114868 655986
rect 113868 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 114868 655954
rect 113868 655634 114868 655718
rect 113868 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 114868 655634
rect 113868 655366 114868 655398
rect 133868 655954 134868 655986
rect 133868 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 134868 655954
rect 133868 655634 134868 655718
rect 133868 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 134868 655634
rect 133868 655366 134868 655398
rect 153868 655954 154868 655986
rect 153868 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 154868 655954
rect 153868 655634 154868 655718
rect 153868 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 154868 655634
rect 153868 655366 154868 655398
rect 173868 655954 174868 655986
rect 173868 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 174868 655954
rect 173868 655634 174868 655718
rect 173868 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 174868 655634
rect 173868 655366 174868 655398
rect 193868 655954 194868 655986
rect 193868 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 194868 655954
rect 193868 655634 194868 655718
rect 193868 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 194868 655634
rect 193868 655366 194868 655398
rect 213868 655954 214868 655986
rect 213868 655718 213930 655954
rect 214166 655718 214250 655954
rect 214486 655718 214570 655954
rect 214806 655718 214868 655954
rect 213868 655634 214868 655718
rect 213868 655398 213930 655634
rect 214166 655398 214250 655634
rect 214486 655398 214570 655634
rect 214806 655398 214868 655634
rect 213868 655366 214868 655398
rect 233868 655954 234868 655986
rect 233868 655718 233930 655954
rect 234166 655718 234250 655954
rect 234486 655718 234570 655954
rect 234806 655718 234868 655954
rect 233868 655634 234868 655718
rect 233868 655398 233930 655634
rect 234166 655398 234250 655634
rect 234486 655398 234570 655634
rect 234806 655398 234868 655634
rect 233868 655366 234868 655398
rect 253868 655954 254868 655986
rect 253868 655718 253930 655954
rect 254166 655718 254250 655954
rect 254486 655718 254570 655954
rect 254806 655718 254868 655954
rect 253868 655634 254868 655718
rect 253868 655398 253930 655634
rect 254166 655398 254250 655634
rect 254486 655398 254570 655634
rect 254806 655398 254868 655634
rect 253868 655366 254868 655398
rect 273868 655954 274868 655986
rect 273868 655718 273930 655954
rect 274166 655718 274250 655954
rect 274486 655718 274570 655954
rect 274806 655718 274868 655954
rect 273868 655634 274868 655718
rect 273868 655398 273930 655634
rect 274166 655398 274250 655634
rect 274486 655398 274570 655634
rect 274806 655398 274868 655634
rect 273868 655366 274868 655398
rect 23868 651454 24868 651486
rect 23868 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 24868 651454
rect 23868 651134 24868 651218
rect 23868 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 24868 651134
rect 23868 650866 24868 650898
rect 43868 651454 44868 651486
rect 43868 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 44868 651454
rect 43868 651134 44868 651218
rect 43868 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 44868 651134
rect 43868 650866 44868 650898
rect 63868 651454 64868 651486
rect 63868 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 64868 651454
rect 63868 651134 64868 651218
rect 63868 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 64868 651134
rect 63868 650866 64868 650898
rect 83868 651454 84868 651486
rect 83868 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 84868 651454
rect 83868 651134 84868 651218
rect 83868 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 84868 651134
rect 83868 650866 84868 650898
rect 103868 651454 104868 651486
rect 103868 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 104868 651454
rect 103868 651134 104868 651218
rect 103868 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 104868 651134
rect 103868 650866 104868 650898
rect 123868 651454 124868 651486
rect 123868 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 124868 651454
rect 123868 651134 124868 651218
rect 123868 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 124868 651134
rect 123868 650866 124868 650898
rect 143868 651454 144868 651486
rect 143868 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 144868 651454
rect 143868 651134 144868 651218
rect 143868 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 144868 651134
rect 143868 650866 144868 650898
rect 163868 651454 164868 651486
rect 163868 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 164868 651454
rect 163868 651134 164868 651218
rect 163868 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 164868 651134
rect 163868 650866 164868 650898
rect 183868 651454 184868 651486
rect 183868 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 184868 651454
rect 183868 651134 184868 651218
rect 183868 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 184868 651134
rect 183868 650866 184868 650898
rect 203868 651454 204868 651486
rect 203868 651218 203930 651454
rect 204166 651218 204250 651454
rect 204486 651218 204570 651454
rect 204806 651218 204868 651454
rect 203868 651134 204868 651218
rect 203868 650898 203930 651134
rect 204166 650898 204250 651134
rect 204486 650898 204570 651134
rect 204806 650898 204868 651134
rect 203868 650866 204868 650898
rect 223868 651454 224868 651486
rect 223868 651218 223930 651454
rect 224166 651218 224250 651454
rect 224486 651218 224570 651454
rect 224806 651218 224868 651454
rect 223868 651134 224868 651218
rect 223868 650898 223930 651134
rect 224166 650898 224250 651134
rect 224486 650898 224570 651134
rect 224806 650898 224868 651134
rect 223868 650866 224868 650898
rect 243868 651454 244868 651486
rect 243868 651218 243930 651454
rect 244166 651218 244250 651454
rect 244486 651218 244570 651454
rect 244806 651218 244868 651454
rect 243868 651134 244868 651218
rect 243868 650898 243930 651134
rect 244166 650898 244250 651134
rect 244486 650898 244570 651134
rect 244806 650898 244868 651134
rect 243868 650866 244868 650898
rect 263868 651454 264868 651486
rect 263868 651218 263930 651454
rect 264166 651218 264250 651454
rect 264486 651218 264570 651454
rect 264806 651218 264868 651454
rect 263868 651134 264868 651218
rect 263868 650898 263930 651134
rect 264166 650898 264250 651134
rect 264486 650898 264570 651134
rect 264806 650898 264868 651134
rect 263868 650866 264868 650898
rect 283868 651454 284868 651486
rect 283868 651218 283930 651454
rect 284166 651218 284250 651454
rect 284486 651218 284570 651454
rect 284806 651218 284868 651454
rect 283868 651134 284868 651218
rect 283868 650898 283930 651134
rect 284166 650898 284250 651134
rect 284486 650898 284570 651134
rect 284806 650898 284868 651134
rect 283868 650866 284868 650898
rect 33868 619954 34868 619986
rect 33868 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 34868 619954
rect 33868 619634 34868 619718
rect 33868 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 34868 619634
rect 33868 619366 34868 619398
rect 53868 619954 54868 619986
rect 53868 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 54868 619954
rect 53868 619634 54868 619718
rect 53868 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 54868 619634
rect 53868 619366 54868 619398
rect 73868 619954 74868 619986
rect 73868 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 74868 619954
rect 73868 619634 74868 619718
rect 73868 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 74868 619634
rect 73868 619366 74868 619398
rect 93868 619954 94868 619986
rect 93868 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 94868 619954
rect 93868 619634 94868 619718
rect 93868 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 94868 619634
rect 93868 619366 94868 619398
rect 113868 619954 114868 619986
rect 113868 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 114868 619954
rect 113868 619634 114868 619718
rect 113868 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 114868 619634
rect 113868 619366 114868 619398
rect 133868 619954 134868 619986
rect 133868 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 134868 619954
rect 133868 619634 134868 619718
rect 133868 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 134868 619634
rect 133868 619366 134868 619398
rect 153868 619954 154868 619986
rect 153868 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 154868 619954
rect 153868 619634 154868 619718
rect 153868 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 154868 619634
rect 153868 619366 154868 619398
rect 173868 619954 174868 619986
rect 173868 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 174868 619954
rect 173868 619634 174868 619718
rect 173868 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 174868 619634
rect 173868 619366 174868 619398
rect 193868 619954 194868 619986
rect 193868 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 194868 619954
rect 193868 619634 194868 619718
rect 193868 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 194868 619634
rect 193868 619366 194868 619398
rect 213868 619954 214868 619986
rect 213868 619718 213930 619954
rect 214166 619718 214250 619954
rect 214486 619718 214570 619954
rect 214806 619718 214868 619954
rect 213868 619634 214868 619718
rect 213868 619398 213930 619634
rect 214166 619398 214250 619634
rect 214486 619398 214570 619634
rect 214806 619398 214868 619634
rect 213868 619366 214868 619398
rect 233868 619954 234868 619986
rect 233868 619718 233930 619954
rect 234166 619718 234250 619954
rect 234486 619718 234570 619954
rect 234806 619718 234868 619954
rect 233868 619634 234868 619718
rect 233868 619398 233930 619634
rect 234166 619398 234250 619634
rect 234486 619398 234570 619634
rect 234806 619398 234868 619634
rect 233868 619366 234868 619398
rect 253868 619954 254868 619986
rect 253868 619718 253930 619954
rect 254166 619718 254250 619954
rect 254486 619718 254570 619954
rect 254806 619718 254868 619954
rect 253868 619634 254868 619718
rect 253868 619398 253930 619634
rect 254166 619398 254250 619634
rect 254486 619398 254570 619634
rect 254806 619398 254868 619634
rect 253868 619366 254868 619398
rect 273868 619954 274868 619986
rect 273868 619718 273930 619954
rect 274166 619718 274250 619954
rect 274486 619718 274570 619954
rect 274806 619718 274868 619954
rect 273868 619634 274868 619718
rect 273868 619398 273930 619634
rect 274166 619398 274250 619634
rect 274486 619398 274570 619634
rect 274806 619398 274868 619634
rect 273868 619366 274868 619398
rect 23868 615454 24868 615486
rect 23868 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 24868 615454
rect 23868 615134 24868 615218
rect 23868 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 24868 615134
rect 23868 614866 24868 614898
rect 43868 615454 44868 615486
rect 43868 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 44868 615454
rect 43868 615134 44868 615218
rect 43868 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 44868 615134
rect 43868 614866 44868 614898
rect 63868 615454 64868 615486
rect 63868 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 64868 615454
rect 63868 615134 64868 615218
rect 63868 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 64868 615134
rect 63868 614866 64868 614898
rect 83868 615454 84868 615486
rect 83868 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 84868 615454
rect 83868 615134 84868 615218
rect 83868 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 84868 615134
rect 83868 614866 84868 614898
rect 103868 615454 104868 615486
rect 103868 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 104868 615454
rect 103868 615134 104868 615218
rect 103868 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 104868 615134
rect 103868 614866 104868 614898
rect 123868 615454 124868 615486
rect 123868 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 124868 615454
rect 123868 615134 124868 615218
rect 123868 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 124868 615134
rect 123868 614866 124868 614898
rect 143868 615454 144868 615486
rect 143868 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 144868 615454
rect 143868 615134 144868 615218
rect 143868 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 144868 615134
rect 143868 614866 144868 614898
rect 163868 615454 164868 615486
rect 163868 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 164868 615454
rect 163868 615134 164868 615218
rect 163868 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 164868 615134
rect 163868 614866 164868 614898
rect 183868 615454 184868 615486
rect 183868 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 184868 615454
rect 183868 615134 184868 615218
rect 183868 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 184868 615134
rect 183868 614866 184868 614898
rect 203868 615454 204868 615486
rect 203868 615218 203930 615454
rect 204166 615218 204250 615454
rect 204486 615218 204570 615454
rect 204806 615218 204868 615454
rect 203868 615134 204868 615218
rect 203868 614898 203930 615134
rect 204166 614898 204250 615134
rect 204486 614898 204570 615134
rect 204806 614898 204868 615134
rect 203868 614866 204868 614898
rect 223868 615454 224868 615486
rect 223868 615218 223930 615454
rect 224166 615218 224250 615454
rect 224486 615218 224570 615454
rect 224806 615218 224868 615454
rect 223868 615134 224868 615218
rect 223868 614898 223930 615134
rect 224166 614898 224250 615134
rect 224486 614898 224570 615134
rect 224806 614898 224868 615134
rect 223868 614866 224868 614898
rect 243868 615454 244868 615486
rect 243868 615218 243930 615454
rect 244166 615218 244250 615454
rect 244486 615218 244570 615454
rect 244806 615218 244868 615454
rect 243868 615134 244868 615218
rect 243868 614898 243930 615134
rect 244166 614898 244250 615134
rect 244486 614898 244570 615134
rect 244806 614898 244868 615134
rect 243868 614866 244868 614898
rect 263868 615454 264868 615486
rect 263868 615218 263930 615454
rect 264166 615218 264250 615454
rect 264486 615218 264570 615454
rect 264806 615218 264868 615454
rect 263868 615134 264868 615218
rect 263868 614898 263930 615134
rect 264166 614898 264250 615134
rect 264486 614898 264570 615134
rect 264806 614898 264868 615134
rect 263868 614866 264868 614898
rect 283868 615454 284868 615486
rect 283868 615218 283930 615454
rect 284166 615218 284250 615454
rect 284486 615218 284570 615454
rect 284806 615218 284868 615454
rect 283868 615134 284868 615218
rect 283868 614898 283930 615134
rect 284166 614898 284250 615134
rect 284486 614898 284570 615134
rect 284806 614898 284868 615134
rect 283868 614866 284868 614898
rect 23243 585716 23309 585717
rect 23243 585652 23244 585716
rect 23308 585652 23309 585716
rect 23243 585651 23309 585652
rect 21955 570620 22021 570621
rect 21955 570556 21956 570620
rect 22020 570556 22021 570620
rect 21955 570555 22021 570556
rect 21958 460325 22018 570555
rect 21955 460324 22021 460325
rect 21955 460260 21956 460324
rect 22020 460260 22021 460324
rect 21955 460259 22021 460260
rect 23246 458149 23306 585651
rect 286179 585172 286245 585173
rect 286179 585108 286180 585172
rect 286244 585108 286245 585172
rect 286179 585107 286245 585108
rect 285627 582996 285693 582997
rect 285627 582932 285628 582996
rect 285692 582932 285693 582996
rect 285627 582931 285693 582932
rect 33868 547954 34868 547986
rect 33868 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 34868 547954
rect 33868 547634 34868 547718
rect 33868 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 34868 547634
rect 33868 547366 34868 547398
rect 53868 547954 54868 547986
rect 53868 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 54868 547954
rect 53868 547634 54868 547718
rect 53868 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 54868 547634
rect 53868 547366 54868 547398
rect 73868 547954 74868 547986
rect 73868 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 74868 547954
rect 73868 547634 74868 547718
rect 73868 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 74868 547634
rect 73868 547366 74868 547398
rect 93868 547954 94868 547986
rect 93868 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 94868 547954
rect 93868 547634 94868 547718
rect 93868 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 94868 547634
rect 93868 547366 94868 547398
rect 113868 547954 114868 547986
rect 113868 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 114868 547954
rect 113868 547634 114868 547718
rect 113868 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 114868 547634
rect 113868 547366 114868 547398
rect 133868 547954 134868 547986
rect 133868 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 134868 547954
rect 133868 547634 134868 547718
rect 133868 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 134868 547634
rect 133868 547366 134868 547398
rect 153868 547954 154868 547986
rect 153868 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 154868 547954
rect 153868 547634 154868 547718
rect 153868 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 154868 547634
rect 153868 547366 154868 547398
rect 173868 547954 174868 547986
rect 173868 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 174868 547954
rect 173868 547634 174868 547718
rect 173868 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 174868 547634
rect 173868 547366 174868 547398
rect 193868 547954 194868 547986
rect 193868 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 194868 547954
rect 193868 547634 194868 547718
rect 193868 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 194868 547634
rect 193868 547366 194868 547398
rect 213868 547954 214868 547986
rect 213868 547718 213930 547954
rect 214166 547718 214250 547954
rect 214486 547718 214570 547954
rect 214806 547718 214868 547954
rect 213868 547634 214868 547718
rect 213868 547398 213930 547634
rect 214166 547398 214250 547634
rect 214486 547398 214570 547634
rect 214806 547398 214868 547634
rect 213868 547366 214868 547398
rect 233868 547954 234868 547986
rect 233868 547718 233930 547954
rect 234166 547718 234250 547954
rect 234486 547718 234570 547954
rect 234806 547718 234868 547954
rect 233868 547634 234868 547718
rect 233868 547398 233930 547634
rect 234166 547398 234250 547634
rect 234486 547398 234570 547634
rect 234806 547398 234868 547634
rect 233868 547366 234868 547398
rect 253868 547954 254868 547986
rect 253868 547718 253930 547954
rect 254166 547718 254250 547954
rect 254486 547718 254570 547954
rect 254806 547718 254868 547954
rect 253868 547634 254868 547718
rect 253868 547398 253930 547634
rect 254166 547398 254250 547634
rect 254486 547398 254570 547634
rect 254806 547398 254868 547634
rect 253868 547366 254868 547398
rect 273868 547954 274868 547986
rect 273868 547718 273930 547954
rect 274166 547718 274250 547954
rect 274486 547718 274570 547954
rect 274806 547718 274868 547954
rect 273868 547634 274868 547718
rect 273868 547398 273930 547634
rect 274166 547398 274250 547634
rect 274486 547398 274570 547634
rect 274806 547398 274868 547634
rect 273868 547366 274868 547398
rect 23868 543454 24868 543486
rect 23868 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 24868 543454
rect 23868 543134 24868 543218
rect 23868 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 24868 543134
rect 23868 542866 24868 542898
rect 43868 543454 44868 543486
rect 43868 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 44868 543454
rect 43868 543134 44868 543218
rect 43868 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 44868 543134
rect 43868 542866 44868 542898
rect 63868 543454 64868 543486
rect 63868 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 64868 543454
rect 63868 543134 64868 543218
rect 63868 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 64868 543134
rect 63868 542866 64868 542898
rect 83868 543454 84868 543486
rect 83868 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 84868 543454
rect 83868 543134 84868 543218
rect 83868 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 84868 543134
rect 83868 542866 84868 542898
rect 103868 543454 104868 543486
rect 103868 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 104868 543454
rect 103868 543134 104868 543218
rect 103868 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 104868 543134
rect 103868 542866 104868 542898
rect 123868 543454 124868 543486
rect 123868 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 124868 543454
rect 123868 543134 124868 543218
rect 123868 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 124868 543134
rect 123868 542866 124868 542898
rect 143868 543454 144868 543486
rect 143868 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 144868 543454
rect 143868 543134 144868 543218
rect 143868 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 144868 543134
rect 143868 542866 144868 542898
rect 163868 543454 164868 543486
rect 163868 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 164868 543454
rect 163868 543134 164868 543218
rect 163868 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 164868 543134
rect 163868 542866 164868 542898
rect 183868 543454 184868 543486
rect 183868 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 184868 543454
rect 183868 543134 184868 543218
rect 183868 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 184868 543134
rect 183868 542866 184868 542898
rect 203868 543454 204868 543486
rect 203868 543218 203930 543454
rect 204166 543218 204250 543454
rect 204486 543218 204570 543454
rect 204806 543218 204868 543454
rect 203868 543134 204868 543218
rect 203868 542898 203930 543134
rect 204166 542898 204250 543134
rect 204486 542898 204570 543134
rect 204806 542898 204868 543134
rect 203868 542866 204868 542898
rect 223868 543454 224868 543486
rect 223868 543218 223930 543454
rect 224166 543218 224250 543454
rect 224486 543218 224570 543454
rect 224806 543218 224868 543454
rect 223868 543134 224868 543218
rect 223868 542898 223930 543134
rect 224166 542898 224250 543134
rect 224486 542898 224570 543134
rect 224806 542898 224868 543134
rect 223868 542866 224868 542898
rect 243868 543454 244868 543486
rect 243868 543218 243930 543454
rect 244166 543218 244250 543454
rect 244486 543218 244570 543454
rect 244806 543218 244868 543454
rect 243868 543134 244868 543218
rect 243868 542898 243930 543134
rect 244166 542898 244250 543134
rect 244486 542898 244570 543134
rect 244806 542898 244868 543134
rect 243868 542866 244868 542898
rect 263868 543454 264868 543486
rect 263868 543218 263930 543454
rect 264166 543218 264250 543454
rect 264486 543218 264570 543454
rect 264806 543218 264868 543454
rect 263868 543134 264868 543218
rect 263868 542898 263930 543134
rect 264166 542898 264250 543134
rect 264486 542898 264570 543134
rect 264806 542898 264868 543134
rect 263868 542866 264868 542898
rect 283868 543454 284868 543486
rect 283868 543218 283930 543454
rect 284166 543218 284250 543454
rect 284486 543218 284570 543454
rect 284806 543218 284868 543454
rect 283868 543134 284868 543218
rect 283868 542898 283930 543134
rect 284166 542898 284250 543134
rect 284486 542898 284570 543134
rect 284806 542898 284868 543134
rect 283868 542866 284868 542898
rect 33868 511954 34868 511986
rect 33868 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 34868 511954
rect 33868 511634 34868 511718
rect 33868 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 34868 511634
rect 33868 511366 34868 511398
rect 53868 511954 54868 511986
rect 53868 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 54868 511954
rect 53868 511634 54868 511718
rect 53868 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 54868 511634
rect 53868 511366 54868 511398
rect 73868 511954 74868 511986
rect 73868 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 74868 511954
rect 73868 511634 74868 511718
rect 73868 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 74868 511634
rect 73868 511366 74868 511398
rect 93868 511954 94868 511986
rect 93868 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 94868 511954
rect 93868 511634 94868 511718
rect 93868 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 94868 511634
rect 93868 511366 94868 511398
rect 113868 511954 114868 511986
rect 113868 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 114868 511954
rect 113868 511634 114868 511718
rect 113868 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 114868 511634
rect 113868 511366 114868 511398
rect 133868 511954 134868 511986
rect 133868 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 134868 511954
rect 133868 511634 134868 511718
rect 133868 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 134868 511634
rect 133868 511366 134868 511398
rect 153868 511954 154868 511986
rect 153868 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 154868 511954
rect 153868 511634 154868 511718
rect 153868 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 154868 511634
rect 153868 511366 154868 511398
rect 173868 511954 174868 511986
rect 173868 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 174868 511954
rect 173868 511634 174868 511718
rect 173868 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 174868 511634
rect 173868 511366 174868 511398
rect 193868 511954 194868 511986
rect 193868 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 194868 511954
rect 193868 511634 194868 511718
rect 193868 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 194868 511634
rect 193868 511366 194868 511398
rect 213868 511954 214868 511986
rect 213868 511718 213930 511954
rect 214166 511718 214250 511954
rect 214486 511718 214570 511954
rect 214806 511718 214868 511954
rect 213868 511634 214868 511718
rect 213868 511398 213930 511634
rect 214166 511398 214250 511634
rect 214486 511398 214570 511634
rect 214806 511398 214868 511634
rect 213868 511366 214868 511398
rect 233868 511954 234868 511986
rect 233868 511718 233930 511954
rect 234166 511718 234250 511954
rect 234486 511718 234570 511954
rect 234806 511718 234868 511954
rect 233868 511634 234868 511718
rect 233868 511398 233930 511634
rect 234166 511398 234250 511634
rect 234486 511398 234570 511634
rect 234806 511398 234868 511634
rect 233868 511366 234868 511398
rect 253868 511954 254868 511986
rect 253868 511718 253930 511954
rect 254166 511718 254250 511954
rect 254486 511718 254570 511954
rect 254806 511718 254868 511954
rect 253868 511634 254868 511718
rect 253868 511398 253930 511634
rect 254166 511398 254250 511634
rect 254486 511398 254570 511634
rect 254806 511398 254868 511634
rect 253868 511366 254868 511398
rect 273868 511954 274868 511986
rect 273868 511718 273930 511954
rect 274166 511718 274250 511954
rect 274486 511718 274570 511954
rect 274806 511718 274868 511954
rect 273868 511634 274868 511718
rect 273868 511398 273930 511634
rect 274166 511398 274250 511634
rect 274486 511398 274570 511634
rect 274806 511398 274868 511634
rect 273868 511366 274868 511398
rect 23868 507454 24868 507486
rect 23868 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 24868 507454
rect 23868 507134 24868 507218
rect 23868 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 24868 507134
rect 23868 506866 24868 506898
rect 43868 507454 44868 507486
rect 43868 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 44868 507454
rect 43868 507134 44868 507218
rect 43868 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 44868 507134
rect 43868 506866 44868 506898
rect 63868 507454 64868 507486
rect 63868 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 64868 507454
rect 63868 507134 64868 507218
rect 63868 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 64868 507134
rect 63868 506866 64868 506898
rect 83868 507454 84868 507486
rect 83868 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 84868 507454
rect 83868 507134 84868 507218
rect 83868 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 84868 507134
rect 83868 506866 84868 506898
rect 103868 507454 104868 507486
rect 103868 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 104868 507454
rect 103868 507134 104868 507218
rect 103868 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 104868 507134
rect 103868 506866 104868 506898
rect 123868 507454 124868 507486
rect 123868 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 124868 507454
rect 123868 507134 124868 507218
rect 123868 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 124868 507134
rect 123868 506866 124868 506898
rect 143868 507454 144868 507486
rect 143868 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 144868 507454
rect 143868 507134 144868 507218
rect 143868 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 144868 507134
rect 143868 506866 144868 506898
rect 163868 507454 164868 507486
rect 163868 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 164868 507454
rect 163868 507134 164868 507218
rect 163868 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 164868 507134
rect 163868 506866 164868 506898
rect 183868 507454 184868 507486
rect 183868 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 184868 507454
rect 183868 507134 184868 507218
rect 183868 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 184868 507134
rect 183868 506866 184868 506898
rect 203868 507454 204868 507486
rect 203868 507218 203930 507454
rect 204166 507218 204250 507454
rect 204486 507218 204570 507454
rect 204806 507218 204868 507454
rect 203868 507134 204868 507218
rect 203868 506898 203930 507134
rect 204166 506898 204250 507134
rect 204486 506898 204570 507134
rect 204806 506898 204868 507134
rect 203868 506866 204868 506898
rect 223868 507454 224868 507486
rect 223868 507218 223930 507454
rect 224166 507218 224250 507454
rect 224486 507218 224570 507454
rect 224806 507218 224868 507454
rect 223868 507134 224868 507218
rect 223868 506898 223930 507134
rect 224166 506898 224250 507134
rect 224486 506898 224570 507134
rect 224806 506898 224868 507134
rect 223868 506866 224868 506898
rect 243868 507454 244868 507486
rect 243868 507218 243930 507454
rect 244166 507218 244250 507454
rect 244486 507218 244570 507454
rect 244806 507218 244868 507454
rect 243868 507134 244868 507218
rect 243868 506898 243930 507134
rect 244166 506898 244250 507134
rect 244486 506898 244570 507134
rect 244806 506898 244868 507134
rect 243868 506866 244868 506898
rect 263868 507454 264868 507486
rect 263868 507218 263930 507454
rect 264166 507218 264250 507454
rect 264486 507218 264570 507454
rect 264806 507218 264868 507454
rect 263868 507134 264868 507218
rect 263868 506898 263930 507134
rect 264166 506898 264250 507134
rect 264486 506898 264570 507134
rect 264806 506898 264868 507134
rect 263868 506866 264868 506898
rect 283868 507454 284868 507486
rect 283868 507218 283930 507454
rect 284166 507218 284250 507454
rect 284486 507218 284570 507454
rect 284806 507218 284868 507454
rect 283868 507134 284868 507218
rect 283868 506898 283930 507134
rect 284166 506898 284250 507134
rect 284486 506898 284570 507134
rect 284806 506898 284868 507134
rect 283868 506866 284868 506898
rect 33868 475954 34868 475986
rect 33868 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 34868 475954
rect 33868 475634 34868 475718
rect 33868 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 34868 475634
rect 33868 475366 34868 475398
rect 53868 475954 54868 475986
rect 53868 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 54868 475954
rect 53868 475634 54868 475718
rect 53868 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 54868 475634
rect 53868 475366 54868 475398
rect 73868 475954 74868 475986
rect 73868 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 74868 475954
rect 73868 475634 74868 475718
rect 73868 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 74868 475634
rect 73868 475366 74868 475398
rect 93868 475954 94868 475986
rect 93868 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 94868 475954
rect 93868 475634 94868 475718
rect 93868 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 94868 475634
rect 93868 475366 94868 475398
rect 113868 475954 114868 475986
rect 113868 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 114868 475954
rect 113868 475634 114868 475718
rect 113868 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 114868 475634
rect 113868 475366 114868 475398
rect 133868 475954 134868 475986
rect 133868 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 134868 475954
rect 133868 475634 134868 475718
rect 133868 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 134868 475634
rect 133868 475366 134868 475398
rect 153868 475954 154868 475986
rect 153868 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 154868 475954
rect 153868 475634 154868 475718
rect 153868 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 154868 475634
rect 153868 475366 154868 475398
rect 173868 475954 174868 475986
rect 173868 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 174868 475954
rect 173868 475634 174868 475718
rect 173868 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 174868 475634
rect 173868 475366 174868 475398
rect 193868 475954 194868 475986
rect 193868 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 194868 475954
rect 193868 475634 194868 475718
rect 193868 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 194868 475634
rect 193868 475366 194868 475398
rect 213868 475954 214868 475986
rect 213868 475718 213930 475954
rect 214166 475718 214250 475954
rect 214486 475718 214570 475954
rect 214806 475718 214868 475954
rect 213868 475634 214868 475718
rect 213868 475398 213930 475634
rect 214166 475398 214250 475634
rect 214486 475398 214570 475634
rect 214806 475398 214868 475634
rect 213868 475366 214868 475398
rect 233868 475954 234868 475986
rect 233868 475718 233930 475954
rect 234166 475718 234250 475954
rect 234486 475718 234570 475954
rect 234806 475718 234868 475954
rect 233868 475634 234868 475718
rect 233868 475398 233930 475634
rect 234166 475398 234250 475634
rect 234486 475398 234570 475634
rect 234806 475398 234868 475634
rect 233868 475366 234868 475398
rect 253868 475954 254868 475986
rect 253868 475718 253930 475954
rect 254166 475718 254250 475954
rect 254486 475718 254570 475954
rect 254806 475718 254868 475954
rect 253868 475634 254868 475718
rect 253868 475398 253930 475634
rect 254166 475398 254250 475634
rect 254486 475398 254570 475634
rect 254806 475398 254868 475634
rect 253868 475366 254868 475398
rect 273868 475954 274868 475986
rect 273868 475718 273930 475954
rect 274166 475718 274250 475954
rect 274486 475718 274570 475954
rect 274806 475718 274868 475954
rect 273868 475634 274868 475718
rect 273868 475398 273930 475634
rect 274166 475398 274250 475634
rect 274486 475398 274570 475634
rect 274806 475398 274868 475634
rect 273868 475366 274868 475398
rect 23868 471454 24868 471486
rect 23868 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 24868 471454
rect 23868 471134 24868 471218
rect 23868 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 24868 471134
rect 23868 470866 24868 470898
rect 43868 471454 44868 471486
rect 43868 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 44868 471454
rect 43868 471134 44868 471218
rect 43868 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 44868 471134
rect 43868 470866 44868 470898
rect 63868 471454 64868 471486
rect 63868 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 64868 471454
rect 63868 471134 64868 471218
rect 63868 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 64868 471134
rect 63868 470866 64868 470898
rect 83868 471454 84868 471486
rect 83868 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 84868 471454
rect 83868 471134 84868 471218
rect 83868 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 84868 471134
rect 83868 470866 84868 470898
rect 103868 471454 104868 471486
rect 103868 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 104868 471454
rect 103868 471134 104868 471218
rect 103868 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 104868 471134
rect 103868 470866 104868 470898
rect 123868 471454 124868 471486
rect 123868 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 124868 471454
rect 123868 471134 124868 471218
rect 123868 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 124868 471134
rect 123868 470866 124868 470898
rect 143868 471454 144868 471486
rect 143868 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 144868 471454
rect 143868 471134 144868 471218
rect 143868 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 144868 471134
rect 143868 470866 144868 470898
rect 163868 471454 164868 471486
rect 163868 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 164868 471454
rect 163868 471134 164868 471218
rect 163868 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 164868 471134
rect 163868 470866 164868 470898
rect 183868 471454 184868 471486
rect 183868 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 184868 471454
rect 183868 471134 184868 471218
rect 183868 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 184868 471134
rect 183868 470866 184868 470898
rect 203868 471454 204868 471486
rect 203868 471218 203930 471454
rect 204166 471218 204250 471454
rect 204486 471218 204570 471454
rect 204806 471218 204868 471454
rect 203868 471134 204868 471218
rect 203868 470898 203930 471134
rect 204166 470898 204250 471134
rect 204486 470898 204570 471134
rect 204806 470898 204868 471134
rect 203868 470866 204868 470898
rect 223868 471454 224868 471486
rect 223868 471218 223930 471454
rect 224166 471218 224250 471454
rect 224486 471218 224570 471454
rect 224806 471218 224868 471454
rect 223868 471134 224868 471218
rect 223868 470898 223930 471134
rect 224166 470898 224250 471134
rect 224486 470898 224570 471134
rect 224806 470898 224868 471134
rect 223868 470866 224868 470898
rect 243868 471454 244868 471486
rect 243868 471218 243930 471454
rect 244166 471218 244250 471454
rect 244486 471218 244570 471454
rect 244806 471218 244868 471454
rect 243868 471134 244868 471218
rect 243868 470898 243930 471134
rect 244166 470898 244250 471134
rect 244486 470898 244570 471134
rect 244806 470898 244868 471134
rect 243868 470866 244868 470898
rect 263868 471454 264868 471486
rect 263868 471218 263930 471454
rect 264166 471218 264250 471454
rect 264486 471218 264570 471454
rect 264806 471218 264868 471454
rect 263868 471134 264868 471218
rect 263868 470898 263930 471134
rect 264166 470898 264250 471134
rect 264486 470898 264570 471134
rect 264806 470898 264868 471134
rect 263868 470866 264868 470898
rect 283868 471454 284868 471486
rect 283868 471218 283930 471454
rect 284166 471218 284250 471454
rect 284486 471218 284570 471454
rect 284806 471218 284868 471454
rect 283868 471134 284868 471218
rect 283868 470898 283930 471134
rect 284166 470898 284250 471134
rect 284486 470898 284570 471134
rect 284806 470898 284868 471134
rect 283868 470866 284868 470898
rect 285443 458284 285509 458285
rect 285443 458220 285444 458284
rect 285508 458220 285509 458284
rect 285443 458219 285509 458220
rect 23243 458148 23309 458149
rect 23243 458084 23244 458148
rect 23308 458084 23309 458148
rect 23243 458083 23309 458084
rect 23246 456925 23306 458083
rect 21955 456924 22021 456925
rect 21955 456860 21956 456924
rect 22020 456860 22021 456924
rect 21955 456859 22021 456860
rect 23243 456924 23309 456925
rect 23243 456860 23244 456924
rect 23308 456860 23309 456924
rect 23243 456859 23309 456860
rect 21771 330444 21837 330445
rect 21771 330380 21772 330444
rect 21836 330380 21837 330444
rect 21771 330379 21837 330380
rect 20483 315348 20549 315349
rect 20483 315284 20484 315348
rect 20548 315284 20549 315348
rect 20483 315283 20549 315284
rect 20486 205869 20546 315283
rect 21219 314804 21285 314805
rect 21219 314740 21220 314804
rect 21284 314740 21285 314804
rect 21219 314739 21285 314740
rect 20483 205868 20549 205869
rect 20483 205804 20484 205868
rect 20548 205804 20549 205868
rect 20483 205803 20549 205804
rect 21222 204237 21282 314739
rect 21774 205733 21834 330379
rect 21958 315893 22018 456859
rect 23243 444276 23309 444277
rect 23243 444212 23244 444276
rect 23308 444212 23309 444276
rect 23243 444211 23309 444212
rect 23246 330989 23306 444211
rect 33868 439954 34868 439986
rect 33868 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 34868 439954
rect 33868 439634 34868 439718
rect 33868 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 34868 439634
rect 33868 439366 34868 439398
rect 53868 439954 54868 439986
rect 53868 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 54868 439954
rect 53868 439634 54868 439718
rect 53868 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 54868 439634
rect 53868 439366 54868 439398
rect 73868 439954 74868 439986
rect 73868 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 74868 439954
rect 73868 439634 74868 439718
rect 73868 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 74868 439634
rect 73868 439366 74868 439398
rect 93868 439954 94868 439986
rect 93868 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 94868 439954
rect 93868 439634 94868 439718
rect 93868 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 94868 439634
rect 93868 439366 94868 439398
rect 113868 439954 114868 439986
rect 113868 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 114868 439954
rect 113868 439634 114868 439718
rect 113868 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 114868 439634
rect 113868 439366 114868 439398
rect 133868 439954 134868 439986
rect 133868 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 134868 439954
rect 133868 439634 134868 439718
rect 133868 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 134868 439634
rect 133868 439366 134868 439398
rect 153868 439954 154868 439986
rect 153868 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 154868 439954
rect 153868 439634 154868 439718
rect 153868 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 154868 439634
rect 153868 439366 154868 439398
rect 173868 439954 174868 439986
rect 173868 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 174868 439954
rect 173868 439634 174868 439718
rect 173868 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 174868 439634
rect 173868 439366 174868 439398
rect 193868 439954 194868 439986
rect 193868 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 194868 439954
rect 193868 439634 194868 439718
rect 193868 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 194868 439634
rect 193868 439366 194868 439398
rect 213868 439954 214868 439986
rect 213868 439718 213930 439954
rect 214166 439718 214250 439954
rect 214486 439718 214570 439954
rect 214806 439718 214868 439954
rect 213868 439634 214868 439718
rect 213868 439398 213930 439634
rect 214166 439398 214250 439634
rect 214486 439398 214570 439634
rect 214806 439398 214868 439634
rect 213868 439366 214868 439398
rect 233868 439954 234868 439986
rect 233868 439718 233930 439954
rect 234166 439718 234250 439954
rect 234486 439718 234570 439954
rect 234806 439718 234868 439954
rect 233868 439634 234868 439718
rect 233868 439398 233930 439634
rect 234166 439398 234250 439634
rect 234486 439398 234570 439634
rect 234806 439398 234868 439634
rect 233868 439366 234868 439398
rect 253868 439954 254868 439986
rect 253868 439718 253930 439954
rect 254166 439718 254250 439954
rect 254486 439718 254570 439954
rect 254806 439718 254868 439954
rect 253868 439634 254868 439718
rect 253868 439398 253930 439634
rect 254166 439398 254250 439634
rect 254486 439398 254570 439634
rect 254806 439398 254868 439634
rect 253868 439366 254868 439398
rect 273868 439954 274868 439986
rect 273868 439718 273930 439954
rect 274166 439718 274250 439954
rect 274486 439718 274570 439954
rect 274806 439718 274868 439954
rect 273868 439634 274868 439718
rect 273868 439398 273930 439634
rect 274166 439398 274250 439634
rect 274486 439398 274570 439634
rect 274806 439398 274868 439634
rect 273868 439366 274868 439398
rect 23868 435454 24868 435486
rect 23868 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 24868 435454
rect 23868 435134 24868 435218
rect 23868 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 24868 435134
rect 23868 434866 24868 434898
rect 43868 435454 44868 435486
rect 43868 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 44868 435454
rect 43868 435134 44868 435218
rect 43868 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 44868 435134
rect 43868 434866 44868 434898
rect 63868 435454 64868 435486
rect 63868 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 64868 435454
rect 63868 435134 64868 435218
rect 63868 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 64868 435134
rect 63868 434866 64868 434898
rect 83868 435454 84868 435486
rect 83868 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 84868 435454
rect 83868 435134 84868 435218
rect 83868 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 84868 435134
rect 83868 434866 84868 434898
rect 103868 435454 104868 435486
rect 103868 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 104868 435454
rect 103868 435134 104868 435218
rect 103868 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 104868 435134
rect 103868 434866 104868 434898
rect 123868 435454 124868 435486
rect 123868 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 124868 435454
rect 123868 435134 124868 435218
rect 123868 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 124868 435134
rect 123868 434866 124868 434898
rect 143868 435454 144868 435486
rect 143868 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 144868 435454
rect 143868 435134 144868 435218
rect 143868 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 144868 435134
rect 143868 434866 144868 434898
rect 163868 435454 164868 435486
rect 163868 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 164868 435454
rect 163868 435134 164868 435218
rect 163868 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 164868 435134
rect 163868 434866 164868 434898
rect 183868 435454 184868 435486
rect 183868 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 184868 435454
rect 183868 435134 184868 435218
rect 183868 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 184868 435134
rect 183868 434866 184868 434898
rect 203868 435454 204868 435486
rect 203868 435218 203930 435454
rect 204166 435218 204250 435454
rect 204486 435218 204570 435454
rect 204806 435218 204868 435454
rect 203868 435134 204868 435218
rect 203868 434898 203930 435134
rect 204166 434898 204250 435134
rect 204486 434898 204570 435134
rect 204806 434898 204868 435134
rect 203868 434866 204868 434898
rect 223868 435454 224868 435486
rect 223868 435218 223930 435454
rect 224166 435218 224250 435454
rect 224486 435218 224570 435454
rect 224806 435218 224868 435454
rect 223868 435134 224868 435218
rect 223868 434898 223930 435134
rect 224166 434898 224250 435134
rect 224486 434898 224570 435134
rect 224806 434898 224868 435134
rect 223868 434866 224868 434898
rect 243868 435454 244868 435486
rect 243868 435218 243930 435454
rect 244166 435218 244250 435454
rect 244486 435218 244570 435454
rect 244806 435218 244868 435454
rect 243868 435134 244868 435218
rect 243868 434898 243930 435134
rect 244166 434898 244250 435134
rect 244486 434898 244570 435134
rect 244806 434898 244868 435134
rect 243868 434866 244868 434898
rect 263868 435454 264868 435486
rect 263868 435218 263930 435454
rect 264166 435218 264250 435454
rect 264486 435218 264570 435454
rect 264806 435218 264868 435454
rect 263868 435134 264868 435218
rect 263868 434898 263930 435134
rect 264166 434898 264250 435134
rect 264486 434898 264570 435134
rect 264806 434898 264868 435134
rect 263868 434866 264868 434898
rect 283868 435454 284868 435486
rect 283868 435218 283930 435454
rect 284166 435218 284250 435454
rect 284486 435218 284570 435454
rect 284806 435218 284868 435454
rect 283868 435134 284868 435218
rect 283868 434898 283930 435134
rect 284166 434898 284250 435134
rect 284486 434898 284570 435134
rect 284806 434898 284868 435134
rect 283868 434866 284868 434898
rect 285446 433941 285506 458219
rect 285630 458149 285690 582931
rect 286182 461957 286242 585107
rect 286179 461956 286245 461957
rect 286179 461892 286180 461956
rect 286244 461892 286245 461956
rect 286179 461891 286245 461892
rect 286179 460732 286245 460733
rect 286179 460668 286180 460732
rect 286244 460668 286245 460732
rect 286179 460667 286245 460668
rect 285627 458148 285693 458149
rect 285627 458084 285628 458148
rect 285692 458084 285693 458148
rect 285627 458083 285693 458084
rect 285443 433940 285509 433941
rect 285443 433876 285444 433940
rect 285508 433876 285509 433940
rect 285443 433875 285509 433876
rect 33868 403954 34868 403986
rect 33868 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 34868 403954
rect 33868 403634 34868 403718
rect 33868 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 34868 403634
rect 33868 403366 34868 403398
rect 53868 403954 54868 403986
rect 53868 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 54868 403954
rect 53868 403634 54868 403718
rect 53868 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 54868 403634
rect 53868 403366 54868 403398
rect 73868 403954 74868 403986
rect 73868 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 74868 403954
rect 73868 403634 74868 403718
rect 73868 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 74868 403634
rect 73868 403366 74868 403398
rect 93868 403954 94868 403986
rect 93868 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 94868 403954
rect 93868 403634 94868 403718
rect 93868 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 94868 403634
rect 93868 403366 94868 403398
rect 113868 403954 114868 403986
rect 113868 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 114868 403954
rect 113868 403634 114868 403718
rect 113868 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 114868 403634
rect 113868 403366 114868 403398
rect 133868 403954 134868 403986
rect 133868 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 134868 403954
rect 133868 403634 134868 403718
rect 133868 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 134868 403634
rect 133868 403366 134868 403398
rect 153868 403954 154868 403986
rect 153868 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 154868 403954
rect 153868 403634 154868 403718
rect 153868 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 154868 403634
rect 153868 403366 154868 403398
rect 173868 403954 174868 403986
rect 173868 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 174868 403954
rect 173868 403634 174868 403718
rect 173868 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 174868 403634
rect 173868 403366 174868 403398
rect 193868 403954 194868 403986
rect 193868 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 194868 403954
rect 193868 403634 194868 403718
rect 193868 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 194868 403634
rect 193868 403366 194868 403398
rect 213868 403954 214868 403986
rect 213868 403718 213930 403954
rect 214166 403718 214250 403954
rect 214486 403718 214570 403954
rect 214806 403718 214868 403954
rect 213868 403634 214868 403718
rect 213868 403398 213930 403634
rect 214166 403398 214250 403634
rect 214486 403398 214570 403634
rect 214806 403398 214868 403634
rect 213868 403366 214868 403398
rect 233868 403954 234868 403986
rect 233868 403718 233930 403954
rect 234166 403718 234250 403954
rect 234486 403718 234570 403954
rect 234806 403718 234868 403954
rect 233868 403634 234868 403718
rect 233868 403398 233930 403634
rect 234166 403398 234250 403634
rect 234486 403398 234570 403634
rect 234806 403398 234868 403634
rect 233868 403366 234868 403398
rect 253868 403954 254868 403986
rect 253868 403718 253930 403954
rect 254166 403718 254250 403954
rect 254486 403718 254570 403954
rect 254806 403718 254868 403954
rect 253868 403634 254868 403718
rect 253868 403398 253930 403634
rect 254166 403398 254250 403634
rect 254486 403398 254570 403634
rect 254806 403398 254868 403634
rect 253868 403366 254868 403398
rect 273868 403954 274868 403986
rect 273868 403718 273930 403954
rect 274166 403718 274250 403954
rect 274486 403718 274570 403954
rect 274806 403718 274868 403954
rect 273868 403634 274868 403718
rect 273868 403398 273930 403634
rect 274166 403398 274250 403634
rect 274486 403398 274570 403634
rect 274806 403398 274868 403634
rect 273868 403366 274868 403398
rect 23868 399454 24868 399486
rect 23868 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 24868 399454
rect 23868 399134 24868 399218
rect 23868 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 24868 399134
rect 23868 398866 24868 398898
rect 43868 399454 44868 399486
rect 43868 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 44868 399454
rect 43868 399134 44868 399218
rect 43868 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 44868 399134
rect 43868 398866 44868 398898
rect 63868 399454 64868 399486
rect 63868 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 64868 399454
rect 63868 399134 64868 399218
rect 63868 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 64868 399134
rect 63868 398866 64868 398898
rect 83868 399454 84868 399486
rect 83868 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 84868 399454
rect 83868 399134 84868 399218
rect 83868 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 84868 399134
rect 83868 398866 84868 398898
rect 103868 399454 104868 399486
rect 103868 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 104868 399454
rect 103868 399134 104868 399218
rect 103868 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 104868 399134
rect 103868 398866 104868 398898
rect 123868 399454 124868 399486
rect 123868 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 124868 399454
rect 123868 399134 124868 399218
rect 123868 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 124868 399134
rect 123868 398866 124868 398898
rect 143868 399454 144868 399486
rect 143868 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 144868 399454
rect 143868 399134 144868 399218
rect 143868 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 144868 399134
rect 143868 398866 144868 398898
rect 163868 399454 164868 399486
rect 163868 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 164868 399454
rect 163868 399134 164868 399218
rect 163868 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 164868 399134
rect 163868 398866 164868 398898
rect 183868 399454 184868 399486
rect 183868 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 184868 399454
rect 183868 399134 184868 399218
rect 183868 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 184868 399134
rect 183868 398866 184868 398898
rect 203868 399454 204868 399486
rect 203868 399218 203930 399454
rect 204166 399218 204250 399454
rect 204486 399218 204570 399454
rect 204806 399218 204868 399454
rect 203868 399134 204868 399218
rect 203868 398898 203930 399134
rect 204166 398898 204250 399134
rect 204486 398898 204570 399134
rect 204806 398898 204868 399134
rect 203868 398866 204868 398898
rect 223868 399454 224868 399486
rect 223868 399218 223930 399454
rect 224166 399218 224250 399454
rect 224486 399218 224570 399454
rect 224806 399218 224868 399454
rect 223868 399134 224868 399218
rect 223868 398898 223930 399134
rect 224166 398898 224250 399134
rect 224486 398898 224570 399134
rect 224806 398898 224868 399134
rect 223868 398866 224868 398898
rect 243868 399454 244868 399486
rect 243868 399218 243930 399454
rect 244166 399218 244250 399454
rect 244486 399218 244570 399454
rect 244806 399218 244868 399454
rect 243868 399134 244868 399218
rect 243868 398898 243930 399134
rect 244166 398898 244250 399134
rect 244486 398898 244570 399134
rect 244806 398898 244868 399134
rect 243868 398866 244868 398898
rect 263868 399454 264868 399486
rect 263868 399218 263930 399454
rect 264166 399218 264250 399454
rect 264486 399218 264570 399454
rect 264806 399218 264868 399454
rect 263868 399134 264868 399218
rect 263868 398898 263930 399134
rect 264166 398898 264250 399134
rect 264486 398898 264570 399134
rect 264806 398898 264868 399134
rect 263868 398866 264868 398898
rect 283868 399454 284868 399486
rect 283868 399218 283930 399454
rect 284166 399218 284250 399454
rect 284486 399218 284570 399454
rect 284806 399218 284868 399454
rect 283868 399134 284868 399218
rect 283868 398898 283930 399134
rect 284166 398898 284250 399134
rect 284486 398898 284570 399134
rect 284806 398898 284868 399134
rect 283868 398866 284868 398898
rect 33868 367954 34868 367986
rect 33868 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 34868 367954
rect 33868 367634 34868 367718
rect 33868 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 34868 367634
rect 33868 367366 34868 367398
rect 53868 367954 54868 367986
rect 53868 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 54868 367954
rect 53868 367634 54868 367718
rect 53868 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 54868 367634
rect 53868 367366 54868 367398
rect 73868 367954 74868 367986
rect 73868 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 74868 367954
rect 73868 367634 74868 367718
rect 73868 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 74868 367634
rect 73868 367366 74868 367398
rect 93868 367954 94868 367986
rect 93868 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 94868 367954
rect 93868 367634 94868 367718
rect 93868 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 94868 367634
rect 93868 367366 94868 367398
rect 113868 367954 114868 367986
rect 113868 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 114868 367954
rect 113868 367634 114868 367718
rect 113868 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 114868 367634
rect 113868 367366 114868 367398
rect 133868 367954 134868 367986
rect 133868 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 134868 367954
rect 133868 367634 134868 367718
rect 133868 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 134868 367634
rect 133868 367366 134868 367398
rect 153868 367954 154868 367986
rect 153868 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 154868 367954
rect 153868 367634 154868 367718
rect 153868 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 154868 367634
rect 153868 367366 154868 367398
rect 173868 367954 174868 367986
rect 173868 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 174868 367954
rect 173868 367634 174868 367718
rect 173868 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 174868 367634
rect 173868 367366 174868 367398
rect 193868 367954 194868 367986
rect 193868 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 194868 367954
rect 193868 367634 194868 367718
rect 193868 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 194868 367634
rect 193868 367366 194868 367398
rect 213868 367954 214868 367986
rect 213868 367718 213930 367954
rect 214166 367718 214250 367954
rect 214486 367718 214570 367954
rect 214806 367718 214868 367954
rect 213868 367634 214868 367718
rect 213868 367398 213930 367634
rect 214166 367398 214250 367634
rect 214486 367398 214570 367634
rect 214806 367398 214868 367634
rect 213868 367366 214868 367398
rect 233868 367954 234868 367986
rect 233868 367718 233930 367954
rect 234166 367718 234250 367954
rect 234486 367718 234570 367954
rect 234806 367718 234868 367954
rect 233868 367634 234868 367718
rect 233868 367398 233930 367634
rect 234166 367398 234250 367634
rect 234486 367398 234570 367634
rect 234806 367398 234868 367634
rect 233868 367366 234868 367398
rect 253868 367954 254868 367986
rect 253868 367718 253930 367954
rect 254166 367718 254250 367954
rect 254486 367718 254570 367954
rect 254806 367718 254868 367954
rect 253868 367634 254868 367718
rect 253868 367398 253930 367634
rect 254166 367398 254250 367634
rect 254486 367398 254570 367634
rect 254806 367398 254868 367634
rect 253868 367366 254868 367398
rect 273868 367954 274868 367986
rect 273868 367718 273930 367954
rect 274166 367718 274250 367954
rect 274486 367718 274570 367954
rect 274806 367718 274868 367954
rect 273868 367634 274868 367718
rect 273868 367398 273930 367634
rect 274166 367398 274250 367634
rect 274486 367398 274570 367634
rect 274806 367398 274868 367634
rect 273868 367366 274868 367398
rect 23868 363454 24868 363486
rect 23868 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 24868 363454
rect 23868 363134 24868 363218
rect 23868 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 24868 363134
rect 23868 362866 24868 362898
rect 43868 363454 44868 363486
rect 43868 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 44868 363454
rect 43868 363134 44868 363218
rect 43868 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 44868 363134
rect 43868 362866 44868 362898
rect 63868 363454 64868 363486
rect 63868 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 64868 363454
rect 63868 363134 64868 363218
rect 63868 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 64868 363134
rect 63868 362866 64868 362898
rect 83868 363454 84868 363486
rect 83868 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 84868 363454
rect 83868 363134 84868 363218
rect 83868 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 84868 363134
rect 83868 362866 84868 362898
rect 103868 363454 104868 363486
rect 103868 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 104868 363454
rect 103868 363134 104868 363218
rect 103868 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 104868 363134
rect 103868 362866 104868 362898
rect 123868 363454 124868 363486
rect 123868 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 124868 363454
rect 123868 363134 124868 363218
rect 123868 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 124868 363134
rect 123868 362866 124868 362898
rect 143868 363454 144868 363486
rect 143868 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 144868 363454
rect 143868 363134 144868 363218
rect 143868 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 144868 363134
rect 143868 362866 144868 362898
rect 163868 363454 164868 363486
rect 163868 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 164868 363454
rect 163868 363134 164868 363218
rect 163868 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 164868 363134
rect 163868 362866 164868 362898
rect 183868 363454 184868 363486
rect 183868 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 184868 363454
rect 183868 363134 184868 363218
rect 183868 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 184868 363134
rect 183868 362866 184868 362898
rect 203868 363454 204868 363486
rect 203868 363218 203930 363454
rect 204166 363218 204250 363454
rect 204486 363218 204570 363454
rect 204806 363218 204868 363454
rect 203868 363134 204868 363218
rect 203868 362898 203930 363134
rect 204166 362898 204250 363134
rect 204486 362898 204570 363134
rect 204806 362898 204868 363134
rect 203868 362866 204868 362898
rect 223868 363454 224868 363486
rect 223868 363218 223930 363454
rect 224166 363218 224250 363454
rect 224486 363218 224570 363454
rect 224806 363218 224868 363454
rect 223868 363134 224868 363218
rect 223868 362898 223930 363134
rect 224166 362898 224250 363134
rect 224486 362898 224570 363134
rect 224806 362898 224868 363134
rect 223868 362866 224868 362898
rect 243868 363454 244868 363486
rect 243868 363218 243930 363454
rect 244166 363218 244250 363454
rect 244486 363218 244570 363454
rect 244806 363218 244868 363454
rect 243868 363134 244868 363218
rect 243868 362898 243930 363134
rect 244166 362898 244250 363134
rect 244486 362898 244570 363134
rect 244806 362898 244868 363134
rect 243868 362866 244868 362898
rect 263868 363454 264868 363486
rect 263868 363218 263930 363454
rect 264166 363218 264250 363454
rect 264486 363218 264570 363454
rect 264806 363218 264868 363454
rect 263868 363134 264868 363218
rect 263868 362898 263930 363134
rect 264166 362898 264250 363134
rect 264486 362898 264570 363134
rect 264806 362898 264868 363134
rect 263868 362866 264868 362898
rect 283868 363454 284868 363486
rect 283868 363218 283930 363454
rect 284166 363218 284250 363454
rect 284486 363218 284570 363454
rect 284806 363218 284868 363454
rect 283868 363134 284868 363218
rect 283868 362898 283930 363134
rect 284166 362898 284250 363134
rect 284486 362898 284570 363134
rect 284806 362898 284868 363134
rect 283868 362866 284868 362898
rect 286182 332213 286242 460667
rect 286363 456924 286429 456925
rect 286363 456860 286364 456924
rect 286428 456860 286429 456924
rect 286363 456859 286429 456860
rect 286366 334117 286426 456859
rect 286363 334116 286429 334117
rect 286363 334052 286364 334116
rect 286428 334052 286429 334116
rect 286363 334051 286429 334052
rect 286179 332212 286245 332213
rect 286179 332148 286180 332212
rect 286244 332148 286245 332212
rect 286179 332147 286245 332148
rect 23243 330988 23309 330989
rect 23243 330924 23244 330988
rect 23308 330924 23309 330988
rect 23243 330923 23309 330924
rect 21955 315892 22021 315893
rect 21955 315828 21956 315892
rect 22020 315828 22021 315892
rect 21955 315827 22021 315828
rect 21958 314805 22018 315827
rect 21955 314804 22021 314805
rect 21955 314740 21956 314804
rect 22020 314740 22021 314804
rect 21955 314739 22021 314740
rect 21771 205732 21837 205733
rect 21771 205668 21772 205732
rect 21836 205668 21837 205732
rect 21771 205667 21837 205668
rect 19563 204236 19629 204237
rect 19563 204172 19564 204236
rect 19628 204172 19629 204236
rect 19563 204171 19629 204172
rect 21219 204236 21285 204237
rect 21219 204172 21220 204236
rect 21284 204172 21285 204236
rect 21219 204171 21285 204172
rect 19566 75581 19626 204171
rect 21222 200130 21282 204171
rect 22875 202740 22941 202741
rect 22875 202676 22876 202740
rect 22940 202676 22941 202740
rect 22875 202675 22941 202676
rect 21222 200070 22018 200130
rect 21771 186012 21837 186013
rect 21771 185948 21772 186012
rect 21836 185948 21837 186012
rect 21771 185947 21837 185948
rect 21774 77893 21834 185947
rect 21771 77892 21837 77893
rect 21771 77828 21772 77892
rect 21836 77828 21837 77892
rect 21771 77827 21837 77828
rect 19563 75580 19629 75581
rect 19563 75516 19564 75580
rect 19628 75516 19629 75580
rect 19563 75515 19629 75516
rect 19794 57454 20414 76000
rect 21958 75717 22018 200070
rect 22878 75989 22938 202675
rect 23246 202197 23306 330923
rect 286182 325710 286242 332147
rect 286915 331260 286981 331261
rect 286915 331196 286916 331260
rect 286980 331196 286981 331260
rect 286915 331195 286981 331196
rect 286182 325650 286794 325710
rect 285443 316708 285509 316709
rect 285443 316644 285444 316708
rect 285508 316644 285509 316708
rect 285443 316643 285509 316644
rect 285446 305693 285506 316643
rect 285443 305692 285509 305693
rect 285443 305628 285444 305692
rect 285508 305628 285509 305692
rect 285443 305627 285509 305628
rect 33868 295954 34868 295986
rect 33868 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 34868 295954
rect 33868 295634 34868 295718
rect 33868 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 34868 295634
rect 33868 295366 34868 295398
rect 53868 295954 54868 295986
rect 53868 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 54868 295954
rect 53868 295634 54868 295718
rect 53868 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 54868 295634
rect 53868 295366 54868 295398
rect 73868 295954 74868 295986
rect 73868 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 74868 295954
rect 73868 295634 74868 295718
rect 73868 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 74868 295634
rect 73868 295366 74868 295398
rect 93868 295954 94868 295986
rect 93868 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 94868 295954
rect 93868 295634 94868 295718
rect 93868 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 94868 295634
rect 93868 295366 94868 295398
rect 113868 295954 114868 295986
rect 113868 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 114868 295954
rect 113868 295634 114868 295718
rect 113868 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 114868 295634
rect 113868 295366 114868 295398
rect 133868 295954 134868 295986
rect 133868 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 134868 295954
rect 133868 295634 134868 295718
rect 133868 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 134868 295634
rect 133868 295366 134868 295398
rect 153868 295954 154868 295986
rect 153868 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 154868 295954
rect 153868 295634 154868 295718
rect 153868 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 154868 295634
rect 153868 295366 154868 295398
rect 173868 295954 174868 295986
rect 173868 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 174868 295954
rect 173868 295634 174868 295718
rect 173868 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 174868 295634
rect 173868 295366 174868 295398
rect 193868 295954 194868 295986
rect 193868 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 194868 295954
rect 193868 295634 194868 295718
rect 193868 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 194868 295634
rect 193868 295366 194868 295398
rect 213868 295954 214868 295986
rect 213868 295718 213930 295954
rect 214166 295718 214250 295954
rect 214486 295718 214570 295954
rect 214806 295718 214868 295954
rect 213868 295634 214868 295718
rect 213868 295398 213930 295634
rect 214166 295398 214250 295634
rect 214486 295398 214570 295634
rect 214806 295398 214868 295634
rect 213868 295366 214868 295398
rect 233868 295954 234868 295986
rect 233868 295718 233930 295954
rect 234166 295718 234250 295954
rect 234486 295718 234570 295954
rect 234806 295718 234868 295954
rect 233868 295634 234868 295718
rect 233868 295398 233930 295634
rect 234166 295398 234250 295634
rect 234486 295398 234570 295634
rect 234806 295398 234868 295634
rect 233868 295366 234868 295398
rect 253868 295954 254868 295986
rect 253868 295718 253930 295954
rect 254166 295718 254250 295954
rect 254486 295718 254570 295954
rect 254806 295718 254868 295954
rect 253868 295634 254868 295718
rect 253868 295398 253930 295634
rect 254166 295398 254250 295634
rect 254486 295398 254570 295634
rect 254806 295398 254868 295634
rect 253868 295366 254868 295398
rect 273868 295954 274868 295986
rect 273868 295718 273930 295954
rect 274166 295718 274250 295954
rect 274486 295718 274570 295954
rect 274806 295718 274868 295954
rect 273868 295634 274868 295718
rect 273868 295398 273930 295634
rect 274166 295398 274250 295634
rect 274486 295398 274570 295634
rect 274806 295398 274868 295634
rect 273868 295366 274868 295398
rect 23868 291454 24868 291486
rect 23868 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 24868 291454
rect 23868 291134 24868 291218
rect 23868 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 24868 291134
rect 23868 290866 24868 290898
rect 43868 291454 44868 291486
rect 43868 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 44868 291454
rect 43868 291134 44868 291218
rect 43868 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 44868 291134
rect 43868 290866 44868 290898
rect 63868 291454 64868 291486
rect 63868 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 64868 291454
rect 63868 291134 64868 291218
rect 63868 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 64868 291134
rect 63868 290866 64868 290898
rect 83868 291454 84868 291486
rect 83868 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 84868 291454
rect 83868 291134 84868 291218
rect 83868 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 84868 291134
rect 83868 290866 84868 290898
rect 103868 291454 104868 291486
rect 103868 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 104868 291454
rect 103868 291134 104868 291218
rect 103868 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 104868 291134
rect 103868 290866 104868 290898
rect 123868 291454 124868 291486
rect 123868 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 124868 291454
rect 123868 291134 124868 291218
rect 123868 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 124868 291134
rect 123868 290866 124868 290898
rect 143868 291454 144868 291486
rect 143868 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 144868 291454
rect 143868 291134 144868 291218
rect 143868 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 144868 291134
rect 143868 290866 144868 290898
rect 163868 291454 164868 291486
rect 163868 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 164868 291454
rect 163868 291134 164868 291218
rect 163868 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 164868 291134
rect 163868 290866 164868 290898
rect 183868 291454 184868 291486
rect 183868 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 184868 291454
rect 183868 291134 184868 291218
rect 183868 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 184868 291134
rect 183868 290866 184868 290898
rect 203868 291454 204868 291486
rect 203868 291218 203930 291454
rect 204166 291218 204250 291454
rect 204486 291218 204570 291454
rect 204806 291218 204868 291454
rect 203868 291134 204868 291218
rect 203868 290898 203930 291134
rect 204166 290898 204250 291134
rect 204486 290898 204570 291134
rect 204806 290898 204868 291134
rect 203868 290866 204868 290898
rect 223868 291454 224868 291486
rect 223868 291218 223930 291454
rect 224166 291218 224250 291454
rect 224486 291218 224570 291454
rect 224806 291218 224868 291454
rect 223868 291134 224868 291218
rect 223868 290898 223930 291134
rect 224166 290898 224250 291134
rect 224486 290898 224570 291134
rect 224806 290898 224868 291134
rect 223868 290866 224868 290898
rect 243868 291454 244868 291486
rect 243868 291218 243930 291454
rect 244166 291218 244250 291454
rect 244486 291218 244570 291454
rect 244806 291218 244868 291454
rect 243868 291134 244868 291218
rect 243868 290898 243930 291134
rect 244166 290898 244250 291134
rect 244486 290898 244570 291134
rect 244806 290898 244868 291134
rect 243868 290866 244868 290898
rect 263868 291454 264868 291486
rect 263868 291218 263930 291454
rect 264166 291218 264250 291454
rect 264486 291218 264570 291454
rect 264806 291218 264868 291454
rect 263868 291134 264868 291218
rect 263868 290898 263930 291134
rect 264166 290898 264250 291134
rect 264486 290898 264570 291134
rect 264806 290898 264868 291134
rect 263868 290866 264868 290898
rect 283868 291454 284868 291486
rect 283868 291218 283930 291454
rect 284166 291218 284250 291454
rect 284486 291218 284570 291454
rect 284806 291218 284868 291454
rect 283868 291134 284868 291218
rect 283868 290898 283930 291134
rect 284166 290898 284250 291134
rect 284486 290898 284570 291134
rect 284806 290898 284868 291134
rect 283868 290866 284868 290898
rect 33868 259954 34868 259986
rect 33868 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 34868 259954
rect 33868 259634 34868 259718
rect 33868 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 34868 259634
rect 33868 259366 34868 259398
rect 53868 259954 54868 259986
rect 53868 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 54868 259954
rect 53868 259634 54868 259718
rect 53868 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 54868 259634
rect 53868 259366 54868 259398
rect 73868 259954 74868 259986
rect 73868 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 74868 259954
rect 73868 259634 74868 259718
rect 73868 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 74868 259634
rect 73868 259366 74868 259398
rect 93868 259954 94868 259986
rect 93868 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 94868 259954
rect 93868 259634 94868 259718
rect 93868 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 94868 259634
rect 93868 259366 94868 259398
rect 113868 259954 114868 259986
rect 113868 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 114868 259954
rect 113868 259634 114868 259718
rect 113868 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 114868 259634
rect 113868 259366 114868 259398
rect 133868 259954 134868 259986
rect 133868 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 134868 259954
rect 133868 259634 134868 259718
rect 133868 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 134868 259634
rect 133868 259366 134868 259398
rect 153868 259954 154868 259986
rect 153868 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 154868 259954
rect 153868 259634 154868 259718
rect 153868 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 154868 259634
rect 153868 259366 154868 259398
rect 173868 259954 174868 259986
rect 173868 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 174868 259954
rect 173868 259634 174868 259718
rect 173868 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 174868 259634
rect 173868 259366 174868 259398
rect 193868 259954 194868 259986
rect 193868 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 194868 259954
rect 193868 259634 194868 259718
rect 193868 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 194868 259634
rect 193868 259366 194868 259398
rect 213868 259954 214868 259986
rect 213868 259718 213930 259954
rect 214166 259718 214250 259954
rect 214486 259718 214570 259954
rect 214806 259718 214868 259954
rect 213868 259634 214868 259718
rect 213868 259398 213930 259634
rect 214166 259398 214250 259634
rect 214486 259398 214570 259634
rect 214806 259398 214868 259634
rect 213868 259366 214868 259398
rect 233868 259954 234868 259986
rect 233868 259718 233930 259954
rect 234166 259718 234250 259954
rect 234486 259718 234570 259954
rect 234806 259718 234868 259954
rect 233868 259634 234868 259718
rect 233868 259398 233930 259634
rect 234166 259398 234250 259634
rect 234486 259398 234570 259634
rect 234806 259398 234868 259634
rect 233868 259366 234868 259398
rect 253868 259954 254868 259986
rect 253868 259718 253930 259954
rect 254166 259718 254250 259954
rect 254486 259718 254570 259954
rect 254806 259718 254868 259954
rect 253868 259634 254868 259718
rect 253868 259398 253930 259634
rect 254166 259398 254250 259634
rect 254486 259398 254570 259634
rect 254806 259398 254868 259634
rect 253868 259366 254868 259398
rect 273868 259954 274868 259986
rect 273868 259718 273930 259954
rect 274166 259718 274250 259954
rect 274486 259718 274570 259954
rect 274806 259718 274868 259954
rect 273868 259634 274868 259718
rect 273868 259398 273930 259634
rect 274166 259398 274250 259634
rect 274486 259398 274570 259634
rect 274806 259398 274868 259634
rect 273868 259366 274868 259398
rect 23868 255454 24868 255486
rect 23868 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 24868 255454
rect 23868 255134 24868 255218
rect 23868 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 24868 255134
rect 23868 254866 24868 254898
rect 43868 255454 44868 255486
rect 43868 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 44868 255454
rect 43868 255134 44868 255218
rect 43868 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 44868 255134
rect 43868 254866 44868 254898
rect 63868 255454 64868 255486
rect 63868 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 64868 255454
rect 63868 255134 64868 255218
rect 63868 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 64868 255134
rect 63868 254866 64868 254898
rect 83868 255454 84868 255486
rect 83868 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 84868 255454
rect 83868 255134 84868 255218
rect 83868 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 84868 255134
rect 83868 254866 84868 254898
rect 103868 255454 104868 255486
rect 103868 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 104868 255454
rect 103868 255134 104868 255218
rect 103868 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 104868 255134
rect 103868 254866 104868 254898
rect 123868 255454 124868 255486
rect 123868 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 124868 255454
rect 123868 255134 124868 255218
rect 123868 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 124868 255134
rect 123868 254866 124868 254898
rect 143868 255454 144868 255486
rect 143868 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 144868 255454
rect 143868 255134 144868 255218
rect 143868 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 144868 255134
rect 143868 254866 144868 254898
rect 163868 255454 164868 255486
rect 163868 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 164868 255454
rect 163868 255134 164868 255218
rect 163868 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 164868 255134
rect 163868 254866 164868 254898
rect 183868 255454 184868 255486
rect 183868 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 184868 255454
rect 183868 255134 184868 255218
rect 183868 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 184868 255134
rect 183868 254866 184868 254898
rect 203868 255454 204868 255486
rect 203868 255218 203930 255454
rect 204166 255218 204250 255454
rect 204486 255218 204570 255454
rect 204806 255218 204868 255454
rect 203868 255134 204868 255218
rect 203868 254898 203930 255134
rect 204166 254898 204250 255134
rect 204486 254898 204570 255134
rect 204806 254898 204868 255134
rect 203868 254866 204868 254898
rect 223868 255454 224868 255486
rect 223868 255218 223930 255454
rect 224166 255218 224250 255454
rect 224486 255218 224570 255454
rect 224806 255218 224868 255454
rect 223868 255134 224868 255218
rect 223868 254898 223930 255134
rect 224166 254898 224250 255134
rect 224486 254898 224570 255134
rect 224806 254898 224868 255134
rect 223868 254866 224868 254898
rect 243868 255454 244868 255486
rect 243868 255218 243930 255454
rect 244166 255218 244250 255454
rect 244486 255218 244570 255454
rect 244806 255218 244868 255454
rect 243868 255134 244868 255218
rect 243868 254898 243930 255134
rect 244166 254898 244250 255134
rect 244486 254898 244570 255134
rect 244806 254898 244868 255134
rect 243868 254866 244868 254898
rect 263868 255454 264868 255486
rect 263868 255218 263930 255454
rect 264166 255218 264250 255454
rect 264486 255218 264570 255454
rect 264806 255218 264868 255454
rect 263868 255134 264868 255218
rect 263868 254898 263930 255134
rect 264166 254898 264250 255134
rect 264486 254898 264570 255134
rect 264806 254898 264868 255134
rect 263868 254866 264868 254898
rect 283868 255454 284868 255486
rect 283868 255218 283930 255454
rect 284166 255218 284250 255454
rect 284486 255218 284570 255454
rect 284806 255218 284868 255454
rect 283868 255134 284868 255218
rect 283868 254898 283930 255134
rect 284166 254898 284250 255134
rect 284486 254898 284570 255134
rect 284806 254898 284868 255134
rect 283868 254866 284868 254898
rect 33868 223954 34868 223986
rect 33868 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 34868 223954
rect 33868 223634 34868 223718
rect 33868 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 34868 223634
rect 33868 223366 34868 223398
rect 53868 223954 54868 223986
rect 53868 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 54868 223954
rect 53868 223634 54868 223718
rect 53868 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 54868 223634
rect 53868 223366 54868 223398
rect 73868 223954 74868 223986
rect 73868 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 74868 223954
rect 73868 223634 74868 223718
rect 73868 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 74868 223634
rect 73868 223366 74868 223398
rect 93868 223954 94868 223986
rect 93868 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 94868 223954
rect 93868 223634 94868 223718
rect 93868 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 94868 223634
rect 93868 223366 94868 223398
rect 113868 223954 114868 223986
rect 113868 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 114868 223954
rect 113868 223634 114868 223718
rect 113868 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 114868 223634
rect 113868 223366 114868 223398
rect 133868 223954 134868 223986
rect 133868 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 134868 223954
rect 133868 223634 134868 223718
rect 133868 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 134868 223634
rect 133868 223366 134868 223398
rect 153868 223954 154868 223986
rect 153868 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 154868 223954
rect 153868 223634 154868 223718
rect 153868 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 154868 223634
rect 153868 223366 154868 223398
rect 173868 223954 174868 223986
rect 173868 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 174868 223954
rect 173868 223634 174868 223718
rect 173868 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 174868 223634
rect 173868 223366 174868 223398
rect 193868 223954 194868 223986
rect 193868 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 194868 223954
rect 193868 223634 194868 223718
rect 193868 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 194868 223634
rect 193868 223366 194868 223398
rect 213868 223954 214868 223986
rect 213868 223718 213930 223954
rect 214166 223718 214250 223954
rect 214486 223718 214570 223954
rect 214806 223718 214868 223954
rect 213868 223634 214868 223718
rect 213868 223398 213930 223634
rect 214166 223398 214250 223634
rect 214486 223398 214570 223634
rect 214806 223398 214868 223634
rect 213868 223366 214868 223398
rect 233868 223954 234868 223986
rect 233868 223718 233930 223954
rect 234166 223718 234250 223954
rect 234486 223718 234570 223954
rect 234806 223718 234868 223954
rect 233868 223634 234868 223718
rect 233868 223398 233930 223634
rect 234166 223398 234250 223634
rect 234486 223398 234570 223634
rect 234806 223398 234868 223634
rect 233868 223366 234868 223398
rect 253868 223954 254868 223986
rect 253868 223718 253930 223954
rect 254166 223718 254250 223954
rect 254486 223718 254570 223954
rect 254806 223718 254868 223954
rect 253868 223634 254868 223718
rect 253868 223398 253930 223634
rect 254166 223398 254250 223634
rect 254486 223398 254570 223634
rect 254806 223398 254868 223634
rect 253868 223366 254868 223398
rect 273868 223954 274868 223986
rect 273868 223718 273930 223954
rect 274166 223718 274250 223954
rect 274486 223718 274570 223954
rect 274806 223718 274868 223954
rect 273868 223634 274868 223718
rect 273868 223398 273930 223634
rect 274166 223398 274250 223634
rect 274486 223398 274570 223634
rect 274806 223398 274868 223634
rect 273868 223366 274868 223398
rect 23868 219454 24868 219486
rect 23868 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 24868 219454
rect 23868 219134 24868 219218
rect 23868 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 24868 219134
rect 23868 218866 24868 218898
rect 43868 219454 44868 219486
rect 43868 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 44868 219454
rect 43868 219134 44868 219218
rect 43868 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 44868 219134
rect 43868 218866 44868 218898
rect 63868 219454 64868 219486
rect 63868 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 64868 219454
rect 63868 219134 64868 219218
rect 63868 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 64868 219134
rect 63868 218866 64868 218898
rect 83868 219454 84868 219486
rect 83868 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 84868 219454
rect 83868 219134 84868 219218
rect 83868 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 84868 219134
rect 83868 218866 84868 218898
rect 103868 219454 104868 219486
rect 103868 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 104868 219454
rect 103868 219134 104868 219218
rect 103868 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 104868 219134
rect 103868 218866 104868 218898
rect 123868 219454 124868 219486
rect 123868 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 124868 219454
rect 123868 219134 124868 219218
rect 123868 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 124868 219134
rect 123868 218866 124868 218898
rect 143868 219454 144868 219486
rect 143868 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 144868 219454
rect 143868 219134 144868 219218
rect 143868 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 144868 219134
rect 143868 218866 144868 218898
rect 163868 219454 164868 219486
rect 163868 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 164868 219454
rect 163868 219134 164868 219218
rect 163868 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 164868 219134
rect 163868 218866 164868 218898
rect 183868 219454 184868 219486
rect 183868 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 184868 219454
rect 183868 219134 184868 219218
rect 183868 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 184868 219134
rect 183868 218866 184868 218898
rect 203868 219454 204868 219486
rect 203868 219218 203930 219454
rect 204166 219218 204250 219454
rect 204486 219218 204570 219454
rect 204806 219218 204868 219454
rect 203868 219134 204868 219218
rect 203868 218898 203930 219134
rect 204166 218898 204250 219134
rect 204486 218898 204570 219134
rect 204806 218898 204868 219134
rect 203868 218866 204868 218898
rect 223868 219454 224868 219486
rect 223868 219218 223930 219454
rect 224166 219218 224250 219454
rect 224486 219218 224570 219454
rect 224806 219218 224868 219454
rect 223868 219134 224868 219218
rect 223868 218898 223930 219134
rect 224166 218898 224250 219134
rect 224486 218898 224570 219134
rect 224806 218898 224868 219134
rect 223868 218866 224868 218898
rect 243868 219454 244868 219486
rect 243868 219218 243930 219454
rect 244166 219218 244250 219454
rect 244486 219218 244570 219454
rect 244806 219218 244868 219454
rect 243868 219134 244868 219218
rect 243868 218898 243930 219134
rect 244166 218898 244250 219134
rect 244486 218898 244570 219134
rect 244806 218898 244868 219134
rect 243868 218866 244868 218898
rect 263868 219454 264868 219486
rect 263868 219218 263930 219454
rect 264166 219218 264250 219454
rect 264486 219218 264570 219454
rect 264806 219218 264868 219454
rect 263868 219134 264868 219218
rect 263868 218898 263930 219134
rect 264166 218898 264250 219134
rect 264486 218898 264570 219134
rect 264806 218898 264868 219134
rect 263868 218866 264868 218898
rect 283868 219454 284868 219486
rect 283868 219218 283930 219454
rect 284166 219218 284250 219454
rect 284486 219218 284570 219454
rect 284806 219218 284868 219454
rect 283868 219134 284868 219218
rect 283868 218898 283930 219134
rect 284166 218898 284250 219134
rect 284486 218898 284570 219134
rect 284806 218898 284868 219134
rect 283868 218866 284868 218898
rect 286734 203693 286794 325650
rect 286731 203692 286797 203693
rect 286731 203628 286732 203692
rect 286796 203628 286797 203692
rect 286731 203627 286797 203628
rect 23243 202196 23309 202197
rect 23243 202132 23244 202196
rect 23308 202132 23309 202196
rect 23243 202131 23309 202132
rect 285259 188324 285325 188325
rect 285259 188260 285260 188324
rect 285324 188260 285325 188324
rect 285259 188259 285325 188260
rect 23059 186420 23125 186421
rect 23059 186356 23060 186420
rect 23124 186356 23125 186420
rect 23059 186355 23125 186356
rect 22875 75988 22941 75989
rect 22875 75924 22876 75988
rect 22940 75924 22941 75988
rect 22875 75923 22941 75924
rect 23062 75853 23122 186355
rect 23868 183454 24868 183486
rect 23868 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 24868 183454
rect 23868 183134 24868 183218
rect 23868 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 24868 183134
rect 23868 182866 24868 182898
rect 43868 183454 44868 183486
rect 43868 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 44868 183454
rect 43868 183134 44868 183218
rect 43868 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 44868 183134
rect 43868 182866 44868 182898
rect 63868 183454 64868 183486
rect 63868 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 64868 183454
rect 63868 183134 64868 183218
rect 63868 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 64868 183134
rect 63868 182866 64868 182898
rect 83868 183454 84868 183486
rect 83868 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 84868 183454
rect 83868 183134 84868 183218
rect 83868 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 84868 183134
rect 83868 182866 84868 182898
rect 103868 183454 104868 183486
rect 103868 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 104868 183454
rect 103868 183134 104868 183218
rect 103868 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 104868 183134
rect 103868 182866 104868 182898
rect 123868 183454 124868 183486
rect 123868 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 124868 183454
rect 123868 183134 124868 183218
rect 123868 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 124868 183134
rect 123868 182866 124868 182898
rect 143868 183454 144868 183486
rect 143868 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 144868 183454
rect 143868 183134 144868 183218
rect 143868 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 144868 183134
rect 143868 182866 144868 182898
rect 163868 183454 164868 183486
rect 163868 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 164868 183454
rect 163868 183134 164868 183218
rect 163868 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 164868 183134
rect 163868 182866 164868 182898
rect 183868 183454 184868 183486
rect 183868 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 184868 183454
rect 183868 183134 184868 183218
rect 183868 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 184868 183134
rect 183868 182866 184868 182898
rect 203868 183454 204868 183486
rect 203868 183218 203930 183454
rect 204166 183218 204250 183454
rect 204486 183218 204570 183454
rect 204806 183218 204868 183454
rect 203868 183134 204868 183218
rect 203868 182898 203930 183134
rect 204166 182898 204250 183134
rect 204486 182898 204570 183134
rect 204806 182898 204868 183134
rect 203868 182866 204868 182898
rect 223868 183454 224868 183486
rect 223868 183218 223930 183454
rect 224166 183218 224250 183454
rect 224486 183218 224570 183454
rect 224806 183218 224868 183454
rect 223868 183134 224868 183218
rect 223868 182898 223930 183134
rect 224166 182898 224250 183134
rect 224486 182898 224570 183134
rect 224806 182898 224868 183134
rect 223868 182866 224868 182898
rect 243868 183454 244868 183486
rect 243868 183218 243930 183454
rect 244166 183218 244250 183454
rect 244486 183218 244570 183454
rect 244806 183218 244868 183454
rect 243868 183134 244868 183218
rect 243868 182898 243930 183134
rect 244166 182898 244250 183134
rect 244486 182898 244570 183134
rect 244806 182898 244868 183134
rect 243868 182866 244868 182898
rect 263868 183454 264868 183486
rect 263868 183218 263930 183454
rect 264166 183218 264250 183454
rect 264486 183218 264570 183454
rect 264806 183218 264868 183454
rect 263868 183134 264868 183218
rect 263868 182898 263930 183134
rect 264166 182898 264250 183134
rect 264486 182898 264570 183134
rect 264806 182898 264868 183134
rect 263868 182866 264868 182898
rect 283868 183454 284868 183486
rect 283868 183218 283930 183454
rect 284166 183218 284250 183454
rect 284486 183218 284570 183454
rect 284806 183218 284868 183454
rect 283868 183134 284868 183218
rect 283868 182898 283930 183134
rect 284166 182898 284250 183134
rect 284486 182898 284570 183134
rect 284806 182898 284868 183134
rect 283868 182866 284868 182898
rect 285262 177989 285322 188259
rect 286179 186148 286245 186149
rect 286179 186084 286180 186148
rect 286244 186084 286245 186148
rect 286179 186083 286245 186084
rect 285259 177988 285325 177989
rect 285259 177924 285260 177988
rect 285324 177924 285325 177988
rect 285259 177923 285325 177924
rect 33868 151954 34868 151986
rect 33868 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 34868 151954
rect 33868 151634 34868 151718
rect 33868 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 34868 151634
rect 33868 151366 34868 151398
rect 53868 151954 54868 151986
rect 53868 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 54868 151954
rect 53868 151634 54868 151718
rect 53868 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 54868 151634
rect 53868 151366 54868 151398
rect 73868 151954 74868 151986
rect 73868 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 74868 151954
rect 73868 151634 74868 151718
rect 73868 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 74868 151634
rect 73868 151366 74868 151398
rect 93868 151954 94868 151986
rect 93868 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 94868 151954
rect 93868 151634 94868 151718
rect 93868 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 94868 151634
rect 93868 151366 94868 151398
rect 113868 151954 114868 151986
rect 113868 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 114868 151954
rect 113868 151634 114868 151718
rect 113868 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 114868 151634
rect 113868 151366 114868 151398
rect 133868 151954 134868 151986
rect 133868 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 134868 151954
rect 133868 151634 134868 151718
rect 133868 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 134868 151634
rect 133868 151366 134868 151398
rect 153868 151954 154868 151986
rect 153868 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 154868 151954
rect 153868 151634 154868 151718
rect 153868 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 154868 151634
rect 153868 151366 154868 151398
rect 173868 151954 174868 151986
rect 173868 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 174868 151954
rect 173868 151634 174868 151718
rect 173868 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 174868 151634
rect 173868 151366 174868 151398
rect 193868 151954 194868 151986
rect 193868 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 194868 151954
rect 193868 151634 194868 151718
rect 193868 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 194868 151634
rect 193868 151366 194868 151398
rect 213868 151954 214868 151986
rect 213868 151718 213930 151954
rect 214166 151718 214250 151954
rect 214486 151718 214570 151954
rect 214806 151718 214868 151954
rect 213868 151634 214868 151718
rect 213868 151398 213930 151634
rect 214166 151398 214250 151634
rect 214486 151398 214570 151634
rect 214806 151398 214868 151634
rect 213868 151366 214868 151398
rect 233868 151954 234868 151986
rect 233868 151718 233930 151954
rect 234166 151718 234250 151954
rect 234486 151718 234570 151954
rect 234806 151718 234868 151954
rect 233868 151634 234868 151718
rect 233868 151398 233930 151634
rect 234166 151398 234250 151634
rect 234486 151398 234570 151634
rect 234806 151398 234868 151634
rect 233868 151366 234868 151398
rect 253868 151954 254868 151986
rect 253868 151718 253930 151954
rect 254166 151718 254250 151954
rect 254486 151718 254570 151954
rect 254806 151718 254868 151954
rect 253868 151634 254868 151718
rect 253868 151398 253930 151634
rect 254166 151398 254250 151634
rect 254486 151398 254570 151634
rect 254806 151398 254868 151634
rect 253868 151366 254868 151398
rect 273868 151954 274868 151986
rect 273868 151718 273930 151954
rect 274166 151718 274250 151954
rect 274486 151718 274570 151954
rect 274806 151718 274868 151954
rect 273868 151634 274868 151718
rect 273868 151398 273930 151634
rect 274166 151398 274250 151634
rect 274486 151398 274570 151634
rect 274806 151398 274868 151634
rect 273868 151366 274868 151398
rect 23868 147454 24868 147486
rect 23868 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 24868 147454
rect 23868 147134 24868 147218
rect 23868 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 24868 147134
rect 23868 146866 24868 146898
rect 43868 147454 44868 147486
rect 43868 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 44868 147454
rect 43868 147134 44868 147218
rect 43868 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 44868 147134
rect 43868 146866 44868 146898
rect 63868 147454 64868 147486
rect 63868 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 64868 147454
rect 63868 147134 64868 147218
rect 63868 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 64868 147134
rect 63868 146866 64868 146898
rect 83868 147454 84868 147486
rect 83868 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 84868 147454
rect 83868 147134 84868 147218
rect 83868 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 84868 147134
rect 83868 146866 84868 146898
rect 103868 147454 104868 147486
rect 103868 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 104868 147454
rect 103868 147134 104868 147218
rect 103868 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 104868 147134
rect 103868 146866 104868 146898
rect 123868 147454 124868 147486
rect 123868 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 124868 147454
rect 123868 147134 124868 147218
rect 123868 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 124868 147134
rect 123868 146866 124868 146898
rect 143868 147454 144868 147486
rect 143868 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 144868 147454
rect 143868 147134 144868 147218
rect 143868 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 144868 147134
rect 143868 146866 144868 146898
rect 163868 147454 164868 147486
rect 163868 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 164868 147454
rect 163868 147134 164868 147218
rect 163868 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 164868 147134
rect 163868 146866 164868 146898
rect 183868 147454 184868 147486
rect 183868 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 184868 147454
rect 183868 147134 184868 147218
rect 183868 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 184868 147134
rect 183868 146866 184868 146898
rect 203868 147454 204868 147486
rect 203868 147218 203930 147454
rect 204166 147218 204250 147454
rect 204486 147218 204570 147454
rect 204806 147218 204868 147454
rect 203868 147134 204868 147218
rect 203868 146898 203930 147134
rect 204166 146898 204250 147134
rect 204486 146898 204570 147134
rect 204806 146898 204868 147134
rect 203868 146866 204868 146898
rect 223868 147454 224868 147486
rect 223868 147218 223930 147454
rect 224166 147218 224250 147454
rect 224486 147218 224570 147454
rect 224806 147218 224868 147454
rect 223868 147134 224868 147218
rect 223868 146898 223930 147134
rect 224166 146898 224250 147134
rect 224486 146898 224570 147134
rect 224806 146898 224868 147134
rect 223868 146866 224868 146898
rect 243868 147454 244868 147486
rect 243868 147218 243930 147454
rect 244166 147218 244250 147454
rect 244486 147218 244570 147454
rect 244806 147218 244868 147454
rect 243868 147134 244868 147218
rect 243868 146898 243930 147134
rect 244166 146898 244250 147134
rect 244486 146898 244570 147134
rect 244806 146898 244868 147134
rect 243868 146866 244868 146898
rect 263868 147454 264868 147486
rect 263868 147218 263930 147454
rect 264166 147218 264250 147454
rect 264486 147218 264570 147454
rect 264806 147218 264868 147454
rect 263868 147134 264868 147218
rect 263868 146898 263930 147134
rect 264166 146898 264250 147134
rect 264486 146898 264570 147134
rect 264806 146898 264868 147134
rect 263868 146866 264868 146898
rect 283868 147454 284868 147486
rect 283868 147218 283930 147454
rect 284166 147218 284250 147454
rect 284486 147218 284570 147454
rect 284806 147218 284868 147454
rect 283868 147134 284868 147218
rect 283868 146898 283930 147134
rect 284166 146898 284250 147134
rect 284486 146898 284570 147134
rect 284806 146898 284868 147134
rect 283868 146866 284868 146898
rect 33868 115954 34868 115986
rect 33868 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 34868 115954
rect 33868 115634 34868 115718
rect 33868 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 34868 115634
rect 33868 115366 34868 115398
rect 53868 115954 54868 115986
rect 53868 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 54868 115954
rect 53868 115634 54868 115718
rect 53868 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 54868 115634
rect 53868 115366 54868 115398
rect 73868 115954 74868 115986
rect 73868 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 74868 115954
rect 73868 115634 74868 115718
rect 73868 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 74868 115634
rect 73868 115366 74868 115398
rect 93868 115954 94868 115986
rect 93868 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 94868 115954
rect 93868 115634 94868 115718
rect 93868 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 94868 115634
rect 93868 115366 94868 115398
rect 113868 115954 114868 115986
rect 113868 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 114868 115954
rect 113868 115634 114868 115718
rect 113868 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 114868 115634
rect 113868 115366 114868 115398
rect 133868 115954 134868 115986
rect 133868 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 134868 115954
rect 133868 115634 134868 115718
rect 133868 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 134868 115634
rect 133868 115366 134868 115398
rect 153868 115954 154868 115986
rect 153868 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 154868 115954
rect 153868 115634 154868 115718
rect 153868 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 154868 115634
rect 153868 115366 154868 115398
rect 173868 115954 174868 115986
rect 173868 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 174868 115954
rect 173868 115634 174868 115718
rect 173868 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 174868 115634
rect 173868 115366 174868 115398
rect 193868 115954 194868 115986
rect 193868 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 194868 115954
rect 193868 115634 194868 115718
rect 193868 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 194868 115634
rect 193868 115366 194868 115398
rect 213868 115954 214868 115986
rect 213868 115718 213930 115954
rect 214166 115718 214250 115954
rect 214486 115718 214570 115954
rect 214806 115718 214868 115954
rect 213868 115634 214868 115718
rect 213868 115398 213930 115634
rect 214166 115398 214250 115634
rect 214486 115398 214570 115634
rect 214806 115398 214868 115634
rect 213868 115366 214868 115398
rect 233868 115954 234868 115986
rect 233868 115718 233930 115954
rect 234166 115718 234250 115954
rect 234486 115718 234570 115954
rect 234806 115718 234868 115954
rect 233868 115634 234868 115718
rect 233868 115398 233930 115634
rect 234166 115398 234250 115634
rect 234486 115398 234570 115634
rect 234806 115398 234868 115634
rect 233868 115366 234868 115398
rect 253868 115954 254868 115986
rect 253868 115718 253930 115954
rect 254166 115718 254250 115954
rect 254486 115718 254570 115954
rect 254806 115718 254868 115954
rect 253868 115634 254868 115718
rect 253868 115398 253930 115634
rect 254166 115398 254250 115634
rect 254486 115398 254570 115634
rect 254806 115398 254868 115634
rect 253868 115366 254868 115398
rect 273868 115954 274868 115986
rect 273868 115718 273930 115954
rect 274166 115718 274250 115954
rect 274486 115718 274570 115954
rect 274806 115718 274868 115954
rect 273868 115634 274868 115718
rect 273868 115398 273930 115634
rect 274166 115398 274250 115634
rect 274486 115398 274570 115634
rect 274806 115398 274868 115634
rect 273868 115366 274868 115398
rect 23868 111454 24868 111486
rect 23868 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 24868 111454
rect 23868 111134 24868 111218
rect 23868 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 24868 111134
rect 23868 110866 24868 110898
rect 43868 111454 44868 111486
rect 43868 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 44868 111454
rect 43868 111134 44868 111218
rect 43868 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 44868 111134
rect 43868 110866 44868 110898
rect 63868 111454 64868 111486
rect 63868 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 64868 111454
rect 63868 111134 64868 111218
rect 63868 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 64868 111134
rect 63868 110866 64868 110898
rect 83868 111454 84868 111486
rect 83868 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 84868 111454
rect 83868 111134 84868 111218
rect 83868 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 84868 111134
rect 83868 110866 84868 110898
rect 103868 111454 104868 111486
rect 103868 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 104868 111454
rect 103868 111134 104868 111218
rect 103868 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 104868 111134
rect 103868 110866 104868 110898
rect 123868 111454 124868 111486
rect 123868 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 124868 111454
rect 123868 111134 124868 111218
rect 123868 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 124868 111134
rect 123868 110866 124868 110898
rect 143868 111454 144868 111486
rect 143868 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 144868 111454
rect 143868 111134 144868 111218
rect 143868 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 144868 111134
rect 143868 110866 144868 110898
rect 163868 111454 164868 111486
rect 163868 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 164868 111454
rect 163868 111134 164868 111218
rect 163868 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 164868 111134
rect 163868 110866 164868 110898
rect 183868 111454 184868 111486
rect 183868 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 184868 111454
rect 183868 111134 184868 111218
rect 183868 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 184868 111134
rect 183868 110866 184868 110898
rect 203868 111454 204868 111486
rect 203868 111218 203930 111454
rect 204166 111218 204250 111454
rect 204486 111218 204570 111454
rect 204806 111218 204868 111454
rect 203868 111134 204868 111218
rect 203868 110898 203930 111134
rect 204166 110898 204250 111134
rect 204486 110898 204570 111134
rect 204806 110898 204868 111134
rect 203868 110866 204868 110898
rect 223868 111454 224868 111486
rect 223868 111218 223930 111454
rect 224166 111218 224250 111454
rect 224486 111218 224570 111454
rect 224806 111218 224868 111454
rect 223868 111134 224868 111218
rect 223868 110898 223930 111134
rect 224166 110898 224250 111134
rect 224486 110898 224570 111134
rect 224806 110898 224868 111134
rect 223868 110866 224868 110898
rect 243868 111454 244868 111486
rect 243868 111218 243930 111454
rect 244166 111218 244250 111454
rect 244486 111218 244570 111454
rect 244806 111218 244868 111454
rect 243868 111134 244868 111218
rect 243868 110898 243930 111134
rect 244166 110898 244250 111134
rect 244486 110898 244570 111134
rect 244806 110898 244868 111134
rect 243868 110866 244868 110898
rect 263868 111454 264868 111486
rect 263868 111218 263930 111454
rect 264166 111218 264250 111454
rect 264486 111218 264570 111454
rect 264806 111218 264868 111454
rect 263868 111134 264868 111218
rect 263868 110898 263930 111134
rect 264166 110898 264250 111134
rect 264486 110898 264570 111134
rect 264806 110898 264868 111134
rect 263868 110866 264868 110898
rect 283868 111454 284868 111486
rect 283868 111218 283930 111454
rect 284166 111218 284250 111454
rect 284486 111218 284570 111454
rect 284806 111218 284868 111454
rect 283868 111134 284868 111218
rect 283868 110898 283930 111134
rect 284166 110898 284250 111134
rect 284486 110898 284570 111134
rect 284806 110898 284868 111134
rect 283868 110866 284868 110898
rect 23059 75852 23125 75853
rect 23059 75788 23060 75852
rect 23124 75788 23125 75852
rect 23059 75787 23125 75788
rect 21955 75716 22021 75717
rect 21955 75652 21956 75716
rect 22020 75652 22021 75716
rect 21955 75651 22021 75652
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19195 34644 19261 34645
rect 19195 34580 19196 34644
rect 19260 34580 19261 34644
rect 19195 34579 19261 34580
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 61954 24914 76000
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 66454 29414 76000
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 70954 33914 76000
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 75454 38414 76000
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 43954 42914 76000
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 48454 47414 76000
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 52954 51914 76000
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 76000
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 61954 60914 76000
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 66454 65414 76000
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 76000
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 76000
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 43954 78914 76000
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 48454 83414 76000
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 52954 87914 76000
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 76000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 76000
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 76000
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 76000
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 76000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 76000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 76000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 76000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 76000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 76000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 76000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 76000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 76000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 76000
rect 286182 53957 286242 186083
rect 286918 57221 286978 331195
rect 287654 76533 287714 699755
rect 288203 570620 288269 570621
rect 288203 570556 288204 570620
rect 288268 570556 288269 570620
rect 288203 570555 288269 570556
rect 287651 76532 287717 76533
rect 287651 76468 287652 76532
rect 287716 76468 287717 76532
rect 287651 76467 287717 76468
rect 286915 57220 286981 57221
rect 286915 57156 286916 57220
rect 286980 57156 286981 57220
rect 286915 57155 286981 57156
rect 288206 54909 288266 570555
rect 288203 54908 288269 54909
rect 288203 54844 288204 54908
rect 288268 54844 288269 54908
rect 288203 54843 288269 54844
rect 286179 53956 286245 53957
rect 286179 53892 286180 53956
rect 286244 53892 286245 53956
rect 286179 53891 286245 53892
rect 288942 53141 289002 700299
rect 294294 691954 294914 705242
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 700000 303914 700398
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 700000 339914 700398
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 700000 375914 700398
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 700000 411914 700398
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 700000 447914 700398
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 700000 483914 700398
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 700000 519914 700398
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 700000 555914 700398
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 303475 697508 303541 697509
rect 303475 697444 303476 697508
rect 303540 697444 303541 697508
rect 303475 697443 303541 697444
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 292619 585852 292685 585853
rect 292619 585788 292620 585852
rect 292684 585788 292685 585852
rect 292619 585787 292685 585788
rect 292435 585716 292501 585717
rect 292435 585652 292436 585716
rect 292500 585652 292501 585716
rect 292435 585651 292501 585652
rect 290043 580276 290109 580277
rect 290043 580212 290044 580276
rect 290108 580212 290109 580276
rect 290043 580211 290109 580212
rect 290046 460189 290106 580211
rect 290043 460188 290109 460189
rect 290043 460124 290044 460188
rect 290108 460124 290109 460188
rect 290043 460123 290109 460124
rect 289859 459644 289925 459645
rect 289859 459580 289860 459644
rect 289924 459580 289925 459644
rect 289859 459579 289925 459580
rect 289123 443596 289189 443597
rect 289123 443532 289124 443596
rect 289188 443532 289189 443596
rect 289123 443531 289189 443532
rect 289126 54501 289186 443531
rect 289862 332485 289922 459579
rect 290043 443868 290109 443869
rect 290043 443804 290044 443868
rect 290108 443804 290109 443868
rect 290043 443803 290109 443804
rect 289859 332484 289925 332485
rect 289859 332420 289860 332484
rect 289924 332420 289925 332484
rect 289859 332419 289925 332420
rect 289859 331804 289925 331805
rect 289859 331740 289860 331804
rect 289924 331740 289925 331804
rect 289859 331739 289925 331740
rect 289862 54637 289922 331739
rect 290046 316709 290106 443803
rect 291147 443732 291213 443733
rect 291147 443668 291148 443732
rect 291212 443668 291213 443732
rect 291147 443667 291213 443668
rect 290043 316708 290109 316709
rect 290043 316644 290044 316708
rect 290108 316644 290109 316708
rect 290043 316643 290109 316644
rect 290043 315348 290109 315349
rect 290043 315284 290044 315348
rect 290108 315284 290109 315348
rect 290043 315283 290109 315284
rect 290046 57357 290106 315283
rect 291150 57493 291210 443667
rect 292438 76397 292498 585651
rect 292435 76396 292501 76397
rect 292435 76332 292436 76396
rect 292500 76332 292501 76396
rect 292435 76331 292501 76332
rect 291147 57492 291213 57493
rect 291147 57428 291148 57492
rect 291212 57428 291213 57492
rect 291147 57427 291213 57428
rect 290043 57356 290109 57357
rect 290043 57292 290044 57356
rect 290108 57292 290109 57356
rect 290043 57291 290109 57292
rect 292622 54773 292682 585787
rect 294294 583954 294914 619398
rect 297955 585852 298021 585853
rect 297955 585788 297956 585852
rect 298020 585788 298021 585852
rect 297955 585787 298021 585788
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 292803 571980 292869 571981
rect 292803 571916 292804 571980
rect 292868 571916 292869 571980
rect 292803 571915 292869 571916
rect 292806 59941 292866 571915
rect 294294 547954 294914 583398
rect 295931 572116 295997 572117
rect 295931 572052 295932 572116
rect 295996 572052 295997 572116
rect 295931 572051 295997 572052
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 295011 458828 295077 458829
rect 295011 458764 295012 458828
rect 295076 458764 295077 458828
rect 295011 458763 295077 458764
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 292803 59940 292869 59941
rect 292803 59876 292804 59940
rect 292868 59876 292869 59940
rect 292803 59875 292869 59876
rect 292619 54772 292685 54773
rect 292619 54708 292620 54772
rect 292684 54708 292685 54772
rect 292619 54707 292685 54708
rect 289859 54636 289925 54637
rect 289859 54572 289860 54636
rect 289924 54572 289925 54636
rect 289859 54571 289925 54572
rect 289123 54500 289189 54501
rect 289123 54436 289124 54500
rect 289188 54436 289189 54500
rect 289123 54435 289189 54436
rect 294294 54000 294914 79398
rect 295014 76805 295074 458763
rect 295011 76804 295077 76805
rect 295011 76740 295012 76804
rect 295076 76740 295077 76804
rect 295011 76739 295077 76740
rect 295934 59941 295994 572051
rect 297771 444004 297837 444005
rect 297771 443940 297772 444004
rect 297836 443940 297837 444004
rect 297771 443939 297837 443940
rect 296115 329084 296181 329085
rect 296115 329020 296116 329084
rect 296180 329020 296181 329084
rect 296115 329019 296181 329020
rect 296118 73813 296178 329019
rect 296115 73812 296181 73813
rect 296115 73748 296116 73812
rect 296180 73748 296181 73812
rect 296115 73747 296181 73748
rect 295931 59940 295997 59941
rect 295931 59876 295932 59940
rect 295996 59876 295997 59940
rect 295931 59875 295997 59876
rect 297774 57357 297834 443939
rect 297958 76941 298018 585787
rect 301635 580276 301701 580277
rect 301635 580212 301636 580276
rect 301700 580212 301701 580276
rect 301635 580211 301701 580212
rect 301638 459509 301698 580211
rect 302187 571980 302253 571981
rect 302187 571916 302188 571980
rect 302252 571916 302253 571980
rect 302187 571915 302253 571916
rect 302190 547890 302250 571915
rect 302006 547830 302250 547890
rect 302006 461821 302066 547830
rect 303478 461957 303538 697443
rect 313868 691954 314868 691986
rect 313868 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 314868 691954
rect 313868 691634 314868 691718
rect 313868 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 314868 691634
rect 313868 691366 314868 691398
rect 333868 691954 334868 691986
rect 333868 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 334868 691954
rect 333868 691634 334868 691718
rect 333868 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 334868 691634
rect 333868 691366 334868 691398
rect 353868 691954 354868 691986
rect 353868 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 354868 691954
rect 353868 691634 354868 691718
rect 353868 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 354868 691634
rect 353868 691366 354868 691398
rect 373868 691954 374868 691986
rect 373868 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 374868 691954
rect 373868 691634 374868 691718
rect 373868 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 374868 691634
rect 373868 691366 374868 691398
rect 393868 691954 394868 691986
rect 393868 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 394868 691954
rect 393868 691634 394868 691718
rect 393868 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 394868 691634
rect 393868 691366 394868 691398
rect 413868 691954 414868 691986
rect 413868 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 414868 691954
rect 413868 691634 414868 691718
rect 413868 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 414868 691634
rect 413868 691366 414868 691398
rect 433868 691954 434868 691986
rect 433868 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 434868 691954
rect 433868 691634 434868 691718
rect 433868 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 434868 691634
rect 433868 691366 434868 691398
rect 453868 691954 454868 691986
rect 453868 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 454868 691954
rect 453868 691634 454868 691718
rect 453868 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 454868 691634
rect 453868 691366 454868 691398
rect 473868 691954 474868 691986
rect 473868 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 474868 691954
rect 473868 691634 474868 691718
rect 473868 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 474868 691634
rect 473868 691366 474868 691398
rect 493868 691954 494868 691986
rect 493868 691718 493930 691954
rect 494166 691718 494250 691954
rect 494486 691718 494570 691954
rect 494806 691718 494868 691954
rect 493868 691634 494868 691718
rect 493868 691398 493930 691634
rect 494166 691398 494250 691634
rect 494486 691398 494570 691634
rect 494806 691398 494868 691634
rect 493868 691366 494868 691398
rect 513868 691954 514868 691986
rect 513868 691718 513930 691954
rect 514166 691718 514250 691954
rect 514486 691718 514570 691954
rect 514806 691718 514868 691954
rect 513868 691634 514868 691718
rect 513868 691398 513930 691634
rect 514166 691398 514250 691634
rect 514486 691398 514570 691634
rect 514806 691398 514868 691634
rect 513868 691366 514868 691398
rect 533868 691954 534868 691986
rect 533868 691718 533930 691954
rect 534166 691718 534250 691954
rect 534486 691718 534570 691954
rect 534806 691718 534868 691954
rect 533868 691634 534868 691718
rect 533868 691398 533930 691634
rect 534166 691398 534250 691634
rect 534486 691398 534570 691634
rect 534806 691398 534868 691634
rect 533868 691366 534868 691398
rect 553868 691954 554868 691986
rect 553868 691718 553930 691954
rect 554166 691718 554250 691954
rect 554486 691718 554570 691954
rect 554806 691718 554868 691954
rect 553868 691634 554868 691718
rect 553868 691398 553930 691634
rect 554166 691398 554250 691634
rect 554486 691398 554570 691634
rect 554806 691398 554868 691634
rect 553868 691366 554868 691398
rect 303868 687454 304868 687486
rect 303868 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 304868 687454
rect 303868 687134 304868 687218
rect 303868 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 304868 687134
rect 303868 686866 304868 686898
rect 323868 687454 324868 687486
rect 323868 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 324868 687454
rect 323868 687134 324868 687218
rect 323868 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 324868 687134
rect 323868 686866 324868 686898
rect 343868 687454 344868 687486
rect 343868 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 344868 687454
rect 343868 687134 344868 687218
rect 343868 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 344868 687134
rect 343868 686866 344868 686898
rect 363868 687454 364868 687486
rect 363868 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 364868 687454
rect 363868 687134 364868 687218
rect 363868 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 364868 687134
rect 363868 686866 364868 686898
rect 383868 687454 384868 687486
rect 383868 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 384868 687454
rect 383868 687134 384868 687218
rect 383868 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 384868 687134
rect 383868 686866 384868 686898
rect 403868 687454 404868 687486
rect 403868 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 404868 687454
rect 403868 687134 404868 687218
rect 403868 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 404868 687134
rect 403868 686866 404868 686898
rect 423868 687454 424868 687486
rect 423868 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 424868 687454
rect 423868 687134 424868 687218
rect 423868 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 424868 687134
rect 423868 686866 424868 686898
rect 443868 687454 444868 687486
rect 443868 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 444868 687454
rect 443868 687134 444868 687218
rect 443868 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 444868 687134
rect 443868 686866 444868 686898
rect 463868 687454 464868 687486
rect 463868 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 464868 687454
rect 463868 687134 464868 687218
rect 463868 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 464868 687134
rect 463868 686866 464868 686898
rect 483868 687454 484868 687486
rect 483868 687218 483930 687454
rect 484166 687218 484250 687454
rect 484486 687218 484570 687454
rect 484806 687218 484868 687454
rect 483868 687134 484868 687218
rect 483868 686898 483930 687134
rect 484166 686898 484250 687134
rect 484486 686898 484570 687134
rect 484806 686898 484868 687134
rect 483868 686866 484868 686898
rect 503868 687454 504868 687486
rect 503868 687218 503930 687454
rect 504166 687218 504250 687454
rect 504486 687218 504570 687454
rect 504806 687218 504868 687454
rect 503868 687134 504868 687218
rect 503868 686898 503930 687134
rect 504166 686898 504250 687134
rect 504486 686898 504570 687134
rect 504806 686898 504868 687134
rect 503868 686866 504868 686898
rect 523868 687454 524868 687486
rect 523868 687218 523930 687454
rect 524166 687218 524250 687454
rect 524486 687218 524570 687454
rect 524806 687218 524868 687454
rect 523868 687134 524868 687218
rect 523868 686898 523930 687134
rect 524166 686898 524250 687134
rect 524486 686898 524570 687134
rect 524806 686898 524868 687134
rect 523868 686866 524868 686898
rect 543868 687454 544868 687486
rect 543868 687218 543930 687454
rect 544166 687218 544250 687454
rect 544486 687218 544570 687454
rect 544806 687218 544868 687454
rect 543868 687134 544868 687218
rect 543868 686898 543930 687134
rect 544166 686898 544250 687134
rect 544486 686898 544570 687134
rect 544806 686898 544868 687134
rect 543868 686866 544868 686898
rect 563868 687454 564868 687486
rect 563868 687218 563930 687454
rect 564166 687218 564250 687454
rect 564486 687218 564570 687454
rect 564806 687218 564868 687454
rect 563868 687134 564868 687218
rect 563868 686898 563930 687134
rect 564166 686898 564250 687134
rect 564486 686898 564570 687134
rect 564806 686898 564868 687134
rect 563868 686866 564868 686898
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 313868 655954 314868 655986
rect 313868 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 314868 655954
rect 313868 655634 314868 655718
rect 313868 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 314868 655634
rect 313868 655366 314868 655398
rect 333868 655954 334868 655986
rect 333868 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 334868 655954
rect 333868 655634 334868 655718
rect 333868 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 334868 655634
rect 333868 655366 334868 655398
rect 353868 655954 354868 655986
rect 353868 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 354868 655954
rect 353868 655634 354868 655718
rect 353868 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 354868 655634
rect 353868 655366 354868 655398
rect 373868 655954 374868 655986
rect 373868 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 374868 655954
rect 373868 655634 374868 655718
rect 373868 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 374868 655634
rect 373868 655366 374868 655398
rect 393868 655954 394868 655986
rect 393868 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 394868 655954
rect 393868 655634 394868 655718
rect 393868 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 394868 655634
rect 393868 655366 394868 655398
rect 413868 655954 414868 655986
rect 413868 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 414868 655954
rect 413868 655634 414868 655718
rect 413868 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 414868 655634
rect 413868 655366 414868 655398
rect 433868 655954 434868 655986
rect 433868 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 434868 655954
rect 433868 655634 434868 655718
rect 433868 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 434868 655634
rect 433868 655366 434868 655398
rect 453868 655954 454868 655986
rect 453868 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 454868 655954
rect 453868 655634 454868 655718
rect 453868 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 454868 655634
rect 453868 655366 454868 655398
rect 473868 655954 474868 655986
rect 473868 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 474868 655954
rect 473868 655634 474868 655718
rect 473868 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 474868 655634
rect 473868 655366 474868 655398
rect 493868 655954 494868 655986
rect 493868 655718 493930 655954
rect 494166 655718 494250 655954
rect 494486 655718 494570 655954
rect 494806 655718 494868 655954
rect 493868 655634 494868 655718
rect 493868 655398 493930 655634
rect 494166 655398 494250 655634
rect 494486 655398 494570 655634
rect 494806 655398 494868 655634
rect 493868 655366 494868 655398
rect 513868 655954 514868 655986
rect 513868 655718 513930 655954
rect 514166 655718 514250 655954
rect 514486 655718 514570 655954
rect 514806 655718 514868 655954
rect 513868 655634 514868 655718
rect 513868 655398 513930 655634
rect 514166 655398 514250 655634
rect 514486 655398 514570 655634
rect 514806 655398 514868 655634
rect 513868 655366 514868 655398
rect 533868 655954 534868 655986
rect 533868 655718 533930 655954
rect 534166 655718 534250 655954
rect 534486 655718 534570 655954
rect 534806 655718 534868 655954
rect 533868 655634 534868 655718
rect 533868 655398 533930 655634
rect 534166 655398 534250 655634
rect 534486 655398 534570 655634
rect 534806 655398 534868 655634
rect 533868 655366 534868 655398
rect 553868 655954 554868 655986
rect 553868 655718 553930 655954
rect 554166 655718 554250 655954
rect 554486 655718 554570 655954
rect 554806 655718 554868 655954
rect 553868 655634 554868 655718
rect 553868 655398 553930 655634
rect 554166 655398 554250 655634
rect 554486 655398 554570 655634
rect 554806 655398 554868 655634
rect 553868 655366 554868 655398
rect 303868 651454 304868 651486
rect 303868 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 304868 651454
rect 303868 651134 304868 651218
rect 303868 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 304868 651134
rect 303868 650866 304868 650898
rect 323868 651454 324868 651486
rect 323868 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 324868 651454
rect 323868 651134 324868 651218
rect 323868 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 324868 651134
rect 323868 650866 324868 650898
rect 343868 651454 344868 651486
rect 343868 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 344868 651454
rect 343868 651134 344868 651218
rect 343868 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 344868 651134
rect 343868 650866 344868 650898
rect 363868 651454 364868 651486
rect 363868 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 364868 651454
rect 363868 651134 364868 651218
rect 363868 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 364868 651134
rect 363868 650866 364868 650898
rect 383868 651454 384868 651486
rect 383868 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 384868 651454
rect 383868 651134 384868 651218
rect 383868 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 384868 651134
rect 383868 650866 384868 650898
rect 403868 651454 404868 651486
rect 403868 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 404868 651454
rect 403868 651134 404868 651218
rect 403868 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 404868 651134
rect 403868 650866 404868 650898
rect 423868 651454 424868 651486
rect 423868 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 424868 651454
rect 423868 651134 424868 651218
rect 423868 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 424868 651134
rect 423868 650866 424868 650898
rect 443868 651454 444868 651486
rect 443868 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 444868 651454
rect 443868 651134 444868 651218
rect 443868 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 444868 651134
rect 443868 650866 444868 650898
rect 463868 651454 464868 651486
rect 463868 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 464868 651454
rect 463868 651134 464868 651218
rect 463868 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 464868 651134
rect 463868 650866 464868 650898
rect 483868 651454 484868 651486
rect 483868 651218 483930 651454
rect 484166 651218 484250 651454
rect 484486 651218 484570 651454
rect 484806 651218 484868 651454
rect 483868 651134 484868 651218
rect 483868 650898 483930 651134
rect 484166 650898 484250 651134
rect 484486 650898 484570 651134
rect 484806 650898 484868 651134
rect 483868 650866 484868 650898
rect 503868 651454 504868 651486
rect 503868 651218 503930 651454
rect 504166 651218 504250 651454
rect 504486 651218 504570 651454
rect 504806 651218 504868 651454
rect 503868 651134 504868 651218
rect 503868 650898 503930 651134
rect 504166 650898 504250 651134
rect 504486 650898 504570 651134
rect 504806 650898 504868 651134
rect 503868 650866 504868 650898
rect 523868 651454 524868 651486
rect 523868 651218 523930 651454
rect 524166 651218 524250 651454
rect 524486 651218 524570 651454
rect 524806 651218 524868 651454
rect 523868 651134 524868 651218
rect 523868 650898 523930 651134
rect 524166 650898 524250 651134
rect 524486 650898 524570 651134
rect 524806 650898 524868 651134
rect 523868 650866 524868 650898
rect 543868 651454 544868 651486
rect 543868 651218 543930 651454
rect 544166 651218 544250 651454
rect 544486 651218 544570 651454
rect 544806 651218 544868 651454
rect 543868 651134 544868 651218
rect 543868 650898 543930 651134
rect 544166 650898 544250 651134
rect 544486 650898 544570 651134
rect 544806 650898 544868 651134
rect 543868 650866 544868 650898
rect 563868 651454 564868 651486
rect 563868 651218 563930 651454
rect 564166 651218 564250 651454
rect 564486 651218 564570 651454
rect 564806 651218 564868 651454
rect 563868 651134 564868 651218
rect 563868 650898 563930 651134
rect 564166 650898 564250 651134
rect 564486 650898 564570 651134
rect 564806 650898 564868 651134
rect 563868 650866 564868 650898
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 313868 619954 314868 619986
rect 313868 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 314868 619954
rect 313868 619634 314868 619718
rect 313868 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 314868 619634
rect 313868 619366 314868 619398
rect 333868 619954 334868 619986
rect 333868 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 334868 619954
rect 333868 619634 334868 619718
rect 333868 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 334868 619634
rect 333868 619366 334868 619398
rect 353868 619954 354868 619986
rect 353868 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 354868 619954
rect 353868 619634 354868 619718
rect 353868 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 354868 619634
rect 353868 619366 354868 619398
rect 373868 619954 374868 619986
rect 373868 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 374868 619954
rect 373868 619634 374868 619718
rect 373868 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 374868 619634
rect 373868 619366 374868 619398
rect 393868 619954 394868 619986
rect 393868 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 394868 619954
rect 393868 619634 394868 619718
rect 393868 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 394868 619634
rect 393868 619366 394868 619398
rect 413868 619954 414868 619986
rect 413868 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 414868 619954
rect 413868 619634 414868 619718
rect 413868 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 414868 619634
rect 413868 619366 414868 619398
rect 433868 619954 434868 619986
rect 433868 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 434868 619954
rect 433868 619634 434868 619718
rect 433868 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 434868 619634
rect 433868 619366 434868 619398
rect 453868 619954 454868 619986
rect 453868 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 454868 619954
rect 453868 619634 454868 619718
rect 453868 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 454868 619634
rect 453868 619366 454868 619398
rect 473868 619954 474868 619986
rect 473868 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 474868 619954
rect 473868 619634 474868 619718
rect 473868 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 474868 619634
rect 473868 619366 474868 619398
rect 493868 619954 494868 619986
rect 493868 619718 493930 619954
rect 494166 619718 494250 619954
rect 494486 619718 494570 619954
rect 494806 619718 494868 619954
rect 493868 619634 494868 619718
rect 493868 619398 493930 619634
rect 494166 619398 494250 619634
rect 494486 619398 494570 619634
rect 494806 619398 494868 619634
rect 493868 619366 494868 619398
rect 513868 619954 514868 619986
rect 513868 619718 513930 619954
rect 514166 619718 514250 619954
rect 514486 619718 514570 619954
rect 514806 619718 514868 619954
rect 513868 619634 514868 619718
rect 513868 619398 513930 619634
rect 514166 619398 514250 619634
rect 514486 619398 514570 619634
rect 514806 619398 514868 619634
rect 513868 619366 514868 619398
rect 533868 619954 534868 619986
rect 533868 619718 533930 619954
rect 534166 619718 534250 619954
rect 534486 619718 534570 619954
rect 534806 619718 534868 619954
rect 533868 619634 534868 619718
rect 533868 619398 533930 619634
rect 534166 619398 534250 619634
rect 534486 619398 534570 619634
rect 534806 619398 534868 619634
rect 533868 619366 534868 619398
rect 553868 619954 554868 619986
rect 553868 619718 553930 619954
rect 554166 619718 554250 619954
rect 554486 619718 554570 619954
rect 554806 619718 554868 619954
rect 553868 619634 554868 619718
rect 553868 619398 553930 619634
rect 554166 619398 554250 619634
rect 554486 619398 554570 619634
rect 554806 619398 554868 619634
rect 553868 619366 554868 619398
rect 303868 615454 304868 615486
rect 303868 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 304868 615454
rect 303868 615134 304868 615218
rect 303868 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 304868 615134
rect 303868 614866 304868 614898
rect 323868 615454 324868 615486
rect 323868 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 324868 615454
rect 323868 615134 324868 615218
rect 323868 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 324868 615134
rect 323868 614866 324868 614898
rect 343868 615454 344868 615486
rect 343868 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 344868 615454
rect 343868 615134 344868 615218
rect 343868 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 344868 615134
rect 343868 614866 344868 614898
rect 363868 615454 364868 615486
rect 363868 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 364868 615454
rect 363868 615134 364868 615218
rect 363868 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 364868 615134
rect 363868 614866 364868 614898
rect 383868 615454 384868 615486
rect 383868 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 384868 615454
rect 383868 615134 384868 615218
rect 383868 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 384868 615134
rect 383868 614866 384868 614898
rect 403868 615454 404868 615486
rect 403868 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 404868 615454
rect 403868 615134 404868 615218
rect 403868 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 404868 615134
rect 403868 614866 404868 614898
rect 423868 615454 424868 615486
rect 423868 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 424868 615454
rect 423868 615134 424868 615218
rect 423868 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 424868 615134
rect 423868 614866 424868 614898
rect 443868 615454 444868 615486
rect 443868 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 444868 615454
rect 443868 615134 444868 615218
rect 443868 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 444868 615134
rect 443868 614866 444868 614898
rect 463868 615454 464868 615486
rect 463868 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 464868 615454
rect 463868 615134 464868 615218
rect 463868 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 464868 615134
rect 463868 614866 464868 614898
rect 483868 615454 484868 615486
rect 483868 615218 483930 615454
rect 484166 615218 484250 615454
rect 484486 615218 484570 615454
rect 484806 615218 484868 615454
rect 483868 615134 484868 615218
rect 483868 614898 483930 615134
rect 484166 614898 484250 615134
rect 484486 614898 484570 615134
rect 484806 614898 484868 615134
rect 483868 614866 484868 614898
rect 503868 615454 504868 615486
rect 503868 615218 503930 615454
rect 504166 615218 504250 615454
rect 504486 615218 504570 615454
rect 504806 615218 504868 615454
rect 503868 615134 504868 615218
rect 503868 614898 503930 615134
rect 504166 614898 504250 615134
rect 504486 614898 504570 615134
rect 504806 614898 504868 615134
rect 503868 614866 504868 614898
rect 523868 615454 524868 615486
rect 523868 615218 523930 615454
rect 524166 615218 524250 615454
rect 524486 615218 524570 615454
rect 524806 615218 524868 615454
rect 523868 615134 524868 615218
rect 523868 614898 523930 615134
rect 524166 614898 524250 615134
rect 524486 614898 524570 615134
rect 524806 614898 524868 615134
rect 523868 614866 524868 614898
rect 543868 615454 544868 615486
rect 543868 615218 543930 615454
rect 544166 615218 544250 615454
rect 544486 615218 544570 615454
rect 544806 615218 544868 615454
rect 543868 615134 544868 615218
rect 543868 614898 543930 615134
rect 544166 614898 544250 615134
rect 544486 614898 544570 615134
rect 544806 614898 544868 615134
rect 543868 614866 544868 614898
rect 563868 615454 564868 615486
rect 563868 615218 563930 615454
rect 564166 615218 564250 615454
rect 564486 615218 564570 615454
rect 564806 615218 564868 615454
rect 563868 615134 564868 615218
rect 563868 614898 563930 615134
rect 564166 614898 564250 615134
rect 564486 614898 564570 615134
rect 564806 614898 564868 615134
rect 563868 614866 564868 614898
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 571379 585716 571445 585717
rect 571379 585652 571380 585716
rect 571444 585652 571445 585716
rect 571379 585651 571445 585652
rect 566963 585172 567029 585173
rect 566963 585108 566964 585172
rect 567028 585108 567029 585172
rect 566963 585107 567029 585108
rect 565859 583132 565925 583133
rect 565859 583068 565860 583132
rect 565924 583068 565925 583132
rect 565859 583067 565925 583068
rect 313868 547954 314868 547986
rect 313868 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 314868 547954
rect 313868 547634 314868 547718
rect 313868 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 314868 547634
rect 313868 547366 314868 547398
rect 333868 547954 334868 547986
rect 333868 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 334868 547954
rect 333868 547634 334868 547718
rect 333868 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 334868 547634
rect 333868 547366 334868 547398
rect 353868 547954 354868 547986
rect 353868 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 354868 547954
rect 353868 547634 354868 547718
rect 353868 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 354868 547634
rect 353868 547366 354868 547398
rect 373868 547954 374868 547986
rect 373868 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 374868 547954
rect 373868 547634 374868 547718
rect 373868 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 374868 547634
rect 373868 547366 374868 547398
rect 393868 547954 394868 547986
rect 393868 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 394868 547954
rect 393868 547634 394868 547718
rect 393868 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 394868 547634
rect 393868 547366 394868 547398
rect 413868 547954 414868 547986
rect 413868 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 414868 547954
rect 413868 547634 414868 547718
rect 413868 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 414868 547634
rect 413868 547366 414868 547398
rect 433868 547954 434868 547986
rect 433868 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 434868 547954
rect 433868 547634 434868 547718
rect 433868 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 434868 547634
rect 433868 547366 434868 547398
rect 453868 547954 454868 547986
rect 453868 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 454868 547954
rect 453868 547634 454868 547718
rect 453868 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 454868 547634
rect 453868 547366 454868 547398
rect 473868 547954 474868 547986
rect 473868 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 474868 547954
rect 473868 547634 474868 547718
rect 473868 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 474868 547634
rect 473868 547366 474868 547398
rect 493868 547954 494868 547986
rect 493868 547718 493930 547954
rect 494166 547718 494250 547954
rect 494486 547718 494570 547954
rect 494806 547718 494868 547954
rect 493868 547634 494868 547718
rect 493868 547398 493930 547634
rect 494166 547398 494250 547634
rect 494486 547398 494570 547634
rect 494806 547398 494868 547634
rect 493868 547366 494868 547398
rect 513868 547954 514868 547986
rect 513868 547718 513930 547954
rect 514166 547718 514250 547954
rect 514486 547718 514570 547954
rect 514806 547718 514868 547954
rect 513868 547634 514868 547718
rect 513868 547398 513930 547634
rect 514166 547398 514250 547634
rect 514486 547398 514570 547634
rect 514806 547398 514868 547634
rect 513868 547366 514868 547398
rect 533868 547954 534868 547986
rect 533868 547718 533930 547954
rect 534166 547718 534250 547954
rect 534486 547718 534570 547954
rect 534806 547718 534868 547954
rect 533868 547634 534868 547718
rect 533868 547398 533930 547634
rect 534166 547398 534250 547634
rect 534486 547398 534570 547634
rect 534806 547398 534868 547634
rect 533868 547366 534868 547398
rect 553868 547954 554868 547986
rect 553868 547718 553930 547954
rect 554166 547718 554250 547954
rect 554486 547718 554570 547954
rect 554806 547718 554868 547954
rect 553868 547634 554868 547718
rect 553868 547398 553930 547634
rect 554166 547398 554250 547634
rect 554486 547398 554570 547634
rect 554806 547398 554868 547634
rect 553868 547366 554868 547398
rect 303868 543454 304868 543486
rect 303868 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 304868 543454
rect 303868 543134 304868 543218
rect 303868 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 304868 543134
rect 303868 542866 304868 542898
rect 323868 543454 324868 543486
rect 323868 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 324868 543454
rect 323868 543134 324868 543218
rect 323868 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 324868 543134
rect 323868 542866 324868 542898
rect 343868 543454 344868 543486
rect 343868 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 344868 543454
rect 343868 543134 344868 543218
rect 343868 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 344868 543134
rect 343868 542866 344868 542898
rect 363868 543454 364868 543486
rect 363868 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 364868 543454
rect 363868 543134 364868 543218
rect 363868 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 364868 543134
rect 363868 542866 364868 542898
rect 383868 543454 384868 543486
rect 383868 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 384868 543454
rect 383868 543134 384868 543218
rect 383868 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 384868 543134
rect 383868 542866 384868 542898
rect 403868 543454 404868 543486
rect 403868 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 404868 543454
rect 403868 543134 404868 543218
rect 403868 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 404868 543134
rect 403868 542866 404868 542898
rect 423868 543454 424868 543486
rect 423868 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 424868 543454
rect 423868 543134 424868 543218
rect 423868 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 424868 543134
rect 423868 542866 424868 542898
rect 443868 543454 444868 543486
rect 443868 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 444868 543454
rect 443868 543134 444868 543218
rect 443868 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 444868 543134
rect 443868 542866 444868 542898
rect 463868 543454 464868 543486
rect 463868 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 464868 543454
rect 463868 543134 464868 543218
rect 463868 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 464868 543134
rect 463868 542866 464868 542898
rect 483868 543454 484868 543486
rect 483868 543218 483930 543454
rect 484166 543218 484250 543454
rect 484486 543218 484570 543454
rect 484806 543218 484868 543454
rect 483868 543134 484868 543218
rect 483868 542898 483930 543134
rect 484166 542898 484250 543134
rect 484486 542898 484570 543134
rect 484806 542898 484868 543134
rect 483868 542866 484868 542898
rect 503868 543454 504868 543486
rect 503868 543218 503930 543454
rect 504166 543218 504250 543454
rect 504486 543218 504570 543454
rect 504806 543218 504868 543454
rect 503868 543134 504868 543218
rect 503868 542898 503930 543134
rect 504166 542898 504250 543134
rect 504486 542898 504570 543134
rect 504806 542898 504868 543134
rect 503868 542866 504868 542898
rect 523868 543454 524868 543486
rect 523868 543218 523930 543454
rect 524166 543218 524250 543454
rect 524486 543218 524570 543454
rect 524806 543218 524868 543454
rect 523868 543134 524868 543218
rect 523868 542898 523930 543134
rect 524166 542898 524250 543134
rect 524486 542898 524570 543134
rect 524806 542898 524868 543134
rect 523868 542866 524868 542898
rect 543868 543454 544868 543486
rect 543868 543218 543930 543454
rect 544166 543218 544250 543454
rect 544486 543218 544570 543454
rect 544806 543218 544868 543454
rect 543868 543134 544868 543218
rect 543868 542898 543930 543134
rect 544166 542898 544250 543134
rect 544486 542898 544570 543134
rect 544806 542898 544868 543134
rect 543868 542866 544868 542898
rect 563868 543454 564868 543486
rect 563868 543218 563930 543454
rect 564166 543218 564250 543454
rect 564486 543218 564570 543454
rect 564806 543218 564868 543454
rect 563868 543134 564868 543218
rect 563868 542898 563930 543134
rect 564166 542898 564250 543134
rect 564486 542898 564570 543134
rect 564806 542898 564868 543134
rect 563868 542866 564868 542898
rect 313868 511954 314868 511986
rect 313868 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 314868 511954
rect 313868 511634 314868 511718
rect 313868 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 314868 511634
rect 313868 511366 314868 511398
rect 333868 511954 334868 511986
rect 333868 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 334868 511954
rect 333868 511634 334868 511718
rect 333868 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 334868 511634
rect 333868 511366 334868 511398
rect 353868 511954 354868 511986
rect 353868 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 354868 511954
rect 353868 511634 354868 511718
rect 353868 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 354868 511634
rect 353868 511366 354868 511398
rect 373868 511954 374868 511986
rect 373868 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 374868 511954
rect 373868 511634 374868 511718
rect 373868 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 374868 511634
rect 373868 511366 374868 511398
rect 393868 511954 394868 511986
rect 393868 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 394868 511954
rect 393868 511634 394868 511718
rect 393868 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 394868 511634
rect 393868 511366 394868 511398
rect 413868 511954 414868 511986
rect 413868 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 414868 511954
rect 413868 511634 414868 511718
rect 413868 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 414868 511634
rect 413868 511366 414868 511398
rect 433868 511954 434868 511986
rect 433868 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 434868 511954
rect 433868 511634 434868 511718
rect 433868 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 434868 511634
rect 433868 511366 434868 511398
rect 453868 511954 454868 511986
rect 453868 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 454868 511954
rect 453868 511634 454868 511718
rect 453868 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 454868 511634
rect 453868 511366 454868 511398
rect 473868 511954 474868 511986
rect 473868 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 474868 511954
rect 473868 511634 474868 511718
rect 473868 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 474868 511634
rect 473868 511366 474868 511398
rect 493868 511954 494868 511986
rect 493868 511718 493930 511954
rect 494166 511718 494250 511954
rect 494486 511718 494570 511954
rect 494806 511718 494868 511954
rect 493868 511634 494868 511718
rect 493868 511398 493930 511634
rect 494166 511398 494250 511634
rect 494486 511398 494570 511634
rect 494806 511398 494868 511634
rect 493868 511366 494868 511398
rect 513868 511954 514868 511986
rect 513868 511718 513930 511954
rect 514166 511718 514250 511954
rect 514486 511718 514570 511954
rect 514806 511718 514868 511954
rect 513868 511634 514868 511718
rect 513868 511398 513930 511634
rect 514166 511398 514250 511634
rect 514486 511398 514570 511634
rect 514806 511398 514868 511634
rect 513868 511366 514868 511398
rect 533868 511954 534868 511986
rect 533868 511718 533930 511954
rect 534166 511718 534250 511954
rect 534486 511718 534570 511954
rect 534806 511718 534868 511954
rect 533868 511634 534868 511718
rect 533868 511398 533930 511634
rect 534166 511398 534250 511634
rect 534486 511398 534570 511634
rect 534806 511398 534868 511634
rect 533868 511366 534868 511398
rect 553868 511954 554868 511986
rect 553868 511718 553930 511954
rect 554166 511718 554250 511954
rect 554486 511718 554570 511954
rect 554806 511718 554868 511954
rect 553868 511634 554868 511718
rect 553868 511398 553930 511634
rect 554166 511398 554250 511634
rect 554486 511398 554570 511634
rect 554806 511398 554868 511634
rect 553868 511366 554868 511398
rect 303868 507454 304868 507486
rect 303868 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 304868 507454
rect 303868 507134 304868 507218
rect 303868 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 304868 507134
rect 303868 506866 304868 506898
rect 323868 507454 324868 507486
rect 323868 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 324868 507454
rect 323868 507134 324868 507218
rect 323868 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 324868 507134
rect 323868 506866 324868 506898
rect 343868 507454 344868 507486
rect 343868 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 344868 507454
rect 343868 507134 344868 507218
rect 343868 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 344868 507134
rect 343868 506866 344868 506898
rect 363868 507454 364868 507486
rect 363868 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 364868 507454
rect 363868 507134 364868 507218
rect 363868 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 364868 507134
rect 363868 506866 364868 506898
rect 383868 507454 384868 507486
rect 383868 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 384868 507454
rect 383868 507134 384868 507218
rect 383868 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 384868 507134
rect 383868 506866 384868 506898
rect 403868 507454 404868 507486
rect 403868 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 404868 507454
rect 403868 507134 404868 507218
rect 403868 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 404868 507134
rect 403868 506866 404868 506898
rect 423868 507454 424868 507486
rect 423868 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 424868 507454
rect 423868 507134 424868 507218
rect 423868 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 424868 507134
rect 423868 506866 424868 506898
rect 443868 507454 444868 507486
rect 443868 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 444868 507454
rect 443868 507134 444868 507218
rect 443868 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 444868 507134
rect 443868 506866 444868 506898
rect 463868 507454 464868 507486
rect 463868 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 464868 507454
rect 463868 507134 464868 507218
rect 463868 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 464868 507134
rect 463868 506866 464868 506898
rect 483868 507454 484868 507486
rect 483868 507218 483930 507454
rect 484166 507218 484250 507454
rect 484486 507218 484570 507454
rect 484806 507218 484868 507454
rect 483868 507134 484868 507218
rect 483868 506898 483930 507134
rect 484166 506898 484250 507134
rect 484486 506898 484570 507134
rect 484806 506898 484868 507134
rect 483868 506866 484868 506898
rect 503868 507454 504868 507486
rect 503868 507218 503930 507454
rect 504166 507218 504250 507454
rect 504486 507218 504570 507454
rect 504806 507218 504868 507454
rect 503868 507134 504868 507218
rect 503868 506898 503930 507134
rect 504166 506898 504250 507134
rect 504486 506898 504570 507134
rect 504806 506898 504868 507134
rect 503868 506866 504868 506898
rect 523868 507454 524868 507486
rect 523868 507218 523930 507454
rect 524166 507218 524250 507454
rect 524486 507218 524570 507454
rect 524806 507218 524868 507454
rect 523868 507134 524868 507218
rect 523868 506898 523930 507134
rect 524166 506898 524250 507134
rect 524486 506898 524570 507134
rect 524806 506898 524868 507134
rect 523868 506866 524868 506898
rect 543868 507454 544868 507486
rect 543868 507218 543930 507454
rect 544166 507218 544250 507454
rect 544486 507218 544570 507454
rect 544806 507218 544868 507454
rect 543868 507134 544868 507218
rect 543868 506898 543930 507134
rect 544166 506898 544250 507134
rect 544486 506898 544570 507134
rect 544806 506898 544868 507134
rect 543868 506866 544868 506898
rect 563868 507454 564868 507486
rect 563868 507218 563930 507454
rect 564166 507218 564250 507454
rect 564486 507218 564570 507454
rect 564806 507218 564868 507454
rect 563868 507134 564868 507218
rect 563868 506898 563930 507134
rect 564166 506898 564250 507134
rect 564486 506898 564570 507134
rect 564806 506898 564868 507134
rect 563868 506866 564868 506898
rect 313868 475954 314868 475986
rect 313868 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 314868 475954
rect 313868 475634 314868 475718
rect 313868 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 314868 475634
rect 313868 475366 314868 475398
rect 333868 475954 334868 475986
rect 333868 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 334868 475954
rect 333868 475634 334868 475718
rect 333868 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 334868 475634
rect 333868 475366 334868 475398
rect 353868 475954 354868 475986
rect 353868 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 354868 475954
rect 353868 475634 354868 475718
rect 353868 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 354868 475634
rect 353868 475366 354868 475398
rect 373868 475954 374868 475986
rect 373868 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 374868 475954
rect 373868 475634 374868 475718
rect 373868 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 374868 475634
rect 373868 475366 374868 475398
rect 393868 475954 394868 475986
rect 393868 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 394868 475954
rect 393868 475634 394868 475718
rect 393868 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 394868 475634
rect 393868 475366 394868 475398
rect 413868 475954 414868 475986
rect 413868 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 414868 475954
rect 413868 475634 414868 475718
rect 413868 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 414868 475634
rect 413868 475366 414868 475398
rect 433868 475954 434868 475986
rect 433868 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 434868 475954
rect 433868 475634 434868 475718
rect 433868 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 434868 475634
rect 433868 475366 434868 475398
rect 453868 475954 454868 475986
rect 453868 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 454868 475954
rect 453868 475634 454868 475718
rect 453868 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 454868 475634
rect 453868 475366 454868 475398
rect 473868 475954 474868 475986
rect 473868 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 474868 475954
rect 473868 475634 474868 475718
rect 473868 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 474868 475634
rect 473868 475366 474868 475398
rect 493868 475954 494868 475986
rect 493868 475718 493930 475954
rect 494166 475718 494250 475954
rect 494486 475718 494570 475954
rect 494806 475718 494868 475954
rect 493868 475634 494868 475718
rect 493868 475398 493930 475634
rect 494166 475398 494250 475634
rect 494486 475398 494570 475634
rect 494806 475398 494868 475634
rect 493868 475366 494868 475398
rect 513868 475954 514868 475986
rect 513868 475718 513930 475954
rect 514166 475718 514250 475954
rect 514486 475718 514570 475954
rect 514806 475718 514868 475954
rect 513868 475634 514868 475718
rect 513868 475398 513930 475634
rect 514166 475398 514250 475634
rect 514486 475398 514570 475634
rect 514806 475398 514868 475634
rect 513868 475366 514868 475398
rect 533868 475954 534868 475986
rect 533868 475718 533930 475954
rect 534166 475718 534250 475954
rect 534486 475718 534570 475954
rect 534806 475718 534868 475954
rect 533868 475634 534868 475718
rect 533868 475398 533930 475634
rect 534166 475398 534250 475634
rect 534486 475398 534570 475634
rect 534806 475398 534868 475634
rect 533868 475366 534868 475398
rect 553868 475954 554868 475986
rect 553868 475718 553930 475954
rect 554166 475718 554250 475954
rect 554486 475718 554570 475954
rect 554806 475718 554868 475954
rect 553868 475634 554868 475718
rect 553868 475398 553930 475634
rect 554166 475398 554250 475634
rect 554486 475398 554570 475634
rect 554806 475398 554868 475634
rect 553868 475366 554868 475398
rect 303868 471454 304868 471486
rect 303868 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 304868 471454
rect 303868 471134 304868 471218
rect 303868 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 304868 471134
rect 303868 470866 304868 470898
rect 323868 471454 324868 471486
rect 323868 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 324868 471454
rect 323868 471134 324868 471218
rect 323868 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 324868 471134
rect 323868 470866 324868 470898
rect 343868 471454 344868 471486
rect 343868 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 344868 471454
rect 343868 471134 344868 471218
rect 343868 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 344868 471134
rect 343868 470866 344868 470898
rect 363868 471454 364868 471486
rect 363868 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 364868 471454
rect 363868 471134 364868 471218
rect 363868 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 364868 471134
rect 363868 470866 364868 470898
rect 383868 471454 384868 471486
rect 383868 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 384868 471454
rect 383868 471134 384868 471218
rect 383868 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 384868 471134
rect 383868 470866 384868 470898
rect 403868 471454 404868 471486
rect 403868 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 404868 471454
rect 403868 471134 404868 471218
rect 403868 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 404868 471134
rect 403868 470866 404868 470898
rect 423868 471454 424868 471486
rect 423868 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 424868 471454
rect 423868 471134 424868 471218
rect 423868 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 424868 471134
rect 423868 470866 424868 470898
rect 443868 471454 444868 471486
rect 443868 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 444868 471454
rect 443868 471134 444868 471218
rect 443868 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 444868 471134
rect 443868 470866 444868 470898
rect 463868 471454 464868 471486
rect 463868 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 464868 471454
rect 463868 471134 464868 471218
rect 463868 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 464868 471134
rect 463868 470866 464868 470898
rect 483868 471454 484868 471486
rect 483868 471218 483930 471454
rect 484166 471218 484250 471454
rect 484486 471218 484570 471454
rect 484806 471218 484868 471454
rect 483868 471134 484868 471218
rect 483868 470898 483930 471134
rect 484166 470898 484250 471134
rect 484486 470898 484570 471134
rect 484806 470898 484868 471134
rect 483868 470866 484868 470898
rect 503868 471454 504868 471486
rect 503868 471218 503930 471454
rect 504166 471218 504250 471454
rect 504486 471218 504570 471454
rect 504806 471218 504868 471454
rect 503868 471134 504868 471218
rect 503868 470898 503930 471134
rect 504166 470898 504250 471134
rect 504486 470898 504570 471134
rect 504806 470898 504868 471134
rect 503868 470866 504868 470898
rect 523868 471454 524868 471486
rect 523868 471218 523930 471454
rect 524166 471218 524250 471454
rect 524486 471218 524570 471454
rect 524806 471218 524868 471454
rect 523868 471134 524868 471218
rect 523868 470898 523930 471134
rect 524166 470898 524250 471134
rect 524486 470898 524570 471134
rect 524806 470898 524868 471134
rect 523868 470866 524868 470898
rect 543868 471454 544868 471486
rect 543868 471218 543930 471454
rect 544166 471218 544250 471454
rect 544486 471218 544570 471454
rect 544806 471218 544868 471454
rect 543868 471134 544868 471218
rect 543868 470898 543930 471134
rect 544166 470898 544250 471134
rect 544486 470898 544570 471134
rect 544806 470898 544868 471134
rect 543868 470866 544868 470898
rect 563868 471454 564868 471486
rect 563868 471218 563930 471454
rect 564166 471218 564250 471454
rect 564486 471218 564570 471454
rect 564806 471218 564868 471454
rect 563868 471134 564868 471218
rect 563868 470898 563930 471134
rect 564166 470898 564250 471134
rect 564486 470898 564570 471134
rect 564806 470898 564868 471134
rect 563868 470866 564868 470898
rect 303475 461956 303541 461957
rect 303475 461892 303476 461956
rect 303540 461892 303541 461956
rect 303475 461891 303541 461892
rect 302003 461820 302069 461821
rect 302003 461756 302004 461820
rect 302068 461756 302069 461820
rect 302003 461755 302069 461756
rect 301635 459508 301701 459509
rect 301635 459444 301636 459508
rect 301700 459444 301701 459508
rect 301635 459443 301701 459444
rect 299979 458964 300045 458965
rect 299979 458900 299980 458964
rect 300044 458900 300045 458964
rect 299979 458899 300045 458900
rect 301451 458964 301517 458965
rect 301451 458900 301452 458964
rect 301516 458900 301517 458964
rect 301451 458899 301517 458900
rect 298691 443732 298757 443733
rect 298691 443668 298692 443732
rect 298756 443668 298757 443732
rect 298691 443667 298757 443668
rect 298694 442917 298754 443667
rect 298691 442916 298757 442917
rect 298691 442852 298692 442916
rect 298756 442852 298757 442916
rect 298691 442851 298757 442852
rect 298694 330581 298754 442851
rect 298691 330580 298757 330581
rect 298691 330516 298692 330580
rect 298756 330516 298757 330580
rect 298691 330515 298757 330516
rect 298691 329764 298757 329765
rect 298691 329700 298692 329764
rect 298756 329700 298757 329764
rect 298691 329699 298757 329700
rect 298694 201245 298754 329699
rect 299243 307732 299309 307733
rect 299243 307668 299244 307732
rect 299308 307668 299309 307732
rect 299243 307667 299309 307668
rect 299246 206005 299306 307667
rect 299243 206004 299309 206005
rect 299243 205940 299244 206004
rect 299308 205940 299309 206004
rect 299243 205939 299309 205940
rect 298691 201244 298757 201245
rect 298691 201180 298692 201244
rect 298756 201180 298757 201244
rect 298691 201179 298757 201180
rect 298875 200700 298941 200701
rect 298875 200636 298876 200700
rect 298940 200636 298941 200700
rect 298875 200635 298941 200636
rect 298691 185876 298757 185877
rect 298691 185812 298692 185876
rect 298756 185812 298757 185876
rect 298691 185811 298757 185812
rect 297955 76940 298021 76941
rect 297955 76876 297956 76940
rect 298020 76876 298021 76940
rect 297955 76875 298021 76876
rect 298694 68237 298754 185811
rect 298878 73949 298938 200635
rect 298875 73948 298941 73949
rect 298875 73884 298876 73948
rect 298940 73884 298941 73948
rect 298875 73883 298941 73884
rect 298691 68236 298757 68237
rect 298691 68172 298692 68236
rect 298756 68172 298757 68236
rect 298691 68171 298757 68172
rect 297771 57356 297837 57357
rect 297771 57292 297772 57356
rect 297836 57292 297837 57356
rect 297771 57291 297837 57292
rect 299982 54637 300042 458899
rect 300163 315484 300229 315485
rect 300163 315420 300164 315484
rect 300228 315420 300229 315484
rect 300163 315419 300229 315420
rect 299979 54636 300045 54637
rect 299979 54572 299980 54636
rect 300044 54572 300045 54636
rect 299979 54571 300045 54572
rect 300166 54501 300226 315419
rect 301454 204917 301514 458899
rect 301638 458285 301698 459443
rect 302739 459100 302805 459101
rect 302739 459036 302740 459100
rect 302804 459036 302805 459100
rect 302739 459035 302805 459036
rect 565675 459100 565741 459101
rect 565675 459036 565676 459100
rect 565740 459036 565741 459100
rect 565675 459035 565741 459036
rect 301635 458284 301701 458285
rect 301635 458220 301636 458284
rect 301700 458220 301701 458284
rect 301635 458219 301701 458220
rect 302003 442916 302069 442917
rect 302003 442852 302004 442916
rect 302068 442852 302069 442916
rect 302003 442851 302069 442852
rect 302006 334117 302066 442851
rect 302003 334116 302069 334117
rect 302003 334052 302004 334116
rect 302068 334052 302069 334116
rect 302003 334051 302069 334052
rect 301635 331940 301701 331941
rect 301635 331876 301636 331940
rect 301700 331876 301701 331940
rect 301635 331875 301701 331876
rect 301638 205733 301698 331875
rect 301635 205732 301701 205733
rect 301635 205668 301636 205732
rect 301700 205668 301701 205732
rect 301635 205667 301701 205668
rect 301451 204916 301517 204917
rect 301451 204852 301452 204916
rect 301516 204852 301517 204916
rect 301451 204851 301517 204852
rect 301635 203556 301701 203557
rect 301635 203492 301636 203556
rect 301700 203492 301701 203556
rect 301635 203491 301701 203492
rect 301638 76669 301698 203491
rect 302003 187644 302069 187645
rect 302003 187580 302004 187644
rect 302068 187580 302069 187644
rect 302003 187579 302069 187580
rect 302006 77757 302066 187579
rect 302003 77756 302069 77757
rect 302003 77692 302004 77756
rect 302068 77692 302069 77756
rect 302003 77691 302069 77692
rect 302742 76805 302802 459035
rect 313868 439954 314868 439986
rect 313868 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 314868 439954
rect 313868 439634 314868 439718
rect 313868 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 314868 439634
rect 313868 439366 314868 439398
rect 333868 439954 334868 439986
rect 333868 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 334868 439954
rect 333868 439634 334868 439718
rect 333868 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 334868 439634
rect 333868 439366 334868 439398
rect 353868 439954 354868 439986
rect 353868 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 354868 439954
rect 353868 439634 354868 439718
rect 353868 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 354868 439634
rect 353868 439366 354868 439398
rect 373868 439954 374868 439986
rect 373868 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 374868 439954
rect 373868 439634 374868 439718
rect 373868 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 374868 439634
rect 373868 439366 374868 439398
rect 393868 439954 394868 439986
rect 393868 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 394868 439954
rect 393868 439634 394868 439718
rect 393868 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 394868 439634
rect 393868 439366 394868 439398
rect 413868 439954 414868 439986
rect 413868 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 414868 439954
rect 413868 439634 414868 439718
rect 413868 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 414868 439634
rect 413868 439366 414868 439398
rect 433868 439954 434868 439986
rect 433868 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 434868 439954
rect 433868 439634 434868 439718
rect 433868 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 434868 439634
rect 433868 439366 434868 439398
rect 453868 439954 454868 439986
rect 453868 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 454868 439954
rect 453868 439634 454868 439718
rect 453868 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 454868 439634
rect 453868 439366 454868 439398
rect 473868 439954 474868 439986
rect 473868 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 474868 439954
rect 473868 439634 474868 439718
rect 473868 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 474868 439634
rect 473868 439366 474868 439398
rect 493868 439954 494868 439986
rect 493868 439718 493930 439954
rect 494166 439718 494250 439954
rect 494486 439718 494570 439954
rect 494806 439718 494868 439954
rect 493868 439634 494868 439718
rect 493868 439398 493930 439634
rect 494166 439398 494250 439634
rect 494486 439398 494570 439634
rect 494806 439398 494868 439634
rect 493868 439366 494868 439398
rect 513868 439954 514868 439986
rect 513868 439718 513930 439954
rect 514166 439718 514250 439954
rect 514486 439718 514570 439954
rect 514806 439718 514868 439954
rect 513868 439634 514868 439718
rect 513868 439398 513930 439634
rect 514166 439398 514250 439634
rect 514486 439398 514570 439634
rect 514806 439398 514868 439634
rect 513868 439366 514868 439398
rect 533868 439954 534868 439986
rect 533868 439718 533930 439954
rect 534166 439718 534250 439954
rect 534486 439718 534570 439954
rect 534806 439718 534868 439954
rect 533868 439634 534868 439718
rect 533868 439398 533930 439634
rect 534166 439398 534250 439634
rect 534486 439398 534570 439634
rect 534806 439398 534868 439634
rect 533868 439366 534868 439398
rect 553868 439954 554868 439986
rect 553868 439718 553930 439954
rect 554166 439718 554250 439954
rect 554486 439718 554570 439954
rect 554806 439718 554868 439954
rect 553868 439634 554868 439718
rect 553868 439398 553930 439634
rect 554166 439398 554250 439634
rect 554486 439398 554570 439634
rect 554806 439398 554868 439634
rect 553868 439366 554868 439398
rect 303868 435454 304868 435486
rect 303868 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 304868 435454
rect 303868 435134 304868 435218
rect 303868 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 304868 435134
rect 303868 434866 304868 434898
rect 323868 435454 324868 435486
rect 323868 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 324868 435454
rect 323868 435134 324868 435218
rect 323868 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 324868 435134
rect 323868 434866 324868 434898
rect 343868 435454 344868 435486
rect 343868 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 344868 435454
rect 343868 435134 344868 435218
rect 343868 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 344868 435134
rect 343868 434866 344868 434898
rect 363868 435454 364868 435486
rect 363868 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 364868 435454
rect 363868 435134 364868 435218
rect 363868 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 364868 435134
rect 363868 434866 364868 434898
rect 383868 435454 384868 435486
rect 383868 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 384868 435454
rect 383868 435134 384868 435218
rect 383868 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 384868 435134
rect 383868 434866 384868 434898
rect 403868 435454 404868 435486
rect 403868 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 404868 435454
rect 403868 435134 404868 435218
rect 403868 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 404868 435134
rect 403868 434866 404868 434898
rect 423868 435454 424868 435486
rect 423868 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 424868 435454
rect 423868 435134 424868 435218
rect 423868 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 424868 435134
rect 423868 434866 424868 434898
rect 443868 435454 444868 435486
rect 443868 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 444868 435454
rect 443868 435134 444868 435218
rect 443868 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 444868 435134
rect 443868 434866 444868 434898
rect 463868 435454 464868 435486
rect 463868 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 464868 435454
rect 463868 435134 464868 435218
rect 463868 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 464868 435134
rect 463868 434866 464868 434898
rect 483868 435454 484868 435486
rect 483868 435218 483930 435454
rect 484166 435218 484250 435454
rect 484486 435218 484570 435454
rect 484806 435218 484868 435454
rect 483868 435134 484868 435218
rect 483868 434898 483930 435134
rect 484166 434898 484250 435134
rect 484486 434898 484570 435134
rect 484806 434898 484868 435134
rect 483868 434866 484868 434898
rect 503868 435454 504868 435486
rect 503868 435218 503930 435454
rect 504166 435218 504250 435454
rect 504486 435218 504570 435454
rect 504806 435218 504868 435454
rect 503868 435134 504868 435218
rect 503868 434898 503930 435134
rect 504166 434898 504250 435134
rect 504486 434898 504570 435134
rect 504806 434898 504868 435134
rect 503868 434866 504868 434898
rect 523868 435454 524868 435486
rect 523868 435218 523930 435454
rect 524166 435218 524250 435454
rect 524486 435218 524570 435454
rect 524806 435218 524868 435454
rect 523868 435134 524868 435218
rect 523868 434898 523930 435134
rect 524166 434898 524250 435134
rect 524486 434898 524570 435134
rect 524806 434898 524868 435134
rect 523868 434866 524868 434898
rect 543868 435454 544868 435486
rect 543868 435218 543930 435454
rect 544166 435218 544250 435454
rect 544486 435218 544570 435454
rect 544806 435218 544868 435454
rect 543868 435134 544868 435218
rect 543868 434898 543930 435134
rect 544166 434898 544250 435134
rect 544486 434898 544570 435134
rect 544806 434898 544868 435134
rect 543868 434866 544868 434898
rect 563868 435454 564868 435486
rect 563868 435218 563930 435454
rect 564166 435218 564250 435454
rect 564486 435218 564570 435454
rect 564806 435218 564868 435454
rect 563868 435134 564868 435218
rect 563868 434898 563930 435134
rect 564166 434898 564250 435134
rect 564486 434898 564570 435134
rect 564806 434898 564868 435134
rect 563868 434866 564868 434898
rect 565678 433397 565738 459035
rect 565862 458149 565922 583067
rect 566043 582996 566109 582997
rect 566043 582932 566044 582996
rect 566108 582932 566109 582996
rect 566043 582931 566109 582932
rect 565859 458148 565925 458149
rect 565859 458084 565860 458148
rect 565924 458084 565925 458148
rect 565859 458083 565925 458084
rect 565862 451290 565922 458083
rect 566046 457469 566106 582931
rect 566043 457468 566109 457469
rect 566043 457404 566044 457468
rect 566108 457404 566109 457468
rect 566043 457403 566109 457404
rect 565862 451230 566474 451290
rect 565675 433396 565741 433397
rect 565675 433332 565676 433396
rect 565740 433332 565741 433396
rect 565675 433331 565741 433332
rect 313868 403954 314868 403986
rect 313868 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 314868 403954
rect 313868 403634 314868 403718
rect 313868 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 314868 403634
rect 313868 403366 314868 403398
rect 333868 403954 334868 403986
rect 333868 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 334868 403954
rect 333868 403634 334868 403718
rect 333868 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 334868 403634
rect 333868 403366 334868 403398
rect 353868 403954 354868 403986
rect 353868 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 354868 403954
rect 353868 403634 354868 403718
rect 353868 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 354868 403634
rect 353868 403366 354868 403398
rect 373868 403954 374868 403986
rect 373868 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 374868 403954
rect 373868 403634 374868 403718
rect 373868 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 374868 403634
rect 373868 403366 374868 403398
rect 393868 403954 394868 403986
rect 393868 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 394868 403954
rect 393868 403634 394868 403718
rect 393868 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 394868 403634
rect 393868 403366 394868 403398
rect 413868 403954 414868 403986
rect 413868 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 414868 403954
rect 413868 403634 414868 403718
rect 413868 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 414868 403634
rect 413868 403366 414868 403398
rect 433868 403954 434868 403986
rect 433868 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 434868 403954
rect 433868 403634 434868 403718
rect 433868 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 434868 403634
rect 433868 403366 434868 403398
rect 453868 403954 454868 403986
rect 453868 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 454868 403954
rect 453868 403634 454868 403718
rect 453868 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 454868 403634
rect 453868 403366 454868 403398
rect 473868 403954 474868 403986
rect 473868 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 474868 403954
rect 473868 403634 474868 403718
rect 473868 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 474868 403634
rect 473868 403366 474868 403398
rect 493868 403954 494868 403986
rect 493868 403718 493930 403954
rect 494166 403718 494250 403954
rect 494486 403718 494570 403954
rect 494806 403718 494868 403954
rect 493868 403634 494868 403718
rect 493868 403398 493930 403634
rect 494166 403398 494250 403634
rect 494486 403398 494570 403634
rect 494806 403398 494868 403634
rect 493868 403366 494868 403398
rect 513868 403954 514868 403986
rect 513868 403718 513930 403954
rect 514166 403718 514250 403954
rect 514486 403718 514570 403954
rect 514806 403718 514868 403954
rect 513868 403634 514868 403718
rect 513868 403398 513930 403634
rect 514166 403398 514250 403634
rect 514486 403398 514570 403634
rect 514806 403398 514868 403634
rect 513868 403366 514868 403398
rect 533868 403954 534868 403986
rect 533868 403718 533930 403954
rect 534166 403718 534250 403954
rect 534486 403718 534570 403954
rect 534806 403718 534868 403954
rect 533868 403634 534868 403718
rect 533868 403398 533930 403634
rect 534166 403398 534250 403634
rect 534486 403398 534570 403634
rect 534806 403398 534868 403634
rect 533868 403366 534868 403398
rect 553868 403954 554868 403986
rect 553868 403718 553930 403954
rect 554166 403718 554250 403954
rect 554486 403718 554570 403954
rect 554806 403718 554868 403954
rect 553868 403634 554868 403718
rect 553868 403398 553930 403634
rect 554166 403398 554250 403634
rect 554486 403398 554570 403634
rect 554806 403398 554868 403634
rect 553868 403366 554868 403398
rect 303868 399454 304868 399486
rect 303868 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 304868 399454
rect 303868 399134 304868 399218
rect 303868 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 304868 399134
rect 303868 398866 304868 398898
rect 323868 399454 324868 399486
rect 323868 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 324868 399454
rect 323868 399134 324868 399218
rect 323868 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 324868 399134
rect 323868 398866 324868 398898
rect 343868 399454 344868 399486
rect 343868 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 344868 399454
rect 343868 399134 344868 399218
rect 343868 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 344868 399134
rect 343868 398866 344868 398898
rect 363868 399454 364868 399486
rect 363868 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 364868 399454
rect 363868 399134 364868 399218
rect 363868 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 364868 399134
rect 363868 398866 364868 398898
rect 383868 399454 384868 399486
rect 383868 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 384868 399454
rect 383868 399134 384868 399218
rect 383868 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 384868 399134
rect 383868 398866 384868 398898
rect 403868 399454 404868 399486
rect 403868 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 404868 399454
rect 403868 399134 404868 399218
rect 403868 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 404868 399134
rect 403868 398866 404868 398898
rect 423868 399454 424868 399486
rect 423868 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 424868 399454
rect 423868 399134 424868 399218
rect 423868 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 424868 399134
rect 423868 398866 424868 398898
rect 443868 399454 444868 399486
rect 443868 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 444868 399454
rect 443868 399134 444868 399218
rect 443868 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 444868 399134
rect 443868 398866 444868 398898
rect 463868 399454 464868 399486
rect 463868 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 464868 399454
rect 463868 399134 464868 399218
rect 463868 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 464868 399134
rect 463868 398866 464868 398898
rect 483868 399454 484868 399486
rect 483868 399218 483930 399454
rect 484166 399218 484250 399454
rect 484486 399218 484570 399454
rect 484806 399218 484868 399454
rect 483868 399134 484868 399218
rect 483868 398898 483930 399134
rect 484166 398898 484250 399134
rect 484486 398898 484570 399134
rect 484806 398898 484868 399134
rect 483868 398866 484868 398898
rect 503868 399454 504868 399486
rect 503868 399218 503930 399454
rect 504166 399218 504250 399454
rect 504486 399218 504570 399454
rect 504806 399218 504868 399454
rect 503868 399134 504868 399218
rect 503868 398898 503930 399134
rect 504166 398898 504250 399134
rect 504486 398898 504570 399134
rect 504806 398898 504868 399134
rect 503868 398866 504868 398898
rect 523868 399454 524868 399486
rect 523868 399218 523930 399454
rect 524166 399218 524250 399454
rect 524486 399218 524570 399454
rect 524806 399218 524868 399454
rect 523868 399134 524868 399218
rect 523868 398898 523930 399134
rect 524166 398898 524250 399134
rect 524486 398898 524570 399134
rect 524806 398898 524868 399134
rect 523868 398866 524868 398898
rect 543868 399454 544868 399486
rect 543868 399218 543930 399454
rect 544166 399218 544250 399454
rect 544486 399218 544570 399454
rect 544806 399218 544868 399454
rect 543868 399134 544868 399218
rect 543868 398898 543930 399134
rect 544166 398898 544250 399134
rect 544486 398898 544570 399134
rect 544806 398898 544868 399134
rect 543868 398866 544868 398898
rect 563868 399454 564868 399486
rect 563868 399218 563930 399454
rect 564166 399218 564250 399454
rect 564486 399218 564570 399454
rect 564806 399218 564868 399454
rect 563868 399134 564868 399218
rect 563868 398898 563930 399134
rect 564166 398898 564250 399134
rect 564486 398898 564570 399134
rect 564806 398898 564868 399134
rect 563868 398866 564868 398898
rect 313868 367954 314868 367986
rect 313868 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 314868 367954
rect 313868 367634 314868 367718
rect 313868 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 314868 367634
rect 313868 367366 314868 367398
rect 333868 367954 334868 367986
rect 333868 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 334868 367954
rect 333868 367634 334868 367718
rect 333868 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 334868 367634
rect 333868 367366 334868 367398
rect 353868 367954 354868 367986
rect 353868 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 354868 367954
rect 353868 367634 354868 367718
rect 353868 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 354868 367634
rect 353868 367366 354868 367398
rect 373868 367954 374868 367986
rect 373868 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 374868 367954
rect 373868 367634 374868 367718
rect 373868 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 374868 367634
rect 373868 367366 374868 367398
rect 393868 367954 394868 367986
rect 393868 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 394868 367954
rect 393868 367634 394868 367718
rect 393868 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 394868 367634
rect 393868 367366 394868 367398
rect 413868 367954 414868 367986
rect 413868 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 414868 367954
rect 413868 367634 414868 367718
rect 413868 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 414868 367634
rect 413868 367366 414868 367398
rect 433868 367954 434868 367986
rect 433868 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 434868 367954
rect 433868 367634 434868 367718
rect 433868 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 434868 367634
rect 433868 367366 434868 367398
rect 453868 367954 454868 367986
rect 453868 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 454868 367954
rect 453868 367634 454868 367718
rect 453868 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 454868 367634
rect 453868 367366 454868 367398
rect 473868 367954 474868 367986
rect 473868 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 474868 367954
rect 473868 367634 474868 367718
rect 473868 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 474868 367634
rect 473868 367366 474868 367398
rect 493868 367954 494868 367986
rect 493868 367718 493930 367954
rect 494166 367718 494250 367954
rect 494486 367718 494570 367954
rect 494806 367718 494868 367954
rect 493868 367634 494868 367718
rect 493868 367398 493930 367634
rect 494166 367398 494250 367634
rect 494486 367398 494570 367634
rect 494806 367398 494868 367634
rect 493868 367366 494868 367398
rect 513868 367954 514868 367986
rect 513868 367718 513930 367954
rect 514166 367718 514250 367954
rect 514486 367718 514570 367954
rect 514806 367718 514868 367954
rect 513868 367634 514868 367718
rect 513868 367398 513930 367634
rect 514166 367398 514250 367634
rect 514486 367398 514570 367634
rect 514806 367398 514868 367634
rect 513868 367366 514868 367398
rect 533868 367954 534868 367986
rect 533868 367718 533930 367954
rect 534166 367718 534250 367954
rect 534486 367718 534570 367954
rect 534806 367718 534868 367954
rect 533868 367634 534868 367718
rect 533868 367398 533930 367634
rect 534166 367398 534250 367634
rect 534486 367398 534570 367634
rect 534806 367398 534868 367634
rect 533868 367366 534868 367398
rect 553868 367954 554868 367986
rect 553868 367718 553930 367954
rect 554166 367718 554250 367954
rect 554486 367718 554570 367954
rect 554806 367718 554868 367954
rect 553868 367634 554868 367718
rect 553868 367398 553930 367634
rect 554166 367398 554250 367634
rect 554486 367398 554570 367634
rect 554806 367398 554868 367634
rect 553868 367366 554868 367398
rect 303868 363454 304868 363486
rect 303868 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 304868 363454
rect 303868 363134 304868 363218
rect 303868 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 304868 363134
rect 303868 362866 304868 362898
rect 323868 363454 324868 363486
rect 323868 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 324868 363454
rect 323868 363134 324868 363218
rect 323868 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 324868 363134
rect 323868 362866 324868 362898
rect 343868 363454 344868 363486
rect 343868 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 344868 363454
rect 343868 363134 344868 363218
rect 343868 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 344868 363134
rect 343868 362866 344868 362898
rect 363868 363454 364868 363486
rect 363868 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 364868 363454
rect 363868 363134 364868 363218
rect 363868 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 364868 363134
rect 363868 362866 364868 362898
rect 383868 363454 384868 363486
rect 383868 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 384868 363454
rect 383868 363134 384868 363218
rect 383868 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 384868 363134
rect 383868 362866 384868 362898
rect 403868 363454 404868 363486
rect 403868 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 404868 363454
rect 403868 363134 404868 363218
rect 403868 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 404868 363134
rect 403868 362866 404868 362898
rect 423868 363454 424868 363486
rect 423868 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 424868 363454
rect 423868 363134 424868 363218
rect 423868 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 424868 363134
rect 423868 362866 424868 362898
rect 443868 363454 444868 363486
rect 443868 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 444868 363454
rect 443868 363134 444868 363218
rect 443868 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 444868 363134
rect 443868 362866 444868 362898
rect 463868 363454 464868 363486
rect 463868 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 464868 363454
rect 463868 363134 464868 363218
rect 463868 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 464868 363134
rect 463868 362866 464868 362898
rect 483868 363454 484868 363486
rect 483868 363218 483930 363454
rect 484166 363218 484250 363454
rect 484486 363218 484570 363454
rect 484806 363218 484868 363454
rect 483868 363134 484868 363218
rect 483868 362898 483930 363134
rect 484166 362898 484250 363134
rect 484486 362898 484570 363134
rect 484806 362898 484868 363134
rect 483868 362866 484868 362898
rect 503868 363454 504868 363486
rect 503868 363218 503930 363454
rect 504166 363218 504250 363454
rect 504486 363218 504570 363454
rect 504806 363218 504868 363454
rect 503868 363134 504868 363218
rect 503868 362898 503930 363134
rect 504166 362898 504250 363134
rect 504486 362898 504570 363134
rect 504806 362898 504868 363134
rect 503868 362866 504868 362898
rect 523868 363454 524868 363486
rect 523868 363218 523930 363454
rect 524166 363218 524250 363454
rect 524486 363218 524570 363454
rect 524806 363218 524868 363454
rect 523868 363134 524868 363218
rect 523868 362898 523930 363134
rect 524166 362898 524250 363134
rect 524486 362898 524570 363134
rect 524806 362898 524868 363134
rect 523868 362866 524868 362898
rect 543868 363454 544868 363486
rect 543868 363218 543930 363454
rect 544166 363218 544250 363454
rect 544486 363218 544570 363454
rect 544806 363218 544868 363454
rect 543868 363134 544868 363218
rect 543868 362898 543930 363134
rect 544166 362898 544250 363134
rect 544486 362898 544570 363134
rect 544806 362898 544868 363134
rect 543868 362866 544868 362898
rect 563868 363454 564868 363486
rect 563868 363218 563930 363454
rect 564166 363218 564250 363454
rect 564486 363218 564570 363454
rect 564806 363218 564868 363454
rect 563868 363134 564868 363218
rect 563868 362898 563930 363134
rect 564166 362898 564250 363134
rect 564486 362898 564570 363134
rect 564806 362898 564868 363134
rect 563868 362866 564868 362898
rect 565859 331396 565925 331397
rect 565859 331332 565860 331396
rect 565924 331332 565925 331396
rect 565859 331331 565925 331332
rect 303475 318068 303541 318069
rect 303475 318004 303476 318068
rect 303540 318004 303541 318068
rect 303475 318003 303541 318004
rect 303478 205597 303538 318003
rect 313868 295954 314868 295986
rect 313868 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 314868 295954
rect 313868 295634 314868 295718
rect 313868 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 314868 295634
rect 313868 295366 314868 295398
rect 333868 295954 334868 295986
rect 333868 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 334868 295954
rect 333868 295634 334868 295718
rect 333868 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 334868 295634
rect 333868 295366 334868 295398
rect 353868 295954 354868 295986
rect 353868 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 354868 295954
rect 353868 295634 354868 295718
rect 353868 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 354868 295634
rect 353868 295366 354868 295398
rect 373868 295954 374868 295986
rect 373868 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 374868 295954
rect 373868 295634 374868 295718
rect 373868 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 374868 295634
rect 373868 295366 374868 295398
rect 393868 295954 394868 295986
rect 393868 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 394868 295954
rect 393868 295634 394868 295718
rect 393868 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 394868 295634
rect 393868 295366 394868 295398
rect 413868 295954 414868 295986
rect 413868 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 414868 295954
rect 413868 295634 414868 295718
rect 413868 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 414868 295634
rect 413868 295366 414868 295398
rect 433868 295954 434868 295986
rect 433868 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 434868 295954
rect 433868 295634 434868 295718
rect 433868 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 434868 295634
rect 433868 295366 434868 295398
rect 453868 295954 454868 295986
rect 453868 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 454868 295954
rect 453868 295634 454868 295718
rect 453868 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 454868 295634
rect 453868 295366 454868 295398
rect 473868 295954 474868 295986
rect 473868 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 474868 295954
rect 473868 295634 474868 295718
rect 473868 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 474868 295634
rect 473868 295366 474868 295398
rect 493868 295954 494868 295986
rect 493868 295718 493930 295954
rect 494166 295718 494250 295954
rect 494486 295718 494570 295954
rect 494806 295718 494868 295954
rect 493868 295634 494868 295718
rect 493868 295398 493930 295634
rect 494166 295398 494250 295634
rect 494486 295398 494570 295634
rect 494806 295398 494868 295634
rect 493868 295366 494868 295398
rect 513868 295954 514868 295986
rect 513868 295718 513930 295954
rect 514166 295718 514250 295954
rect 514486 295718 514570 295954
rect 514806 295718 514868 295954
rect 513868 295634 514868 295718
rect 513868 295398 513930 295634
rect 514166 295398 514250 295634
rect 514486 295398 514570 295634
rect 514806 295398 514868 295634
rect 513868 295366 514868 295398
rect 533868 295954 534868 295986
rect 533868 295718 533930 295954
rect 534166 295718 534250 295954
rect 534486 295718 534570 295954
rect 534806 295718 534868 295954
rect 533868 295634 534868 295718
rect 533868 295398 533930 295634
rect 534166 295398 534250 295634
rect 534486 295398 534570 295634
rect 534806 295398 534868 295634
rect 533868 295366 534868 295398
rect 553868 295954 554868 295986
rect 553868 295718 553930 295954
rect 554166 295718 554250 295954
rect 554486 295718 554570 295954
rect 554806 295718 554868 295954
rect 553868 295634 554868 295718
rect 553868 295398 553930 295634
rect 554166 295398 554250 295634
rect 554486 295398 554570 295634
rect 554806 295398 554868 295634
rect 553868 295366 554868 295398
rect 303868 291454 304868 291486
rect 303868 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 304868 291454
rect 303868 291134 304868 291218
rect 303868 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 304868 291134
rect 303868 290866 304868 290898
rect 323868 291454 324868 291486
rect 323868 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 324868 291454
rect 323868 291134 324868 291218
rect 323868 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 324868 291134
rect 323868 290866 324868 290898
rect 343868 291454 344868 291486
rect 343868 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 344868 291454
rect 343868 291134 344868 291218
rect 343868 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 344868 291134
rect 343868 290866 344868 290898
rect 363868 291454 364868 291486
rect 363868 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 364868 291454
rect 363868 291134 364868 291218
rect 363868 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 364868 291134
rect 363868 290866 364868 290898
rect 383868 291454 384868 291486
rect 383868 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 384868 291454
rect 383868 291134 384868 291218
rect 383868 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 384868 291134
rect 383868 290866 384868 290898
rect 403868 291454 404868 291486
rect 403868 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 404868 291454
rect 403868 291134 404868 291218
rect 403868 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 404868 291134
rect 403868 290866 404868 290898
rect 423868 291454 424868 291486
rect 423868 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 424868 291454
rect 423868 291134 424868 291218
rect 423868 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 424868 291134
rect 423868 290866 424868 290898
rect 443868 291454 444868 291486
rect 443868 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 444868 291454
rect 443868 291134 444868 291218
rect 443868 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 444868 291134
rect 443868 290866 444868 290898
rect 463868 291454 464868 291486
rect 463868 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 464868 291454
rect 463868 291134 464868 291218
rect 463868 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 464868 291134
rect 463868 290866 464868 290898
rect 483868 291454 484868 291486
rect 483868 291218 483930 291454
rect 484166 291218 484250 291454
rect 484486 291218 484570 291454
rect 484806 291218 484868 291454
rect 483868 291134 484868 291218
rect 483868 290898 483930 291134
rect 484166 290898 484250 291134
rect 484486 290898 484570 291134
rect 484806 290898 484868 291134
rect 483868 290866 484868 290898
rect 503868 291454 504868 291486
rect 503868 291218 503930 291454
rect 504166 291218 504250 291454
rect 504486 291218 504570 291454
rect 504806 291218 504868 291454
rect 503868 291134 504868 291218
rect 503868 290898 503930 291134
rect 504166 290898 504250 291134
rect 504486 290898 504570 291134
rect 504806 290898 504868 291134
rect 503868 290866 504868 290898
rect 523868 291454 524868 291486
rect 523868 291218 523930 291454
rect 524166 291218 524250 291454
rect 524486 291218 524570 291454
rect 524806 291218 524868 291454
rect 523868 291134 524868 291218
rect 523868 290898 523930 291134
rect 524166 290898 524250 291134
rect 524486 290898 524570 291134
rect 524806 290898 524868 291134
rect 523868 290866 524868 290898
rect 543868 291454 544868 291486
rect 543868 291218 543930 291454
rect 544166 291218 544250 291454
rect 544486 291218 544570 291454
rect 544806 291218 544868 291454
rect 543868 291134 544868 291218
rect 543868 290898 543930 291134
rect 544166 290898 544250 291134
rect 544486 290898 544570 291134
rect 544806 290898 544868 291134
rect 543868 290866 544868 290898
rect 563868 291454 564868 291486
rect 563868 291218 563930 291454
rect 564166 291218 564250 291454
rect 564486 291218 564570 291454
rect 564806 291218 564868 291454
rect 563868 291134 564868 291218
rect 563868 290898 563930 291134
rect 564166 290898 564250 291134
rect 564486 290898 564570 291134
rect 564806 290898 564868 291134
rect 563868 290866 564868 290898
rect 313868 259954 314868 259986
rect 313868 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 314868 259954
rect 313868 259634 314868 259718
rect 313868 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 314868 259634
rect 313868 259366 314868 259398
rect 333868 259954 334868 259986
rect 333868 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 334868 259954
rect 333868 259634 334868 259718
rect 333868 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 334868 259634
rect 333868 259366 334868 259398
rect 353868 259954 354868 259986
rect 353868 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 354868 259954
rect 353868 259634 354868 259718
rect 353868 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 354868 259634
rect 353868 259366 354868 259398
rect 373868 259954 374868 259986
rect 373868 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 374868 259954
rect 373868 259634 374868 259718
rect 373868 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 374868 259634
rect 373868 259366 374868 259398
rect 393868 259954 394868 259986
rect 393868 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 394868 259954
rect 393868 259634 394868 259718
rect 393868 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 394868 259634
rect 393868 259366 394868 259398
rect 413868 259954 414868 259986
rect 413868 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 414868 259954
rect 413868 259634 414868 259718
rect 413868 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 414868 259634
rect 413868 259366 414868 259398
rect 433868 259954 434868 259986
rect 433868 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 434868 259954
rect 433868 259634 434868 259718
rect 433868 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 434868 259634
rect 433868 259366 434868 259398
rect 453868 259954 454868 259986
rect 453868 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 454868 259954
rect 453868 259634 454868 259718
rect 453868 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 454868 259634
rect 453868 259366 454868 259398
rect 473868 259954 474868 259986
rect 473868 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 474868 259954
rect 473868 259634 474868 259718
rect 473868 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 474868 259634
rect 473868 259366 474868 259398
rect 493868 259954 494868 259986
rect 493868 259718 493930 259954
rect 494166 259718 494250 259954
rect 494486 259718 494570 259954
rect 494806 259718 494868 259954
rect 493868 259634 494868 259718
rect 493868 259398 493930 259634
rect 494166 259398 494250 259634
rect 494486 259398 494570 259634
rect 494806 259398 494868 259634
rect 493868 259366 494868 259398
rect 513868 259954 514868 259986
rect 513868 259718 513930 259954
rect 514166 259718 514250 259954
rect 514486 259718 514570 259954
rect 514806 259718 514868 259954
rect 513868 259634 514868 259718
rect 513868 259398 513930 259634
rect 514166 259398 514250 259634
rect 514486 259398 514570 259634
rect 514806 259398 514868 259634
rect 513868 259366 514868 259398
rect 533868 259954 534868 259986
rect 533868 259718 533930 259954
rect 534166 259718 534250 259954
rect 534486 259718 534570 259954
rect 534806 259718 534868 259954
rect 533868 259634 534868 259718
rect 533868 259398 533930 259634
rect 534166 259398 534250 259634
rect 534486 259398 534570 259634
rect 534806 259398 534868 259634
rect 533868 259366 534868 259398
rect 553868 259954 554868 259986
rect 553868 259718 553930 259954
rect 554166 259718 554250 259954
rect 554486 259718 554570 259954
rect 554806 259718 554868 259954
rect 553868 259634 554868 259718
rect 553868 259398 553930 259634
rect 554166 259398 554250 259634
rect 554486 259398 554570 259634
rect 554806 259398 554868 259634
rect 553868 259366 554868 259398
rect 303868 255454 304868 255486
rect 303868 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 304868 255454
rect 303868 255134 304868 255218
rect 303868 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 304868 255134
rect 303868 254866 304868 254898
rect 323868 255454 324868 255486
rect 323868 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 324868 255454
rect 323868 255134 324868 255218
rect 323868 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 324868 255134
rect 323868 254866 324868 254898
rect 343868 255454 344868 255486
rect 343868 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 344868 255454
rect 343868 255134 344868 255218
rect 343868 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 344868 255134
rect 343868 254866 344868 254898
rect 363868 255454 364868 255486
rect 363868 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 364868 255454
rect 363868 255134 364868 255218
rect 363868 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 364868 255134
rect 363868 254866 364868 254898
rect 383868 255454 384868 255486
rect 383868 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 384868 255454
rect 383868 255134 384868 255218
rect 383868 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 384868 255134
rect 383868 254866 384868 254898
rect 403868 255454 404868 255486
rect 403868 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 404868 255454
rect 403868 255134 404868 255218
rect 403868 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 404868 255134
rect 403868 254866 404868 254898
rect 423868 255454 424868 255486
rect 423868 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 424868 255454
rect 423868 255134 424868 255218
rect 423868 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 424868 255134
rect 423868 254866 424868 254898
rect 443868 255454 444868 255486
rect 443868 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 444868 255454
rect 443868 255134 444868 255218
rect 443868 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 444868 255134
rect 443868 254866 444868 254898
rect 463868 255454 464868 255486
rect 463868 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 464868 255454
rect 463868 255134 464868 255218
rect 463868 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 464868 255134
rect 463868 254866 464868 254898
rect 483868 255454 484868 255486
rect 483868 255218 483930 255454
rect 484166 255218 484250 255454
rect 484486 255218 484570 255454
rect 484806 255218 484868 255454
rect 483868 255134 484868 255218
rect 483868 254898 483930 255134
rect 484166 254898 484250 255134
rect 484486 254898 484570 255134
rect 484806 254898 484868 255134
rect 483868 254866 484868 254898
rect 503868 255454 504868 255486
rect 503868 255218 503930 255454
rect 504166 255218 504250 255454
rect 504486 255218 504570 255454
rect 504806 255218 504868 255454
rect 503868 255134 504868 255218
rect 503868 254898 503930 255134
rect 504166 254898 504250 255134
rect 504486 254898 504570 255134
rect 504806 254898 504868 255134
rect 503868 254866 504868 254898
rect 523868 255454 524868 255486
rect 523868 255218 523930 255454
rect 524166 255218 524250 255454
rect 524486 255218 524570 255454
rect 524806 255218 524868 255454
rect 523868 255134 524868 255218
rect 523868 254898 523930 255134
rect 524166 254898 524250 255134
rect 524486 254898 524570 255134
rect 524806 254898 524868 255134
rect 523868 254866 524868 254898
rect 543868 255454 544868 255486
rect 543868 255218 543930 255454
rect 544166 255218 544250 255454
rect 544486 255218 544570 255454
rect 544806 255218 544868 255454
rect 543868 255134 544868 255218
rect 543868 254898 543930 255134
rect 544166 254898 544250 255134
rect 544486 254898 544570 255134
rect 544806 254898 544868 255134
rect 543868 254866 544868 254898
rect 563868 255454 564868 255486
rect 563868 255218 563930 255454
rect 564166 255218 564250 255454
rect 564486 255218 564570 255454
rect 564806 255218 564868 255454
rect 563868 255134 564868 255218
rect 563868 254898 563930 255134
rect 564166 254898 564250 255134
rect 564486 254898 564570 255134
rect 564806 254898 564868 255134
rect 563868 254866 564868 254898
rect 313868 223954 314868 223986
rect 313868 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 314868 223954
rect 313868 223634 314868 223718
rect 313868 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 314868 223634
rect 313868 223366 314868 223398
rect 333868 223954 334868 223986
rect 333868 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 334868 223954
rect 333868 223634 334868 223718
rect 333868 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 334868 223634
rect 333868 223366 334868 223398
rect 353868 223954 354868 223986
rect 353868 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 354868 223954
rect 353868 223634 354868 223718
rect 353868 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 354868 223634
rect 353868 223366 354868 223398
rect 373868 223954 374868 223986
rect 373868 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 374868 223954
rect 373868 223634 374868 223718
rect 373868 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 374868 223634
rect 373868 223366 374868 223398
rect 393868 223954 394868 223986
rect 393868 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 394868 223954
rect 393868 223634 394868 223718
rect 393868 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 394868 223634
rect 393868 223366 394868 223398
rect 413868 223954 414868 223986
rect 413868 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 414868 223954
rect 413868 223634 414868 223718
rect 413868 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 414868 223634
rect 413868 223366 414868 223398
rect 433868 223954 434868 223986
rect 433868 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 434868 223954
rect 433868 223634 434868 223718
rect 433868 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 434868 223634
rect 433868 223366 434868 223398
rect 453868 223954 454868 223986
rect 453868 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 454868 223954
rect 453868 223634 454868 223718
rect 453868 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 454868 223634
rect 453868 223366 454868 223398
rect 473868 223954 474868 223986
rect 473868 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 474868 223954
rect 473868 223634 474868 223718
rect 473868 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 474868 223634
rect 473868 223366 474868 223398
rect 493868 223954 494868 223986
rect 493868 223718 493930 223954
rect 494166 223718 494250 223954
rect 494486 223718 494570 223954
rect 494806 223718 494868 223954
rect 493868 223634 494868 223718
rect 493868 223398 493930 223634
rect 494166 223398 494250 223634
rect 494486 223398 494570 223634
rect 494806 223398 494868 223634
rect 493868 223366 494868 223398
rect 513868 223954 514868 223986
rect 513868 223718 513930 223954
rect 514166 223718 514250 223954
rect 514486 223718 514570 223954
rect 514806 223718 514868 223954
rect 513868 223634 514868 223718
rect 513868 223398 513930 223634
rect 514166 223398 514250 223634
rect 514486 223398 514570 223634
rect 514806 223398 514868 223634
rect 513868 223366 514868 223398
rect 533868 223954 534868 223986
rect 533868 223718 533930 223954
rect 534166 223718 534250 223954
rect 534486 223718 534570 223954
rect 534806 223718 534868 223954
rect 533868 223634 534868 223718
rect 533868 223398 533930 223634
rect 534166 223398 534250 223634
rect 534486 223398 534570 223634
rect 534806 223398 534868 223634
rect 533868 223366 534868 223398
rect 553868 223954 554868 223986
rect 553868 223718 553930 223954
rect 554166 223718 554250 223954
rect 554486 223718 554570 223954
rect 554806 223718 554868 223954
rect 553868 223634 554868 223718
rect 553868 223398 553930 223634
rect 554166 223398 554250 223634
rect 554486 223398 554570 223634
rect 554806 223398 554868 223634
rect 553868 223366 554868 223398
rect 303868 219454 304868 219486
rect 303868 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 304868 219454
rect 303868 219134 304868 219218
rect 303868 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 304868 219134
rect 303868 218866 304868 218898
rect 323868 219454 324868 219486
rect 323868 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 324868 219454
rect 323868 219134 324868 219218
rect 323868 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 324868 219134
rect 323868 218866 324868 218898
rect 343868 219454 344868 219486
rect 343868 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 344868 219454
rect 343868 219134 344868 219218
rect 343868 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 344868 219134
rect 343868 218866 344868 218898
rect 363868 219454 364868 219486
rect 363868 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 364868 219454
rect 363868 219134 364868 219218
rect 363868 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 364868 219134
rect 363868 218866 364868 218898
rect 383868 219454 384868 219486
rect 383868 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 384868 219454
rect 383868 219134 384868 219218
rect 383868 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 384868 219134
rect 383868 218866 384868 218898
rect 403868 219454 404868 219486
rect 403868 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 404868 219454
rect 403868 219134 404868 219218
rect 403868 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 404868 219134
rect 403868 218866 404868 218898
rect 423868 219454 424868 219486
rect 423868 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 424868 219454
rect 423868 219134 424868 219218
rect 423868 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 424868 219134
rect 423868 218866 424868 218898
rect 443868 219454 444868 219486
rect 443868 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 444868 219454
rect 443868 219134 444868 219218
rect 443868 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 444868 219134
rect 443868 218866 444868 218898
rect 463868 219454 464868 219486
rect 463868 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 464868 219454
rect 463868 219134 464868 219218
rect 463868 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 464868 219134
rect 463868 218866 464868 218898
rect 483868 219454 484868 219486
rect 483868 219218 483930 219454
rect 484166 219218 484250 219454
rect 484486 219218 484570 219454
rect 484806 219218 484868 219454
rect 483868 219134 484868 219218
rect 483868 218898 483930 219134
rect 484166 218898 484250 219134
rect 484486 218898 484570 219134
rect 484806 218898 484868 219134
rect 483868 218866 484868 218898
rect 503868 219454 504868 219486
rect 503868 219218 503930 219454
rect 504166 219218 504250 219454
rect 504486 219218 504570 219454
rect 504806 219218 504868 219454
rect 503868 219134 504868 219218
rect 503868 218898 503930 219134
rect 504166 218898 504250 219134
rect 504486 218898 504570 219134
rect 504806 218898 504868 219134
rect 503868 218866 504868 218898
rect 523868 219454 524868 219486
rect 523868 219218 523930 219454
rect 524166 219218 524250 219454
rect 524486 219218 524570 219454
rect 524806 219218 524868 219454
rect 523868 219134 524868 219218
rect 523868 218898 523930 219134
rect 524166 218898 524250 219134
rect 524486 218898 524570 219134
rect 524806 218898 524868 219134
rect 523868 218866 524868 218898
rect 543868 219454 544868 219486
rect 543868 219218 543930 219454
rect 544166 219218 544250 219454
rect 544486 219218 544570 219454
rect 544806 219218 544868 219454
rect 543868 219134 544868 219218
rect 543868 218898 543930 219134
rect 544166 218898 544250 219134
rect 544486 218898 544570 219134
rect 544806 218898 544868 219134
rect 543868 218866 544868 218898
rect 563868 219454 564868 219486
rect 563868 219218 563930 219454
rect 564166 219218 564250 219454
rect 564486 219218 564570 219454
rect 564806 219218 564868 219454
rect 563868 219134 564868 219218
rect 563868 218898 563930 219134
rect 564166 218898 564250 219134
rect 564486 218898 564570 219134
rect 564806 218898 564868 219134
rect 563868 218866 564868 218898
rect 303475 205596 303541 205597
rect 303475 205532 303476 205596
rect 303540 205532 303541 205596
rect 303475 205531 303541 205532
rect 303475 188324 303541 188325
rect 303475 188260 303476 188324
rect 303540 188260 303541 188324
rect 303475 188259 303541 188260
rect 303478 77893 303538 188259
rect 303868 183454 304868 183486
rect 303868 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 304868 183454
rect 303868 183134 304868 183218
rect 303868 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 304868 183134
rect 303868 182866 304868 182898
rect 323868 183454 324868 183486
rect 323868 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 324868 183454
rect 323868 183134 324868 183218
rect 323868 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 324868 183134
rect 323868 182866 324868 182898
rect 343868 183454 344868 183486
rect 343868 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 344868 183454
rect 343868 183134 344868 183218
rect 343868 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 344868 183134
rect 343868 182866 344868 182898
rect 363868 183454 364868 183486
rect 363868 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 364868 183454
rect 363868 183134 364868 183218
rect 363868 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 364868 183134
rect 363868 182866 364868 182898
rect 383868 183454 384868 183486
rect 383868 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 384868 183454
rect 383868 183134 384868 183218
rect 383868 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 384868 183134
rect 383868 182866 384868 182898
rect 403868 183454 404868 183486
rect 403868 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 404868 183454
rect 403868 183134 404868 183218
rect 403868 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 404868 183134
rect 403868 182866 404868 182898
rect 423868 183454 424868 183486
rect 423868 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 424868 183454
rect 423868 183134 424868 183218
rect 423868 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 424868 183134
rect 423868 182866 424868 182898
rect 443868 183454 444868 183486
rect 443868 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 444868 183454
rect 443868 183134 444868 183218
rect 443868 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 444868 183134
rect 443868 182866 444868 182898
rect 463868 183454 464868 183486
rect 463868 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 464868 183454
rect 463868 183134 464868 183218
rect 463868 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 464868 183134
rect 463868 182866 464868 182898
rect 483868 183454 484868 183486
rect 483868 183218 483930 183454
rect 484166 183218 484250 183454
rect 484486 183218 484570 183454
rect 484806 183218 484868 183454
rect 483868 183134 484868 183218
rect 483868 182898 483930 183134
rect 484166 182898 484250 183134
rect 484486 182898 484570 183134
rect 484806 182898 484868 183134
rect 483868 182866 484868 182898
rect 503868 183454 504868 183486
rect 503868 183218 503930 183454
rect 504166 183218 504250 183454
rect 504486 183218 504570 183454
rect 504806 183218 504868 183454
rect 503868 183134 504868 183218
rect 503868 182898 503930 183134
rect 504166 182898 504250 183134
rect 504486 182898 504570 183134
rect 504806 182898 504868 183134
rect 503868 182866 504868 182898
rect 523868 183454 524868 183486
rect 523868 183218 523930 183454
rect 524166 183218 524250 183454
rect 524486 183218 524570 183454
rect 524806 183218 524868 183454
rect 523868 183134 524868 183218
rect 523868 182898 523930 183134
rect 524166 182898 524250 183134
rect 524486 182898 524570 183134
rect 524806 182898 524868 183134
rect 523868 182866 524868 182898
rect 543868 183454 544868 183486
rect 543868 183218 543930 183454
rect 544166 183218 544250 183454
rect 544486 183218 544570 183454
rect 544806 183218 544868 183454
rect 543868 183134 544868 183218
rect 543868 182898 543930 183134
rect 544166 182898 544250 183134
rect 544486 182898 544570 183134
rect 544806 182898 544868 183134
rect 543868 182866 544868 182898
rect 563868 183454 564868 183486
rect 563868 183218 563930 183454
rect 564166 183218 564250 183454
rect 564486 183218 564570 183454
rect 564806 183218 564868 183454
rect 563868 183134 564868 183218
rect 563868 182898 563930 183134
rect 564166 182898 564250 183134
rect 564486 182898 564570 183134
rect 564806 182898 564868 183134
rect 563868 182866 564868 182898
rect 313868 151954 314868 151986
rect 313868 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 314868 151954
rect 313868 151634 314868 151718
rect 313868 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 314868 151634
rect 313868 151366 314868 151398
rect 333868 151954 334868 151986
rect 333868 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 334868 151954
rect 333868 151634 334868 151718
rect 333868 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 334868 151634
rect 333868 151366 334868 151398
rect 353868 151954 354868 151986
rect 353868 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 354868 151954
rect 353868 151634 354868 151718
rect 353868 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 354868 151634
rect 353868 151366 354868 151398
rect 373868 151954 374868 151986
rect 373868 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 374868 151954
rect 373868 151634 374868 151718
rect 373868 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 374868 151634
rect 373868 151366 374868 151398
rect 393868 151954 394868 151986
rect 393868 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 394868 151954
rect 393868 151634 394868 151718
rect 393868 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 394868 151634
rect 393868 151366 394868 151398
rect 413868 151954 414868 151986
rect 413868 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 414868 151954
rect 413868 151634 414868 151718
rect 413868 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 414868 151634
rect 413868 151366 414868 151398
rect 433868 151954 434868 151986
rect 433868 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 434868 151954
rect 433868 151634 434868 151718
rect 433868 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 434868 151634
rect 433868 151366 434868 151398
rect 453868 151954 454868 151986
rect 453868 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 454868 151954
rect 453868 151634 454868 151718
rect 453868 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 454868 151634
rect 453868 151366 454868 151398
rect 473868 151954 474868 151986
rect 473868 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 474868 151954
rect 473868 151634 474868 151718
rect 473868 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 474868 151634
rect 473868 151366 474868 151398
rect 493868 151954 494868 151986
rect 493868 151718 493930 151954
rect 494166 151718 494250 151954
rect 494486 151718 494570 151954
rect 494806 151718 494868 151954
rect 493868 151634 494868 151718
rect 493868 151398 493930 151634
rect 494166 151398 494250 151634
rect 494486 151398 494570 151634
rect 494806 151398 494868 151634
rect 493868 151366 494868 151398
rect 513868 151954 514868 151986
rect 513868 151718 513930 151954
rect 514166 151718 514250 151954
rect 514486 151718 514570 151954
rect 514806 151718 514868 151954
rect 513868 151634 514868 151718
rect 513868 151398 513930 151634
rect 514166 151398 514250 151634
rect 514486 151398 514570 151634
rect 514806 151398 514868 151634
rect 513868 151366 514868 151398
rect 533868 151954 534868 151986
rect 533868 151718 533930 151954
rect 534166 151718 534250 151954
rect 534486 151718 534570 151954
rect 534806 151718 534868 151954
rect 533868 151634 534868 151718
rect 533868 151398 533930 151634
rect 534166 151398 534250 151634
rect 534486 151398 534570 151634
rect 534806 151398 534868 151634
rect 533868 151366 534868 151398
rect 553868 151954 554868 151986
rect 553868 151718 553930 151954
rect 554166 151718 554250 151954
rect 554486 151718 554570 151954
rect 554806 151718 554868 151954
rect 553868 151634 554868 151718
rect 553868 151398 553930 151634
rect 554166 151398 554250 151634
rect 554486 151398 554570 151634
rect 554806 151398 554868 151634
rect 553868 151366 554868 151398
rect 303868 147454 304868 147486
rect 303868 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 304868 147454
rect 303868 147134 304868 147218
rect 303868 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 304868 147134
rect 303868 146866 304868 146898
rect 323868 147454 324868 147486
rect 323868 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 324868 147454
rect 323868 147134 324868 147218
rect 323868 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 324868 147134
rect 323868 146866 324868 146898
rect 343868 147454 344868 147486
rect 343868 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 344868 147454
rect 343868 147134 344868 147218
rect 343868 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 344868 147134
rect 343868 146866 344868 146898
rect 363868 147454 364868 147486
rect 363868 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 364868 147454
rect 363868 147134 364868 147218
rect 363868 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 364868 147134
rect 363868 146866 364868 146898
rect 383868 147454 384868 147486
rect 383868 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 384868 147454
rect 383868 147134 384868 147218
rect 383868 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 384868 147134
rect 383868 146866 384868 146898
rect 403868 147454 404868 147486
rect 403868 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 404868 147454
rect 403868 147134 404868 147218
rect 403868 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 404868 147134
rect 403868 146866 404868 146898
rect 423868 147454 424868 147486
rect 423868 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 424868 147454
rect 423868 147134 424868 147218
rect 423868 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 424868 147134
rect 423868 146866 424868 146898
rect 443868 147454 444868 147486
rect 443868 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 444868 147454
rect 443868 147134 444868 147218
rect 443868 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 444868 147134
rect 443868 146866 444868 146898
rect 463868 147454 464868 147486
rect 463868 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 464868 147454
rect 463868 147134 464868 147218
rect 463868 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 464868 147134
rect 463868 146866 464868 146898
rect 483868 147454 484868 147486
rect 483868 147218 483930 147454
rect 484166 147218 484250 147454
rect 484486 147218 484570 147454
rect 484806 147218 484868 147454
rect 483868 147134 484868 147218
rect 483868 146898 483930 147134
rect 484166 146898 484250 147134
rect 484486 146898 484570 147134
rect 484806 146898 484868 147134
rect 483868 146866 484868 146898
rect 503868 147454 504868 147486
rect 503868 147218 503930 147454
rect 504166 147218 504250 147454
rect 504486 147218 504570 147454
rect 504806 147218 504868 147454
rect 503868 147134 504868 147218
rect 503868 146898 503930 147134
rect 504166 146898 504250 147134
rect 504486 146898 504570 147134
rect 504806 146898 504868 147134
rect 503868 146866 504868 146898
rect 523868 147454 524868 147486
rect 523868 147218 523930 147454
rect 524166 147218 524250 147454
rect 524486 147218 524570 147454
rect 524806 147218 524868 147454
rect 523868 147134 524868 147218
rect 523868 146898 523930 147134
rect 524166 146898 524250 147134
rect 524486 146898 524570 147134
rect 524806 146898 524868 147134
rect 523868 146866 524868 146898
rect 543868 147454 544868 147486
rect 543868 147218 543930 147454
rect 544166 147218 544250 147454
rect 544486 147218 544570 147454
rect 544806 147218 544868 147454
rect 543868 147134 544868 147218
rect 543868 146898 543930 147134
rect 544166 146898 544250 147134
rect 544486 146898 544570 147134
rect 544806 146898 544868 147134
rect 543868 146866 544868 146898
rect 563868 147454 564868 147486
rect 563868 147218 563930 147454
rect 564166 147218 564250 147454
rect 564486 147218 564570 147454
rect 564806 147218 564868 147454
rect 563868 147134 564868 147218
rect 563868 146898 563930 147134
rect 564166 146898 564250 147134
rect 564486 146898 564570 147134
rect 564806 146898 564868 147134
rect 563868 146866 564868 146898
rect 313868 115954 314868 115986
rect 313868 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 314868 115954
rect 313868 115634 314868 115718
rect 313868 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 314868 115634
rect 313868 115366 314868 115398
rect 333868 115954 334868 115986
rect 333868 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 334868 115954
rect 333868 115634 334868 115718
rect 333868 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 334868 115634
rect 333868 115366 334868 115398
rect 353868 115954 354868 115986
rect 353868 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 354868 115954
rect 353868 115634 354868 115718
rect 353868 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 354868 115634
rect 353868 115366 354868 115398
rect 373868 115954 374868 115986
rect 373868 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 374868 115954
rect 373868 115634 374868 115718
rect 373868 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 374868 115634
rect 373868 115366 374868 115398
rect 393868 115954 394868 115986
rect 393868 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 394868 115954
rect 393868 115634 394868 115718
rect 393868 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 394868 115634
rect 393868 115366 394868 115398
rect 413868 115954 414868 115986
rect 413868 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 414868 115954
rect 413868 115634 414868 115718
rect 413868 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 414868 115634
rect 413868 115366 414868 115398
rect 433868 115954 434868 115986
rect 433868 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 434868 115954
rect 433868 115634 434868 115718
rect 433868 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 434868 115634
rect 433868 115366 434868 115398
rect 453868 115954 454868 115986
rect 453868 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 454868 115954
rect 453868 115634 454868 115718
rect 453868 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 454868 115634
rect 453868 115366 454868 115398
rect 473868 115954 474868 115986
rect 473868 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 474868 115954
rect 473868 115634 474868 115718
rect 473868 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 474868 115634
rect 473868 115366 474868 115398
rect 493868 115954 494868 115986
rect 493868 115718 493930 115954
rect 494166 115718 494250 115954
rect 494486 115718 494570 115954
rect 494806 115718 494868 115954
rect 493868 115634 494868 115718
rect 493868 115398 493930 115634
rect 494166 115398 494250 115634
rect 494486 115398 494570 115634
rect 494806 115398 494868 115634
rect 493868 115366 494868 115398
rect 513868 115954 514868 115986
rect 513868 115718 513930 115954
rect 514166 115718 514250 115954
rect 514486 115718 514570 115954
rect 514806 115718 514868 115954
rect 513868 115634 514868 115718
rect 513868 115398 513930 115634
rect 514166 115398 514250 115634
rect 514486 115398 514570 115634
rect 514806 115398 514868 115634
rect 513868 115366 514868 115398
rect 533868 115954 534868 115986
rect 533868 115718 533930 115954
rect 534166 115718 534250 115954
rect 534486 115718 534570 115954
rect 534806 115718 534868 115954
rect 533868 115634 534868 115718
rect 533868 115398 533930 115634
rect 534166 115398 534250 115634
rect 534486 115398 534570 115634
rect 534806 115398 534868 115634
rect 533868 115366 534868 115398
rect 553868 115954 554868 115986
rect 553868 115718 553930 115954
rect 554166 115718 554250 115954
rect 554486 115718 554570 115954
rect 554806 115718 554868 115954
rect 553868 115634 554868 115718
rect 553868 115398 553930 115634
rect 554166 115398 554250 115634
rect 554486 115398 554570 115634
rect 554806 115398 554868 115634
rect 553868 115366 554868 115398
rect 303868 111454 304868 111486
rect 303868 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 304868 111454
rect 303868 111134 304868 111218
rect 303868 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 304868 111134
rect 303868 110866 304868 110898
rect 323868 111454 324868 111486
rect 323868 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 324868 111454
rect 323868 111134 324868 111218
rect 323868 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 324868 111134
rect 323868 110866 324868 110898
rect 343868 111454 344868 111486
rect 343868 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 344868 111454
rect 343868 111134 344868 111218
rect 343868 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 344868 111134
rect 343868 110866 344868 110898
rect 363868 111454 364868 111486
rect 363868 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 364868 111454
rect 363868 111134 364868 111218
rect 363868 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 364868 111134
rect 363868 110866 364868 110898
rect 383868 111454 384868 111486
rect 383868 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 384868 111454
rect 383868 111134 384868 111218
rect 383868 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 384868 111134
rect 383868 110866 384868 110898
rect 403868 111454 404868 111486
rect 403868 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 404868 111454
rect 403868 111134 404868 111218
rect 403868 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 404868 111134
rect 403868 110866 404868 110898
rect 423868 111454 424868 111486
rect 423868 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 424868 111454
rect 423868 111134 424868 111218
rect 423868 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 424868 111134
rect 423868 110866 424868 110898
rect 443868 111454 444868 111486
rect 443868 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 444868 111454
rect 443868 111134 444868 111218
rect 443868 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 444868 111134
rect 443868 110866 444868 110898
rect 463868 111454 464868 111486
rect 463868 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 464868 111454
rect 463868 111134 464868 111218
rect 463868 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 464868 111134
rect 463868 110866 464868 110898
rect 483868 111454 484868 111486
rect 483868 111218 483930 111454
rect 484166 111218 484250 111454
rect 484486 111218 484570 111454
rect 484806 111218 484868 111454
rect 483868 111134 484868 111218
rect 483868 110898 483930 111134
rect 484166 110898 484250 111134
rect 484486 110898 484570 111134
rect 484806 110898 484868 111134
rect 483868 110866 484868 110898
rect 503868 111454 504868 111486
rect 503868 111218 503930 111454
rect 504166 111218 504250 111454
rect 504486 111218 504570 111454
rect 504806 111218 504868 111454
rect 503868 111134 504868 111218
rect 503868 110898 503930 111134
rect 504166 110898 504250 111134
rect 504486 110898 504570 111134
rect 504806 110898 504868 111134
rect 503868 110866 504868 110898
rect 523868 111454 524868 111486
rect 523868 111218 523930 111454
rect 524166 111218 524250 111454
rect 524486 111218 524570 111454
rect 524806 111218 524868 111454
rect 523868 111134 524868 111218
rect 523868 110898 523930 111134
rect 524166 110898 524250 111134
rect 524486 110898 524570 111134
rect 524806 110898 524868 111134
rect 523868 110866 524868 110898
rect 543868 111454 544868 111486
rect 543868 111218 543930 111454
rect 544166 111218 544250 111454
rect 544486 111218 544570 111454
rect 544806 111218 544868 111454
rect 543868 111134 544868 111218
rect 543868 110898 543930 111134
rect 544166 110898 544250 111134
rect 544486 110898 544570 111134
rect 544806 110898 544868 111134
rect 543868 110866 544868 110898
rect 563868 111454 564868 111486
rect 563868 111218 563930 111454
rect 564166 111218 564250 111454
rect 564486 111218 564570 111454
rect 564806 111218 564868 111454
rect 563868 111134 564868 111218
rect 563868 110898 563930 111134
rect 564166 110898 564250 111134
rect 564486 110898 564570 111134
rect 564806 110898 564868 111134
rect 563868 110866 564868 110898
rect 565307 79388 565373 79389
rect 565307 79324 565308 79388
rect 565372 79324 565373 79388
rect 565307 79323 565373 79324
rect 303475 77892 303541 77893
rect 303475 77828 303476 77892
rect 303540 77828 303541 77892
rect 303475 77827 303541 77828
rect 302739 76804 302805 76805
rect 302739 76740 302740 76804
rect 302804 76740 302805 76804
rect 302739 76739 302805 76740
rect 301635 76668 301701 76669
rect 301635 76604 301636 76668
rect 301700 76604 301701 76668
rect 301635 76603 301701 76604
rect 300163 54500 300229 54501
rect 300163 54436 300164 54500
rect 300228 54436 300229 54500
rect 300163 54435 300229 54436
rect 288939 53140 289005 53141
rect 288939 53076 288940 53140
rect 289004 53076 289005 53140
rect 288939 53075 289005 53076
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 167868 43954 168868 43986
rect 167868 43718 167930 43954
rect 168166 43718 168250 43954
rect 168486 43718 168570 43954
rect 168806 43718 168868 43954
rect 167868 43634 168868 43718
rect 167868 43398 167930 43634
rect 168166 43398 168250 43634
rect 168486 43398 168570 43634
rect 168806 43398 168868 43634
rect 167868 43366 168868 43398
rect 187868 43954 188868 43986
rect 187868 43718 187930 43954
rect 188166 43718 188250 43954
rect 188486 43718 188570 43954
rect 188806 43718 188868 43954
rect 187868 43634 188868 43718
rect 187868 43398 187930 43634
rect 188166 43398 188250 43634
rect 188486 43398 188570 43634
rect 188806 43398 188868 43634
rect 187868 43366 188868 43398
rect 207868 43954 208868 43986
rect 207868 43718 207930 43954
rect 208166 43718 208250 43954
rect 208486 43718 208570 43954
rect 208806 43718 208868 43954
rect 207868 43634 208868 43718
rect 207868 43398 207930 43634
rect 208166 43398 208250 43634
rect 208486 43398 208570 43634
rect 208806 43398 208868 43634
rect 207868 43366 208868 43398
rect 227868 43954 228868 43986
rect 227868 43718 227930 43954
rect 228166 43718 228250 43954
rect 228486 43718 228570 43954
rect 228806 43718 228868 43954
rect 227868 43634 228868 43718
rect 227868 43398 227930 43634
rect 228166 43398 228250 43634
rect 228486 43398 228570 43634
rect 228806 43398 228868 43634
rect 227868 43366 228868 43398
rect 247868 43954 248868 43986
rect 247868 43718 247930 43954
rect 248166 43718 248250 43954
rect 248486 43718 248570 43954
rect 248806 43718 248868 43954
rect 247868 43634 248868 43718
rect 247868 43398 247930 43634
rect 248166 43398 248250 43634
rect 248486 43398 248570 43634
rect 248806 43398 248868 43634
rect 247868 43366 248868 43398
rect 267868 43954 268868 43986
rect 267868 43718 267930 43954
rect 268166 43718 268250 43954
rect 268486 43718 268570 43954
rect 268806 43718 268868 43954
rect 267868 43634 268868 43718
rect 267868 43398 267930 43634
rect 268166 43398 268250 43634
rect 268486 43398 268570 43634
rect 268806 43398 268868 43634
rect 267868 43366 268868 43398
rect 287868 43954 288868 43986
rect 287868 43718 287930 43954
rect 288166 43718 288250 43954
rect 288486 43718 288570 43954
rect 288806 43718 288868 43954
rect 287868 43634 288868 43718
rect 287868 43398 287930 43634
rect 288166 43398 288250 43634
rect 288486 43398 288570 43634
rect 288806 43398 288868 43634
rect 287868 43366 288868 43398
rect 307868 43954 308868 43986
rect 307868 43718 307930 43954
rect 308166 43718 308250 43954
rect 308486 43718 308570 43954
rect 308806 43718 308868 43954
rect 307868 43634 308868 43718
rect 307868 43398 307930 43634
rect 308166 43398 308250 43634
rect 308486 43398 308570 43634
rect 308806 43398 308868 43634
rect 307868 43366 308868 43398
rect 327868 43954 328868 43986
rect 327868 43718 327930 43954
rect 328166 43718 328250 43954
rect 328486 43718 328570 43954
rect 328806 43718 328868 43954
rect 327868 43634 328868 43718
rect 327868 43398 327930 43634
rect 328166 43398 328250 43634
rect 328486 43398 328570 43634
rect 328806 43398 328868 43634
rect 327868 43366 328868 43398
rect 347868 43954 348868 43986
rect 347868 43718 347930 43954
rect 348166 43718 348250 43954
rect 348486 43718 348570 43954
rect 348806 43718 348868 43954
rect 347868 43634 348868 43718
rect 347868 43398 347930 43634
rect 348166 43398 348250 43634
rect 348486 43398 348570 43634
rect 348806 43398 348868 43634
rect 347868 43366 348868 43398
rect 367868 43954 368868 43986
rect 367868 43718 367930 43954
rect 368166 43718 368250 43954
rect 368486 43718 368570 43954
rect 368806 43718 368868 43954
rect 367868 43634 368868 43718
rect 367868 43398 367930 43634
rect 368166 43398 368250 43634
rect 368486 43398 368570 43634
rect 368806 43398 368868 43634
rect 367868 43366 368868 43398
rect 387868 43954 388868 43986
rect 387868 43718 387930 43954
rect 388166 43718 388250 43954
rect 388486 43718 388570 43954
rect 388806 43718 388868 43954
rect 387868 43634 388868 43718
rect 387868 43398 387930 43634
rect 388166 43398 388250 43634
rect 388486 43398 388570 43634
rect 388806 43398 388868 43634
rect 387868 43366 388868 43398
rect 407868 43954 408868 43986
rect 407868 43718 407930 43954
rect 408166 43718 408250 43954
rect 408486 43718 408570 43954
rect 408806 43718 408868 43954
rect 407868 43634 408868 43718
rect 407868 43398 407930 43634
rect 408166 43398 408250 43634
rect 408486 43398 408570 43634
rect 408806 43398 408868 43634
rect 407868 43366 408868 43398
rect 427868 43954 428868 43986
rect 427868 43718 427930 43954
rect 428166 43718 428250 43954
rect 428486 43718 428570 43954
rect 428806 43718 428868 43954
rect 427868 43634 428868 43718
rect 427868 43398 427930 43634
rect 428166 43398 428250 43634
rect 428486 43398 428570 43634
rect 428806 43398 428868 43634
rect 427868 43366 428868 43398
rect 438294 43954 438914 76000
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 157868 39454 158868 39486
rect 157868 39218 157930 39454
rect 158166 39218 158250 39454
rect 158486 39218 158570 39454
rect 158806 39218 158868 39454
rect 157868 39134 158868 39218
rect 157868 38898 157930 39134
rect 158166 38898 158250 39134
rect 158486 38898 158570 39134
rect 158806 38898 158868 39134
rect 157868 38866 158868 38898
rect 177868 39454 178868 39486
rect 177868 39218 177930 39454
rect 178166 39218 178250 39454
rect 178486 39218 178570 39454
rect 178806 39218 178868 39454
rect 177868 39134 178868 39218
rect 177868 38898 177930 39134
rect 178166 38898 178250 39134
rect 178486 38898 178570 39134
rect 178806 38898 178868 39134
rect 177868 38866 178868 38898
rect 197868 39454 198868 39486
rect 197868 39218 197930 39454
rect 198166 39218 198250 39454
rect 198486 39218 198570 39454
rect 198806 39218 198868 39454
rect 197868 39134 198868 39218
rect 197868 38898 197930 39134
rect 198166 38898 198250 39134
rect 198486 38898 198570 39134
rect 198806 38898 198868 39134
rect 197868 38866 198868 38898
rect 217868 39454 218868 39486
rect 217868 39218 217930 39454
rect 218166 39218 218250 39454
rect 218486 39218 218570 39454
rect 218806 39218 218868 39454
rect 217868 39134 218868 39218
rect 217868 38898 217930 39134
rect 218166 38898 218250 39134
rect 218486 38898 218570 39134
rect 218806 38898 218868 39134
rect 217868 38866 218868 38898
rect 237868 39454 238868 39486
rect 237868 39218 237930 39454
rect 238166 39218 238250 39454
rect 238486 39218 238570 39454
rect 238806 39218 238868 39454
rect 237868 39134 238868 39218
rect 237868 38898 237930 39134
rect 238166 38898 238250 39134
rect 238486 38898 238570 39134
rect 238806 38898 238868 39134
rect 237868 38866 238868 38898
rect 257868 39454 258868 39486
rect 257868 39218 257930 39454
rect 258166 39218 258250 39454
rect 258486 39218 258570 39454
rect 258806 39218 258868 39454
rect 257868 39134 258868 39218
rect 257868 38898 257930 39134
rect 258166 38898 258250 39134
rect 258486 38898 258570 39134
rect 258806 38898 258868 39134
rect 257868 38866 258868 38898
rect 277868 39454 278868 39486
rect 277868 39218 277930 39454
rect 278166 39218 278250 39454
rect 278486 39218 278570 39454
rect 278806 39218 278868 39454
rect 277868 39134 278868 39218
rect 277868 38898 277930 39134
rect 278166 38898 278250 39134
rect 278486 38898 278570 39134
rect 278806 38898 278868 39134
rect 277868 38866 278868 38898
rect 297868 39454 298868 39486
rect 297868 39218 297930 39454
rect 298166 39218 298250 39454
rect 298486 39218 298570 39454
rect 298806 39218 298868 39454
rect 297868 39134 298868 39218
rect 297868 38898 297930 39134
rect 298166 38898 298250 39134
rect 298486 38898 298570 39134
rect 298806 38898 298868 39134
rect 297868 38866 298868 38898
rect 317868 39454 318868 39486
rect 317868 39218 317930 39454
rect 318166 39218 318250 39454
rect 318486 39218 318570 39454
rect 318806 39218 318868 39454
rect 317868 39134 318868 39218
rect 317868 38898 317930 39134
rect 318166 38898 318250 39134
rect 318486 38898 318570 39134
rect 318806 38898 318868 39134
rect 317868 38866 318868 38898
rect 337868 39454 338868 39486
rect 337868 39218 337930 39454
rect 338166 39218 338250 39454
rect 338486 39218 338570 39454
rect 338806 39218 338868 39454
rect 337868 39134 338868 39218
rect 337868 38898 337930 39134
rect 338166 38898 338250 39134
rect 338486 38898 338570 39134
rect 338806 38898 338868 39134
rect 337868 38866 338868 38898
rect 357868 39454 358868 39486
rect 357868 39218 357930 39454
rect 358166 39218 358250 39454
rect 358486 39218 358570 39454
rect 358806 39218 358868 39454
rect 357868 39134 358868 39218
rect 357868 38898 357930 39134
rect 358166 38898 358250 39134
rect 358486 38898 358570 39134
rect 358806 38898 358868 39134
rect 357868 38866 358868 38898
rect 377868 39454 378868 39486
rect 377868 39218 377930 39454
rect 378166 39218 378250 39454
rect 378486 39218 378570 39454
rect 378806 39218 378868 39454
rect 377868 39134 378868 39218
rect 377868 38898 377930 39134
rect 378166 38898 378250 39134
rect 378486 38898 378570 39134
rect 378806 38898 378868 39134
rect 377868 38866 378868 38898
rect 397868 39454 398868 39486
rect 397868 39218 397930 39454
rect 398166 39218 398250 39454
rect 398486 39218 398570 39454
rect 398806 39218 398868 39454
rect 397868 39134 398868 39218
rect 397868 38898 397930 39134
rect 398166 38898 398250 39134
rect 398486 38898 398570 39134
rect 398806 38898 398868 39134
rect 397868 38866 398868 38898
rect 417868 39454 418868 39486
rect 417868 39218 417930 39454
rect 418166 39218 418250 39454
rect 418486 39218 418570 39454
rect 418806 39218 418868 39454
rect 417868 39134 418868 39218
rect 417868 38898 417930 39134
rect 418166 38898 418250 39134
rect 418486 38898 418570 39134
rect 418806 38898 418868 39134
rect 417868 38866 418868 38898
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 22000
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 22000
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 22000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 181794 3454 182414 22000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 7954 186914 22000
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 12454 191414 22000
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 22000
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 22000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 217794 3454 218414 22000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 22000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 22000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 22000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 22000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 253794 3454 254414 22000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 22000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 22000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 22000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 22000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 289794 3454 290414 22000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 22000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 22000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 22000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 22000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 325794 3454 326414 22000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 22000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 22000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 22000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 22000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 361794 3454 362414 22000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 22000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 22000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 22000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 22000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 397794 3454 398414 22000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 22000
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 12454 407414 22000
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 16954 411914 22000
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 21454 416414 22000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 433794 3454 434414 22000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 48454 443414 76000
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 52954 447914 76000
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 57454 452414 76000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 76000
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 66454 461414 76000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 70954 465914 76000
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 75454 470414 76000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 43954 474914 76000
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 48454 479414 76000
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 52954 483914 76000
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 57454 488414 76000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 61954 492914 76000
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 66454 497414 76000
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 70954 501914 76000
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 75454 506414 76000
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 43954 510914 76000
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 48454 515414 76000
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 52954 519914 76000
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 57454 524414 76000
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 61954 528914 76000
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 66454 533414 76000
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 70954 537914 76000
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 75454 542414 76000
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 43954 546914 76000
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 48454 551414 76000
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 52954 555914 76000
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 57454 560414 76000
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 61954 564914 76000
rect 565310 68917 565370 79323
rect 565307 68916 565373 68917
rect 565307 68852 565308 68916
rect 565372 68852 565373 68916
rect 565307 68851 565373 68852
rect 565862 62797 565922 331331
rect 566414 315893 566474 451230
rect 566595 442916 566661 442917
rect 566595 442852 566596 442916
rect 566660 442852 566661 442916
rect 566595 442851 566661 442852
rect 566598 331261 566658 442851
rect 566595 331260 566661 331261
rect 566595 331196 566596 331260
rect 566660 331196 566661 331260
rect 566595 331195 566661 331196
rect 566411 315892 566477 315893
rect 566411 315828 566412 315892
rect 566476 315828 566477 315892
rect 566411 315827 566477 315828
rect 566043 313988 566109 313989
rect 566043 313924 566044 313988
rect 566108 313924 566109 313988
rect 566043 313923 566109 313924
rect 566046 69733 566106 313923
rect 566043 69732 566109 69733
rect 566043 69668 566044 69732
rect 566108 69668 566109 69732
rect 566043 69667 566109 69668
rect 565859 62796 565925 62797
rect 565859 62732 565860 62796
rect 565924 62732 565925 62796
rect 565859 62731 565925 62732
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 566966 54501 567026 585107
rect 567331 580412 567397 580413
rect 567331 580348 567332 580412
rect 567396 580348 567397 580412
rect 567331 580347 567397 580348
rect 567334 459101 567394 580347
rect 570091 580276 570157 580277
rect 570091 580212 570092 580276
rect 570156 580212 570157 580276
rect 570091 580211 570157 580212
rect 568619 571980 568685 571981
rect 568619 571916 568620 571980
rect 568684 571916 568685 571980
rect 568619 571915 568685 571916
rect 568622 461005 568682 571915
rect 568619 461004 568685 461005
rect 568619 460940 568620 461004
rect 568684 460940 568685 461004
rect 568619 460939 568685 460940
rect 570094 460325 570154 580211
rect 570091 460324 570157 460325
rect 570091 460260 570092 460324
rect 570156 460260 570157 460324
rect 570091 460259 570157 460260
rect 570091 460188 570157 460189
rect 570091 460124 570092 460188
rect 570156 460124 570157 460188
rect 570091 460123 570157 460124
rect 570094 459645 570154 460123
rect 570091 459644 570157 459645
rect 570091 459580 570092 459644
rect 570156 459580 570157 459644
rect 570091 459579 570157 459580
rect 567331 459100 567397 459101
rect 567331 459036 567332 459100
rect 567396 459036 567397 459100
rect 567331 459035 567397 459036
rect 567331 458828 567397 458829
rect 567331 458764 567332 458828
rect 567396 458764 567397 458828
rect 567331 458763 567397 458764
rect 567334 76669 567394 458763
rect 568619 458692 568685 458693
rect 568619 458628 568620 458692
rect 568684 458628 568685 458692
rect 568619 458627 568685 458628
rect 568622 314669 568682 458627
rect 569171 418300 569237 418301
rect 569171 418236 569172 418300
rect 569236 418236 569237 418300
rect 569171 418235 569237 418236
rect 568619 314668 568685 314669
rect 568619 314604 568620 314668
rect 568684 314604 568685 314668
rect 568619 314603 568685 314604
rect 569174 188325 569234 418235
rect 570094 334661 570154 459579
rect 570091 334660 570157 334661
rect 570091 334596 570092 334660
rect 570156 334596 570157 334660
rect 570091 334595 570157 334596
rect 570091 331804 570157 331805
rect 570091 331740 570092 331804
rect 570156 331740 570157 331804
rect 570091 331739 570157 331740
rect 570094 200130 570154 331739
rect 570275 201380 570341 201381
rect 570275 201316 570276 201380
rect 570340 201316 570341 201380
rect 570275 201315 570341 201316
rect 569910 200070 570154 200130
rect 569171 188324 569237 188325
rect 569171 188260 569172 188324
rect 569236 188260 569237 188324
rect 569171 188259 569237 188260
rect 568619 187644 568685 187645
rect 568619 187580 568620 187644
rect 568684 187580 568685 187644
rect 568619 187579 568685 187580
rect 568622 77893 568682 187579
rect 568619 77892 568685 77893
rect 568619 77828 568620 77892
rect 568684 77828 568685 77892
rect 568619 77827 568685 77828
rect 567331 76668 567397 76669
rect 567331 76604 567332 76668
rect 567396 76604 567397 76668
rect 567331 76603 567397 76604
rect 569910 76533 569970 200070
rect 570278 180810 570338 201315
rect 570094 180750 570338 180810
rect 569907 76532 569973 76533
rect 569907 76468 569908 76532
rect 569972 76468 569973 76532
rect 569907 76467 569973 76468
rect 568794 66454 569414 76000
rect 570094 71773 570154 180750
rect 571382 76125 571442 585651
rect 573294 574954 573914 610398
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 575243 591020 575309 591021
rect 575243 590956 575244 591020
rect 575308 590956 575309 591020
rect 575243 590955 575309 590956
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 571379 76124 571445 76125
rect 571379 76060 571380 76124
rect 571444 76060 571445 76124
rect 571379 76059 571445 76060
rect 570091 71772 570157 71773
rect 570091 71708 570092 71772
rect 570156 71708 570157 71772
rect 570091 71707 570157 71708
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 566963 54500 567029 54501
rect 566963 54436 566964 54500
rect 567028 54436 567029 54500
rect 566963 54435 567029 54436
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 70954 573914 106398
rect 575246 76533 575306 590955
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 575243 76532 575309 76533
rect 575243 76468 575244 76532
rect 575308 76468 575309 76532
rect 575243 76467 575309 76468
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 33930 691718 34166 691954
rect 34250 691718 34486 691954
rect 34570 691718 34806 691954
rect 33930 691398 34166 691634
rect 34250 691398 34486 691634
rect 34570 691398 34806 691634
rect 53930 691718 54166 691954
rect 54250 691718 54486 691954
rect 54570 691718 54806 691954
rect 53930 691398 54166 691634
rect 54250 691398 54486 691634
rect 54570 691398 54806 691634
rect 73930 691718 74166 691954
rect 74250 691718 74486 691954
rect 74570 691718 74806 691954
rect 73930 691398 74166 691634
rect 74250 691398 74486 691634
rect 74570 691398 74806 691634
rect 93930 691718 94166 691954
rect 94250 691718 94486 691954
rect 94570 691718 94806 691954
rect 93930 691398 94166 691634
rect 94250 691398 94486 691634
rect 94570 691398 94806 691634
rect 113930 691718 114166 691954
rect 114250 691718 114486 691954
rect 114570 691718 114806 691954
rect 113930 691398 114166 691634
rect 114250 691398 114486 691634
rect 114570 691398 114806 691634
rect 133930 691718 134166 691954
rect 134250 691718 134486 691954
rect 134570 691718 134806 691954
rect 133930 691398 134166 691634
rect 134250 691398 134486 691634
rect 134570 691398 134806 691634
rect 153930 691718 154166 691954
rect 154250 691718 154486 691954
rect 154570 691718 154806 691954
rect 153930 691398 154166 691634
rect 154250 691398 154486 691634
rect 154570 691398 154806 691634
rect 173930 691718 174166 691954
rect 174250 691718 174486 691954
rect 174570 691718 174806 691954
rect 173930 691398 174166 691634
rect 174250 691398 174486 691634
rect 174570 691398 174806 691634
rect 193930 691718 194166 691954
rect 194250 691718 194486 691954
rect 194570 691718 194806 691954
rect 193930 691398 194166 691634
rect 194250 691398 194486 691634
rect 194570 691398 194806 691634
rect 213930 691718 214166 691954
rect 214250 691718 214486 691954
rect 214570 691718 214806 691954
rect 213930 691398 214166 691634
rect 214250 691398 214486 691634
rect 214570 691398 214806 691634
rect 233930 691718 234166 691954
rect 234250 691718 234486 691954
rect 234570 691718 234806 691954
rect 233930 691398 234166 691634
rect 234250 691398 234486 691634
rect 234570 691398 234806 691634
rect 253930 691718 254166 691954
rect 254250 691718 254486 691954
rect 254570 691718 254806 691954
rect 253930 691398 254166 691634
rect 254250 691398 254486 691634
rect 254570 691398 254806 691634
rect 273930 691718 274166 691954
rect 274250 691718 274486 691954
rect 274570 691718 274806 691954
rect 273930 691398 274166 691634
rect 274250 691398 274486 691634
rect 274570 691398 274806 691634
rect 23930 687218 24166 687454
rect 24250 687218 24486 687454
rect 24570 687218 24806 687454
rect 23930 686898 24166 687134
rect 24250 686898 24486 687134
rect 24570 686898 24806 687134
rect 43930 687218 44166 687454
rect 44250 687218 44486 687454
rect 44570 687218 44806 687454
rect 43930 686898 44166 687134
rect 44250 686898 44486 687134
rect 44570 686898 44806 687134
rect 63930 687218 64166 687454
rect 64250 687218 64486 687454
rect 64570 687218 64806 687454
rect 63930 686898 64166 687134
rect 64250 686898 64486 687134
rect 64570 686898 64806 687134
rect 83930 687218 84166 687454
rect 84250 687218 84486 687454
rect 84570 687218 84806 687454
rect 83930 686898 84166 687134
rect 84250 686898 84486 687134
rect 84570 686898 84806 687134
rect 103930 687218 104166 687454
rect 104250 687218 104486 687454
rect 104570 687218 104806 687454
rect 103930 686898 104166 687134
rect 104250 686898 104486 687134
rect 104570 686898 104806 687134
rect 123930 687218 124166 687454
rect 124250 687218 124486 687454
rect 124570 687218 124806 687454
rect 123930 686898 124166 687134
rect 124250 686898 124486 687134
rect 124570 686898 124806 687134
rect 143930 687218 144166 687454
rect 144250 687218 144486 687454
rect 144570 687218 144806 687454
rect 143930 686898 144166 687134
rect 144250 686898 144486 687134
rect 144570 686898 144806 687134
rect 163930 687218 164166 687454
rect 164250 687218 164486 687454
rect 164570 687218 164806 687454
rect 163930 686898 164166 687134
rect 164250 686898 164486 687134
rect 164570 686898 164806 687134
rect 183930 687218 184166 687454
rect 184250 687218 184486 687454
rect 184570 687218 184806 687454
rect 183930 686898 184166 687134
rect 184250 686898 184486 687134
rect 184570 686898 184806 687134
rect 203930 687218 204166 687454
rect 204250 687218 204486 687454
rect 204570 687218 204806 687454
rect 203930 686898 204166 687134
rect 204250 686898 204486 687134
rect 204570 686898 204806 687134
rect 223930 687218 224166 687454
rect 224250 687218 224486 687454
rect 224570 687218 224806 687454
rect 223930 686898 224166 687134
rect 224250 686898 224486 687134
rect 224570 686898 224806 687134
rect 243930 687218 244166 687454
rect 244250 687218 244486 687454
rect 244570 687218 244806 687454
rect 243930 686898 244166 687134
rect 244250 686898 244486 687134
rect 244570 686898 244806 687134
rect 263930 687218 264166 687454
rect 264250 687218 264486 687454
rect 264570 687218 264806 687454
rect 263930 686898 264166 687134
rect 264250 686898 264486 687134
rect 264570 686898 264806 687134
rect 283930 687218 284166 687454
rect 284250 687218 284486 687454
rect 284570 687218 284806 687454
rect 283930 686898 284166 687134
rect 284250 686898 284486 687134
rect 284570 686898 284806 687134
rect 33930 655718 34166 655954
rect 34250 655718 34486 655954
rect 34570 655718 34806 655954
rect 33930 655398 34166 655634
rect 34250 655398 34486 655634
rect 34570 655398 34806 655634
rect 53930 655718 54166 655954
rect 54250 655718 54486 655954
rect 54570 655718 54806 655954
rect 53930 655398 54166 655634
rect 54250 655398 54486 655634
rect 54570 655398 54806 655634
rect 73930 655718 74166 655954
rect 74250 655718 74486 655954
rect 74570 655718 74806 655954
rect 73930 655398 74166 655634
rect 74250 655398 74486 655634
rect 74570 655398 74806 655634
rect 93930 655718 94166 655954
rect 94250 655718 94486 655954
rect 94570 655718 94806 655954
rect 93930 655398 94166 655634
rect 94250 655398 94486 655634
rect 94570 655398 94806 655634
rect 113930 655718 114166 655954
rect 114250 655718 114486 655954
rect 114570 655718 114806 655954
rect 113930 655398 114166 655634
rect 114250 655398 114486 655634
rect 114570 655398 114806 655634
rect 133930 655718 134166 655954
rect 134250 655718 134486 655954
rect 134570 655718 134806 655954
rect 133930 655398 134166 655634
rect 134250 655398 134486 655634
rect 134570 655398 134806 655634
rect 153930 655718 154166 655954
rect 154250 655718 154486 655954
rect 154570 655718 154806 655954
rect 153930 655398 154166 655634
rect 154250 655398 154486 655634
rect 154570 655398 154806 655634
rect 173930 655718 174166 655954
rect 174250 655718 174486 655954
rect 174570 655718 174806 655954
rect 173930 655398 174166 655634
rect 174250 655398 174486 655634
rect 174570 655398 174806 655634
rect 193930 655718 194166 655954
rect 194250 655718 194486 655954
rect 194570 655718 194806 655954
rect 193930 655398 194166 655634
rect 194250 655398 194486 655634
rect 194570 655398 194806 655634
rect 213930 655718 214166 655954
rect 214250 655718 214486 655954
rect 214570 655718 214806 655954
rect 213930 655398 214166 655634
rect 214250 655398 214486 655634
rect 214570 655398 214806 655634
rect 233930 655718 234166 655954
rect 234250 655718 234486 655954
rect 234570 655718 234806 655954
rect 233930 655398 234166 655634
rect 234250 655398 234486 655634
rect 234570 655398 234806 655634
rect 253930 655718 254166 655954
rect 254250 655718 254486 655954
rect 254570 655718 254806 655954
rect 253930 655398 254166 655634
rect 254250 655398 254486 655634
rect 254570 655398 254806 655634
rect 273930 655718 274166 655954
rect 274250 655718 274486 655954
rect 274570 655718 274806 655954
rect 273930 655398 274166 655634
rect 274250 655398 274486 655634
rect 274570 655398 274806 655634
rect 23930 651218 24166 651454
rect 24250 651218 24486 651454
rect 24570 651218 24806 651454
rect 23930 650898 24166 651134
rect 24250 650898 24486 651134
rect 24570 650898 24806 651134
rect 43930 651218 44166 651454
rect 44250 651218 44486 651454
rect 44570 651218 44806 651454
rect 43930 650898 44166 651134
rect 44250 650898 44486 651134
rect 44570 650898 44806 651134
rect 63930 651218 64166 651454
rect 64250 651218 64486 651454
rect 64570 651218 64806 651454
rect 63930 650898 64166 651134
rect 64250 650898 64486 651134
rect 64570 650898 64806 651134
rect 83930 651218 84166 651454
rect 84250 651218 84486 651454
rect 84570 651218 84806 651454
rect 83930 650898 84166 651134
rect 84250 650898 84486 651134
rect 84570 650898 84806 651134
rect 103930 651218 104166 651454
rect 104250 651218 104486 651454
rect 104570 651218 104806 651454
rect 103930 650898 104166 651134
rect 104250 650898 104486 651134
rect 104570 650898 104806 651134
rect 123930 651218 124166 651454
rect 124250 651218 124486 651454
rect 124570 651218 124806 651454
rect 123930 650898 124166 651134
rect 124250 650898 124486 651134
rect 124570 650898 124806 651134
rect 143930 651218 144166 651454
rect 144250 651218 144486 651454
rect 144570 651218 144806 651454
rect 143930 650898 144166 651134
rect 144250 650898 144486 651134
rect 144570 650898 144806 651134
rect 163930 651218 164166 651454
rect 164250 651218 164486 651454
rect 164570 651218 164806 651454
rect 163930 650898 164166 651134
rect 164250 650898 164486 651134
rect 164570 650898 164806 651134
rect 183930 651218 184166 651454
rect 184250 651218 184486 651454
rect 184570 651218 184806 651454
rect 183930 650898 184166 651134
rect 184250 650898 184486 651134
rect 184570 650898 184806 651134
rect 203930 651218 204166 651454
rect 204250 651218 204486 651454
rect 204570 651218 204806 651454
rect 203930 650898 204166 651134
rect 204250 650898 204486 651134
rect 204570 650898 204806 651134
rect 223930 651218 224166 651454
rect 224250 651218 224486 651454
rect 224570 651218 224806 651454
rect 223930 650898 224166 651134
rect 224250 650898 224486 651134
rect 224570 650898 224806 651134
rect 243930 651218 244166 651454
rect 244250 651218 244486 651454
rect 244570 651218 244806 651454
rect 243930 650898 244166 651134
rect 244250 650898 244486 651134
rect 244570 650898 244806 651134
rect 263930 651218 264166 651454
rect 264250 651218 264486 651454
rect 264570 651218 264806 651454
rect 263930 650898 264166 651134
rect 264250 650898 264486 651134
rect 264570 650898 264806 651134
rect 283930 651218 284166 651454
rect 284250 651218 284486 651454
rect 284570 651218 284806 651454
rect 283930 650898 284166 651134
rect 284250 650898 284486 651134
rect 284570 650898 284806 651134
rect 33930 619718 34166 619954
rect 34250 619718 34486 619954
rect 34570 619718 34806 619954
rect 33930 619398 34166 619634
rect 34250 619398 34486 619634
rect 34570 619398 34806 619634
rect 53930 619718 54166 619954
rect 54250 619718 54486 619954
rect 54570 619718 54806 619954
rect 53930 619398 54166 619634
rect 54250 619398 54486 619634
rect 54570 619398 54806 619634
rect 73930 619718 74166 619954
rect 74250 619718 74486 619954
rect 74570 619718 74806 619954
rect 73930 619398 74166 619634
rect 74250 619398 74486 619634
rect 74570 619398 74806 619634
rect 93930 619718 94166 619954
rect 94250 619718 94486 619954
rect 94570 619718 94806 619954
rect 93930 619398 94166 619634
rect 94250 619398 94486 619634
rect 94570 619398 94806 619634
rect 113930 619718 114166 619954
rect 114250 619718 114486 619954
rect 114570 619718 114806 619954
rect 113930 619398 114166 619634
rect 114250 619398 114486 619634
rect 114570 619398 114806 619634
rect 133930 619718 134166 619954
rect 134250 619718 134486 619954
rect 134570 619718 134806 619954
rect 133930 619398 134166 619634
rect 134250 619398 134486 619634
rect 134570 619398 134806 619634
rect 153930 619718 154166 619954
rect 154250 619718 154486 619954
rect 154570 619718 154806 619954
rect 153930 619398 154166 619634
rect 154250 619398 154486 619634
rect 154570 619398 154806 619634
rect 173930 619718 174166 619954
rect 174250 619718 174486 619954
rect 174570 619718 174806 619954
rect 173930 619398 174166 619634
rect 174250 619398 174486 619634
rect 174570 619398 174806 619634
rect 193930 619718 194166 619954
rect 194250 619718 194486 619954
rect 194570 619718 194806 619954
rect 193930 619398 194166 619634
rect 194250 619398 194486 619634
rect 194570 619398 194806 619634
rect 213930 619718 214166 619954
rect 214250 619718 214486 619954
rect 214570 619718 214806 619954
rect 213930 619398 214166 619634
rect 214250 619398 214486 619634
rect 214570 619398 214806 619634
rect 233930 619718 234166 619954
rect 234250 619718 234486 619954
rect 234570 619718 234806 619954
rect 233930 619398 234166 619634
rect 234250 619398 234486 619634
rect 234570 619398 234806 619634
rect 253930 619718 254166 619954
rect 254250 619718 254486 619954
rect 254570 619718 254806 619954
rect 253930 619398 254166 619634
rect 254250 619398 254486 619634
rect 254570 619398 254806 619634
rect 273930 619718 274166 619954
rect 274250 619718 274486 619954
rect 274570 619718 274806 619954
rect 273930 619398 274166 619634
rect 274250 619398 274486 619634
rect 274570 619398 274806 619634
rect 23930 615218 24166 615454
rect 24250 615218 24486 615454
rect 24570 615218 24806 615454
rect 23930 614898 24166 615134
rect 24250 614898 24486 615134
rect 24570 614898 24806 615134
rect 43930 615218 44166 615454
rect 44250 615218 44486 615454
rect 44570 615218 44806 615454
rect 43930 614898 44166 615134
rect 44250 614898 44486 615134
rect 44570 614898 44806 615134
rect 63930 615218 64166 615454
rect 64250 615218 64486 615454
rect 64570 615218 64806 615454
rect 63930 614898 64166 615134
rect 64250 614898 64486 615134
rect 64570 614898 64806 615134
rect 83930 615218 84166 615454
rect 84250 615218 84486 615454
rect 84570 615218 84806 615454
rect 83930 614898 84166 615134
rect 84250 614898 84486 615134
rect 84570 614898 84806 615134
rect 103930 615218 104166 615454
rect 104250 615218 104486 615454
rect 104570 615218 104806 615454
rect 103930 614898 104166 615134
rect 104250 614898 104486 615134
rect 104570 614898 104806 615134
rect 123930 615218 124166 615454
rect 124250 615218 124486 615454
rect 124570 615218 124806 615454
rect 123930 614898 124166 615134
rect 124250 614898 124486 615134
rect 124570 614898 124806 615134
rect 143930 615218 144166 615454
rect 144250 615218 144486 615454
rect 144570 615218 144806 615454
rect 143930 614898 144166 615134
rect 144250 614898 144486 615134
rect 144570 614898 144806 615134
rect 163930 615218 164166 615454
rect 164250 615218 164486 615454
rect 164570 615218 164806 615454
rect 163930 614898 164166 615134
rect 164250 614898 164486 615134
rect 164570 614898 164806 615134
rect 183930 615218 184166 615454
rect 184250 615218 184486 615454
rect 184570 615218 184806 615454
rect 183930 614898 184166 615134
rect 184250 614898 184486 615134
rect 184570 614898 184806 615134
rect 203930 615218 204166 615454
rect 204250 615218 204486 615454
rect 204570 615218 204806 615454
rect 203930 614898 204166 615134
rect 204250 614898 204486 615134
rect 204570 614898 204806 615134
rect 223930 615218 224166 615454
rect 224250 615218 224486 615454
rect 224570 615218 224806 615454
rect 223930 614898 224166 615134
rect 224250 614898 224486 615134
rect 224570 614898 224806 615134
rect 243930 615218 244166 615454
rect 244250 615218 244486 615454
rect 244570 615218 244806 615454
rect 243930 614898 244166 615134
rect 244250 614898 244486 615134
rect 244570 614898 244806 615134
rect 263930 615218 264166 615454
rect 264250 615218 264486 615454
rect 264570 615218 264806 615454
rect 263930 614898 264166 615134
rect 264250 614898 264486 615134
rect 264570 614898 264806 615134
rect 283930 615218 284166 615454
rect 284250 615218 284486 615454
rect 284570 615218 284806 615454
rect 283930 614898 284166 615134
rect 284250 614898 284486 615134
rect 284570 614898 284806 615134
rect 33930 547718 34166 547954
rect 34250 547718 34486 547954
rect 34570 547718 34806 547954
rect 33930 547398 34166 547634
rect 34250 547398 34486 547634
rect 34570 547398 34806 547634
rect 53930 547718 54166 547954
rect 54250 547718 54486 547954
rect 54570 547718 54806 547954
rect 53930 547398 54166 547634
rect 54250 547398 54486 547634
rect 54570 547398 54806 547634
rect 73930 547718 74166 547954
rect 74250 547718 74486 547954
rect 74570 547718 74806 547954
rect 73930 547398 74166 547634
rect 74250 547398 74486 547634
rect 74570 547398 74806 547634
rect 93930 547718 94166 547954
rect 94250 547718 94486 547954
rect 94570 547718 94806 547954
rect 93930 547398 94166 547634
rect 94250 547398 94486 547634
rect 94570 547398 94806 547634
rect 113930 547718 114166 547954
rect 114250 547718 114486 547954
rect 114570 547718 114806 547954
rect 113930 547398 114166 547634
rect 114250 547398 114486 547634
rect 114570 547398 114806 547634
rect 133930 547718 134166 547954
rect 134250 547718 134486 547954
rect 134570 547718 134806 547954
rect 133930 547398 134166 547634
rect 134250 547398 134486 547634
rect 134570 547398 134806 547634
rect 153930 547718 154166 547954
rect 154250 547718 154486 547954
rect 154570 547718 154806 547954
rect 153930 547398 154166 547634
rect 154250 547398 154486 547634
rect 154570 547398 154806 547634
rect 173930 547718 174166 547954
rect 174250 547718 174486 547954
rect 174570 547718 174806 547954
rect 173930 547398 174166 547634
rect 174250 547398 174486 547634
rect 174570 547398 174806 547634
rect 193930 547718 194166 547954
rect 194250 547718 194486 547954
rect 194570 547718 194806 547954
rect 193930 547398 194166 547634
rect 194250 547398 194486 547634
rect 194570 547398 194806 547634
rect 213930 547718 214166 547954
rect 214250 547718 214486 547954
rect 214570 547718 214806 547954
rect 213930 547398 214166 547634
rect 214250 547398 214486 547634
rect 214570 547398 214806 547634
rect 233930 547718 234166 547954
rect 234250 547718 234486 547954
rect 234570 547718 234806 547954
rect 233930 547398 234166 547634
rect 234250 547398 234486 547634
rect 234570 547398 234806 547634
rect 253930 547718 254166 547954
rect 254250 547718 254486 547954
rect 254570 547718 254806 547954
rect 253930 547398 254166 547634
rect 254250 547398 254486 547634
rect 254570 547398 254806 547634
rect 273930 547718 274166 547954
rect 274250 547718 274486 547954
rect 274570 547718 274806 547954
rect 273930 547398 274166 547634
rect 274250 547398 274486 547634
rect 274570 547398 274806 547634
rect 23930 543218 24166 543454
rect 24250 543218 24486 543454
rect 24570 543218 24806 543454
rect 23930 542898 24166 543134
rect 24250 542898 24486 543134
rect 24570 542898 24806 543134
rect 43930 543218 44166 543454
rect 44250 543218 44486 543454
rect 44570 543218 44806 543454
rect 43930 542898 44166 543134
rect 44250 542898 44486 543134
rect 44570 542898 44806 543134
rect 63930 543218 64166 543454
rect 64250 543218 64486 543454
rect 64570 543218 64806 543454
rect 63930 542898 64166 543134
rect 64250 542898 64486 543134
rect 64570 542898 64806 543134
rect 83930 543218 84166 543454
rect 84250 543218 84486 543454
rect 84570 543218 84806 543454
rect 83930 542898 84166 543134
rect 84250 542898 84486 543134
rect 84570 542898 84806 543134
rect 103930 543218 104166 543454
rect 104250 543218 104486 543454
rect 104570 543218 104806 543454
rect 103930 542898 104166 543134
rect 104250 542898 104486 543134
rect 104570 542898 104806 543134
rect 123930 543218 124166 543454
rect 124250 543218 124486 543454
rect 124570 543218 124806 543454
rect 123930 542898 124166 543134
rect 124250 542898 124486 543134
rect 124570 542898 124806 543134
rect 143930 543218 144166 543454
rect 144250 543218 144486 543454
rect 144570 543218 144806 543454
rect 143930 542898 144166 543134
rect 144250 542898 144486 543134
rect 144570 542898 144806 543134
rect 163930 543218 164166 543454
rect 164250 543218 164486 543454
rect 164570 543218 164806 543454
rect 163930 542898 164166 543134
rect 164250 542898 164486 543134
rect 164570 542898 164806 543134
rect 183930 543218 184166 543454
rect 184250 543218 184486 543454
rect 184570 543218 184806 543454
rect 183930 542898 184166 543134
rect 184250 542898 184486 543134
rect 184570 542898 184806 543134
rect 203930 543218 204166 543454
rect 204250 543218 204486 543454
rect 204570 543218 204806 543454
rect 203930 542898 204166 543134
rect 204250 542898 204486 543134
rect 204570 542898 204806 543134
rect 223930 543218 224166 543454
rect 224250 543218 224486 543454
rect 224570 543218 224806 543454
rect 223930 542898 224166 543134
rect 224250 542898 224486 543134
rect 224570 542898 224806 543134
rect 243930 543218 244166 543454
rect 244250 543218 244486 543454
rect 244570 543218 244806 543454
rect 243930 542898 244166 543134
rect 244250 542898 244486 543134
rect 244570 542898 244806 543134
rect 263930 543218 264166 543454
rect 264250 543218 264486 543454
rect 264570 543218 264806 543454
rect 263930 542898 264166 543134
rect 264250 542898 264486 543134
rect 264570 542898 264806 543134
rect 283930 543218 284166 543454
rect 284250 543218 284486 543454
rect 284570 543218 284806 543454
rect 283930 542898 284166 543134
rect 284250 542898 284486 543134
rect 284570 542898 284806 543134
rect 33930 511718 34166 511954
rect 34250 511718 34486 511954
rect 34570 511718 34806 511954
rect 33930 511398 34166 511634
rect 34250 511398 34486 511634
rect 34570 511398 34806 511634
rect 53930 511718 54166 511954
rect 54250 511718 54486 511954
rect 54570 511718 54806 511954
rect 53930 511398 54166 511634
rect 54250 511398 54486 511634
rect 54570 511398 54806 511634
rect 73930 511718 74166 511954
rect 74250 511718 74486 511954
rect 74570 511718 74806 511954
rect 73930 511398 74166 511634
rect 74250 511398 74486 511634
rect 74570 511398 74806 511634
rect 93930 511718 94166 511954
rect 94250 511718 94486 511954
rect 94570 511718 94806 511954
rect 93930 511398 94166 511634
rect 94250 511398 94486 511634
rect 94570 511398 94806 511634
rect 113930 511718 114166 511954
rect 114250 511718 114486 511954
rect 114570 511718 114806 511954
rect 113930 511398 114166 511634
rect 114250 511398 114486 511634
rect 114570 511398 114806 511634
rect 133930 511718 134166 511954
rect 134250 511718 134486 511954
rect 134570 511718 134806 511954
rect 133930 511398 134166 511634
rect 134250 511398 134486 511634
rect 134570 511398 134806 511634
rect 153930 511718 154166 511954
rect 154250 511718 154486 511954
rect 154570 511718 154806 511954
rect 153930 511398 154166 511634
rect 154250 511398 154486 511634
rect 154570 511398 154806 511634
rect 173930 511718 174166 511954
rect 174250 511718 174486 511954
rect 174570 511718 174806 511954
rect 173930 511398 174166 511634
rect 174250 511398 174486 511634
rect 174570 511398 174806 511634
rect 193930 511718 194166 511954
rect 194250 511718 194486 511954
rect 194570 511718 194806 511954
rect 193930 511398 194166 511634
rect 194250 511398 194486 511634
rect 194570 511398 194806 511634
rect 213930 511718 214166 511954
rect 214250 511718 214486 511954
rect 214570 511718 214806 511954
rect 213930 511398 214166 511634
rect 214250 511398 214486 511634
rect 214570 511398 214806 511634
rect 233930 511718 234166 511954
rect 234250 511718 234486 511954
rect 234570 511718 234806 511954
rect 233930 511398 234166 511634
rect 234250 511398 234486 511634
rect 234570 511398 234806 511634
rect 253930 511718 254166 511954
rect 254250 511718 254486 511954
rect 254570 511718 254806 511954
rect 253930 511398 254166 511634
rect 254250 511398 254486 511634
rect 254570 511398 254806 511634
rect 273930 511718 274166 511954
rect 274250 511718 274486 511954
rect 274570 511718 274806 511954
rect 273930 511398 274166 511634
rect 274250 511398 274486 511634
rect 274570 511398 274806 511634
rect 23930 507218 24166 507454
rect 24250 507218 24486 507454
rect 24570 507218 24806 507454
rect 23930 506898 24166 507134
rect 24250 506898 24486 507134
rect 24570 506898 24806 507134
rect 43930 507218 44166 507454
rect 44250 507218 44486 507454
rect 44570 507218 44806 507454
rect 43930 506898 44166 507134
rect 44250 506898 44486 507134
rect 44570 506898 44806 507134
rect 63930 507218 64166 507454
rect 64250 507218 64486 507454
rect 64570 507218 64806 507454
rect 63930 506898 64166 507134
rect 64250 506898 64486 507134
rect 64570 506898 64806 507134
rect 83930 507218 84166 507454
rect 84250 507218 84486 507454
rect 84570 507218 84806 507454
rect 83930 506898 84166 507134
rect 84250 506898 84486 507134
rect 84570 506898 84806 507134
rect 103930 507218 104166 507454
rect 104250 507218 104486 507454
rect 104570 507218 104806 507454
rect 103930 506898 104166 507134
rect 104250 506898 104486 507134
rect 104570 506898 104806 507134
rect 123930 507218 124166 507454
rect 124250 507218 124486 507454
rect 124570 507218 124806 507454
rect 123930 506898 124166 507134
rect 124250 506898 124486 507134
rect 124570 506898 124806 507134
rect 143930 507218 144166 507454
rect 144250 507218 144486 507454
rect 144570 507218 144806 507454
rect 143930 506898 144166 507134
rect 144250 506898 144486 507134
rect 144570 506898 144806 507134
rect 163930 507218 164166 507454
rect 164250 507218 164486 507454
rect 164570 507218 164806 507454
rect 163930 506898 164166 507134
rect 164250 506898 164486 507134
rect 164570 506898 164806 507134
rect 183930 507218 184166 507454
rect 184250 507218 184486 507454
rect 184570 507218 184806 507454
rect 183930 506898 184166 507134
rect 184250 506898 184486 507134
rect 184570 506898 184806 507134
rect 203930 507218 204166 507454
rect 204250 507218 204486 507454
rect 204570 507218 204806 507454
rect 203930 506898 204166 507134
rect 204250 506898 204486 507134
rect 204570 506898 204806 507134
rect 223930 507218 224166 507454
rect 224250 507218 224486 507454
rect 224570 507218 224806 507454
rect 223930 506898 224166 507134
rect 224250 506898 224486 507134
rect 224570 506898 224806 507134
rect 243930 507218 244166 507454
rect 244250 507218 244486 507454
rect 244570 507218 244806 507454
rect 243930 506898 244166 507134
rect 244250 506898 244486 507134
rect 244570 506898 244806 507134
rect 263930 507218 264166 507454
rect 264250 507218 264486 507454
rect 264570 507218 264806 507454
rect 263930 506898 264166 507134
rect 264250 506898 264486 507134
rect 264570 506898 264806 507134
rect 283930 507218 284166 507454
rect 284250 507218 284486 507454
rect 284570 507218 284806 507454
rect 283930 506898 284166 507134
rect 284250 506898 284486 507134
rect 284570 506898 284806 507134
rect 33930 475718 34166 475954
rect 34250 475718 34486 475954
rect 34570 475718 34806 475954
rect 33930 475398 34166 475634
rect 34250 475398 34486 475634
rect 34570 475398 34806 475634
rect 53930 475718 54166 475954
rect 54250 475718 54486 475954
rect 54570 475718 54806 475954
rect 53930 475398 54166 475634
rect 54250 475398 54486 475634
rect 54570 475398 54806 475634
rect 73930 475718 74166 475954
rect 74250 475718 74486 475954
rect 74570 475718 74806 475954
rect 73930 475398 74166 475634
rect 74250 475398 74486 475634
rect 74570 475398 74806 475634
rect 93930 475718 94166 475954
rect 94250 475718 94486 475954
rect 94570 475718 94806 475954
rect 93930 475398 94166 475634
rect 94250 475398 94486 475634
rect 94570 475398 94806 475634
rect 113930 475718 114166 475954
rect 114250 475718 114486 475954
rect 114570 475718 114806 475954
rect 113930 475398 114166 475634
rect 114250 475398 114486 475634
rect 114570 475398 114806 475634
rect 133930 475718 134166 475954
rect 134250 475718 134486 475954
rect 134570 475718 134806 475954
rect 133930 475398 134166 475634
rect 134250 475398 134486 475634
rect 134570 475398 134806 475634
rect 153930 475718 154166 475954
rect 154250 475718 154486 475954
rect 154570 475718 154806 475954
rect 153930 475398 154166 475634
rect 154250 475398 154486 475634
rect 154570 475398 154806 475634
rect 173930 475718 174166 475954
rect 174250 475718 174486 475954
rect 174570 475718 174806 475954
rect 173930 475398 174166 475634
rect 174250 475398 174486 475634
rect 174570 475398 174806 475634
rect 193930 475718 194166 475954
rect 194250 475718 194486 475954
rect 194570 475718 194806 475954
rect 193930 475398 194166 475634
rect 194250 475398 194486 475634
rect 194570 475398 194806 475634
rect 213930 475718 214166 475954
rect 214250 475718 214486 475954
rect 214570 475718 214806 475954
rect 213930 475398 214166 475634
rect 214250 475398 214486 475634
rect 214570 475398 214806 475634
rect 233930 475718 234166 475954
rect 234250 475718 234486 475954
rect 234570 475718 234806 475954
rect 233930 475398 234166 475634
rect 234250 475398 234486 475634
rect 234570 475398 234806 475634
rect 253930 475718 254166 475954
rect 254250 475718 254486 475954
rect 254570 475718 254806 475954
rect 253930 475398 254166 475634
rect 254250 475398 254486 475634
rect 254570 475398 254806 475634
rect 273930 475718 274166 475954
rect 274250 475718 274486 475954
rect 274570 475718 274806 475954
rect 273930 475398 274166 475634
rect 274250 475398 274486 475634
rect 274570 475398 274806 475634
rect 23930 471218 24166 471454
rect 24250 471218 24486 471454
rect 24570 471218 24806 471454
rect 23930 470898 24166 471134
rect 24250 470898 24486 471134
rect 24570 470898 24806 471134
rect 43930 471218 44166 471454
rect 44250 471218 44486 471454
rect 44570 471218 44806 471454
rect 43930 470898 44166 471134
rect 44250 470898 44486 471134
rect 44570 470898 44806 471134
rect 63930 471218 64166 471454
rect 64250 471218 64486 471454
rect 64570 471218 64806 471454
rect 63930 470898 64166 471134
rect 64250 470898 64486 471134
rect 64570 470898 64806 471134
rect 83930 471218 84166 471454
rect 84250 471218 84486 471454
rect 84570 471218 84806 471454
rect 83930 470898 84166 471134
rect 84250 470898 84486 471134
rect 84570 470898 84806 471134
rect 103930 471218 104166 471454
rect 104250 471218 104486 471454
rect 104570 471218 104806 471454
rect 103930 470898 104166 471134
rect 104250 470898 104486 471134
rect 104570 470898 104806 471134
rect 123930 471218 124166 471454
rect 124250 471218 124486 471454
rect 124570 471218 124806 471454
rect 123930 470898 124166 471134
rect 124250 470898 124486 471134
rect 124570 470898 124806 471134
rect 143930 471218 144166 471454
rect 144250 471218 144486 471454
rect 144570 471218 144806 471454
rect 143930 470898 144166 471134
rect 144250 470898 144486 471134
rect 144570 470898 144806 471134
rect 163930 471218 164166 471454
rect 164250 471218 164486 471454
rect 164570 471218 164806 471454
rect 163930 470898 164166 471134
rect 164250 470898 164486 471134
rect 164570 470898 164806 471134
rect 183930 471218 184166 471454
rect 184250 471218 184486 471454
rect 184570 471218 184806 471454
rect 183930 470898 184166 471134
rect 184250 470898 184486 471134
rect 184570 470898 184806 471134
rect 203930 471218 204166 471454
rect 204250 471218 204486 471454
rect 204570 471218 204806 471454
rect 203930 470898 204166 471134
rect 204250 470898 204486 471134
rect 204570 470898 204806 471134
rect 223930 471218 224166 471454
rect 224250 471218 224486 471454
rect 224570 471218 224806 471454
rect 223930 470898 224166 471134
rect 224250 470898 224486 471134
rect 224570 470898 224806 471134
rect 243930 471218 244166 471454
rect 244250 471218 244486 471454
rect 244570 471218 244806 471454
rect 243930 470898 244166 471134
rect 244250 470898 244486 471134
rect 244570 470898 244806 471134
rect 263930 471218 264166 471454
rect 264250 471218 264486 471454
rect 264570 471218 264806 471454
rect 263930 470898 264166 471134
rect 264250 470898 264486 471134
rect 264570 470898 264806 471134
rect 283930 471218 284166 471454
rect 284250 471218 284486 471454
rect 284570 471218 284806 471454
rect 283930 470898 284166 471134
rect 284250 470898 284486 471134
rect 284570 470898 284806 471134
rect 33930 439718 34166 439954
rect 34250 439718 34486 439954
rect 34570 439718 34806 439954
rect 33930 439398 34166 439634
rect 34250 439398 34486 439634
rect 34570 439398 34806 439634
rect 53930 439718 54166 439954
rect 54250 439718 54486 439954
rect 54570 439718 54806 439954
rect 53930 439398 54166 439634
rect 54250 439398 54486 439634
rect 54570 439398 54806 439634
rect 73930 439718 74166 439954
rect 74250 439718 74486 439954
rect 74570 439718 74806 439954
rect 73930 439398 74166 439634
rect 74250 439398 74486 439634
rect 74570 439398 74806 439634
rect 93930 439718 94166 439954
rect 94250 439718 94486 439954
rect 94570 439718 94806 439954
rect 93930 439398 94166 439634
rect 94250 439398 94486 439634
rect 94570 439398 94806 439634
rect 113930 439718 114166 439954
rect 114250 439718 114486 439954
rect 114570 439718 114806 439954
rect 113930 439398 114166 439634
rect 114250 439398 114486 439634
rect 114570 439398 114806 439634
rect 133930 439718 134166 439954
rect 134250 439718 134486 439954
rect 134570 439718 134806 439954
rect 133930 439398 134166 439634
rect 134250 439398 134486 439634
rect 134570 439398 134806 439634
rect 153930 439718 154166 439954
rect 154250 439718 154486 439954
rect 154570 439718 154806 439954
rect 153930 439398 154166 439634
rect 154250 439398 154486 439634
rect 154570 439398 154806 439634
rect 173930 439718 174166 439954
rect 174250 439718 174486 439954
rect 174570 439718 174806 439954
rect 173930 439398 174166 439634
rect 174250 439398 174486 439634
rect 174570 439398 174806 439634
rect 193930 439718 194166 439954
rect 194250 439718 194486 439954
rect 194570 439718 194806 439954
rect 193930 439398 194166 439634
rect 194250 439398 194486 439634
rect 194570 439398 194806 439634
rect 213930 439718 214166 439954
rect 214250 439718 214486 439954
rect 214570 439718 214806 439954
rect 213930 439398 214166 439634
rect 214250 439398 214486 439634
rect 214570 439398 214806 439634
rect 233930 439718 234166 439954
rect 234250 439718 234486 439954
rect 234570 439718 234806 439954
rect 233930 439398 234166 439634
rect 234250 439398 234486 439634
rect 234570 439398 234806 439634
rect 253930 439718 254166 439954
rect 254250 439718 254486 439954
rect 254570 439718 254806 439954
rect 253930 439398 254166 439634
rect 254250 439398 254486 439634
rect 254570 439398 254806 439634
rect 273930 439718 274166 439954
rect 274250 439718 274486 439954
rect 274570 439718 274806 439954
rect 273930 439398 274166 439634
rect 274250 439398 274486 439634
rect 274570 439398 274806 439634
rect 23930 435218 24166 435454
rect 24250 435218 24486 435454
rect 24570 435218 24806 435454
rect 23930 434898 24166 435134
rect 24250 434898 24486 435134
rect 24570 434898 24806 435134
rect 43930 435218 44166 435454
rect 44250 435218 44486 435454
rect 44570 435218 44806 435454
rect 43930 434898 44166 435134
rect 44250 434898 44486 435134
rect 44570 434898 44806 435134
rect 63930 435218 64166 435454
rect 64250 435218 64486 435454
rect 64570 435218 64806 435454
rect 63930 434898 64166 435134
rect 64250 434898 64486 435134
rect 64570 434898 64806 435134
rect 83930 435218 84166 435454
rect 84250 435218 84486 435454
rect 84570 435218 84806 435454
rect 83930 434898 84166 435134
rect 84250 434898 84486 435134
rect 84570 434898 84806 435134
rect 103930 435218 104166 435454
rect 104250 435218 104486 435454
rect 104570 435218 104806 435454
rect 103930 434898 104166 435134
rect 104250 434898 104486 435134
rect 104570 434898 104806 435134
rect 123930 435218 124166 435454
rect 124250 435218 124486 435454
rect 124570 435218 124806 435454
rect 123930 434898 124166 435134
rect 124250 434898 124486 435134
rect 124570 434898 124806 435134
rect 143930 435218 144166 435454
rect 144250 435218 144486 435454
rect 144570 435218 144806 435454
rect 143930 434898 144166 435134
rect 144250 434898 144486 435134
rect 144570 434898 144806 435134
rect 163930 435218 164166 435454
rect 164250 435218 164486 435454
rect 164570 435218 164806 435454
rect 163930 434898 164166 435134
rect 164250 434898 164486 435134
rect 164570 434898 164806 435134
rect 183930 435218 184166 435454
rect 184250 435218 184486 435454
rect 184570 435218 184806 435454
rect 183930 434898 184166 435134
rect 184250 434898 184486 435134
rect 184570 434898 184806 435134
rect 203930 435218 204166 435454
rect 204250 435218 204486 435454
rect 204570 435218 204806 435454
rect 203930 434898 204166 435134
rect 204250 434898 204486 435134
rect 204570 434898 204806 435134
rect 223930 435218 224166 435454
rect 224250 435218 224486 435454
rect 224570 435218 224806 435454
rect 223930 434898 224166 435134
rect 224250 434898 224486 435134
rect 224570 434898 224806 435134
rect 243930 435218 244166 435454
rect 244250 435218 244486 435454
rect 244570 435218 244806 435454
rect 243930 434898 244166 435134
rect 244250 434898 244486 435134
rect 244570 434898 244806 435134
rect 263930 435218 264166 435454
rect 264250 435218 264486 435454
rect 264570 435218 264806 435454
rect 263930 434898 264166 435134
rect 264250 434898 264486 435134
rect 264570 434898 264806 435134
rect 283930 435218 284166 435454
rect 284250 435218 284486 435454
rect 284570 435218 284806 435454
rect 283930 434898 284166 435134
rect 284250 434898 284486 435134
rect 284570 434898 284806 435134
rect 33930 403718 34166 403954
rect 34250 403718 34486 403954
rect 34570 403718 34806 403954
rect 33930 403398 34166 403634
rect 34250 403398 34486 403634
rect 34570 403398 34806 403634
rect 53930 403718 54166 403954
rect 54250 403718 54486 403954
rect 54570 403718 54806 403954
rect 53930 403398 54166 403634
rect 54250 403398 54486 403634
rect 54570 403398 54806 403634
rect 73930 403718 74166 403954
rect 74250 403718 74486 403954
rect 74570 403718 74806 403954
rect 73930 403398 74166 403634
rect 74250 403398 74486 403634
rect 74570 403398 74806 403634
rect 93930 403718 94166 403954
rect 94250 403718 94486 403954
rect 94570 403718 94806 403954
rect 93930 403398 94166 403634
rect 94250 403398 94486 403634
rect 94570 403398 94806 403634
rect 113930 403718 114166 403954
rect 114250 403718 114486 403954
rect 114570 403718 114806 403954
rect 113930 403398 114166 403634
rect 114250 403398 114486 403634
rect 114570 403398 114806 403634
rect 133930 403718 134166 403954
rect 134250 403718 134486 403954
rect 134570 403718 134806 403954
rect 133930 403398 134166 403634
rect 134250 403398 134486 403634
rect 134570 403398 134806 403634
rect 153930 403718 154166 403954
rect 154250 403718 154486 403954
rect 154570 403718 154806 403954
rect 153930 403398 154166 403634
rect 154250 403398 154486 403634
rect 154570 403398 154806 403634
rect 173930 403718 174166 403954
rect 174250 403718 174486 403954
rect 174570 403718 174806 403954
rect 173930 403398 174166 403634
rect 174250 403398 174486 403634
rect 174570 403398 174806 403634
rect 193930 403718 194166 403954
rect 194250 403718 194486 403954
rect 194570 403718 194806 403954
rect 193930 403398 194166 403634
rect 194250 403398 194486 403634
rect 194570 403398 194806 403634
rect 213930 403718 214166 403954
rect 214250 403718 214486 403954
rect 214570 403718 214806 403954
rect 213930 403398 214166 403634
rect 214250 403398 214486 403634
rect 214570 403398 214806 403634
rect 233930 403718 234166 403954
rect 234250 403718 234486 403954
rect 234570 403718 234806 403954
rect 233930 403398 234166 403634
rect 234250 403398 234486 403634
rect 234570 403398 234806 403634
rect 253930 403718 254166 403954
rect 254250 403718 254486 403954
rect 254570 403718 254806 403954
rect 253930 403398 254166 403634
rect 254250 403398 254486 403634
rect 254570 403398 254806 403634
rect 273930 403718 274166 403954
rect 274250 403718 274486 403954
rect 274570 403718 274806 403954
rect 273930 403398 274166 403634
rect 274250 403398 274486 403634
rect 274570 403398 274806 403634
rect 23930 399218 24166 399454
rect 24250 399218 24486 399454
rect 24570 399218 24806 399454
rect 23930 398898 24166 399134
rect 24250 398898 24486 399134
rect 24570 398898 24806 399134
rect 43930 399218 44166 399454
rect 44250 399218 44486 399454
rect 44570 399218 44806 399454
rect 43930 398898 44166 399134
rect 44250 398898 44486 399134
rect 44570 398898 44806 399134
rect 63930 399218 64166 399454
rect 64250 399218 64486 399454
rect 64570 399218 64806 399454
rect 63930 398898 64166 399134
rect 64250 398898 64486 399134
rect 64570 398898 64806 399134
rect 83930 399218 84166 399454
rect 84250 399218 84486 399454
rect 84570 399218 84806 399454
rect 83930 398898 84166 399134
rect 84250 398898 84486 399134
rect 84570 398898 84806 399134
rect 103930 399218 104166 399454
rect 104250 399218 104486 399454
rect 104570 399218 104806 399454
rect 103930 398898 104166 399134
rect 104250 398898 104486 399134
rect 104570 398898 104806 399134
rect 123930 399218 124166 399454
rect 124250 399218 124486 399454
rect 124570 399218 124806 399454
rect 123930 398898 124166 399134
rect 124250 398898 124486 399134
rect 124570 398898 124806 399134
rect 143930 399218 144166 399454
rect 144250 399218 144486 399454
rect 144570 399218 144806 399454
rect 143930 398898 144166 399134
rect 144250 398898 144486 399134
rect 144570 398898 144806 399134
rect 163930 399218 164166 399454
rect 164250 399218 164486 399454
rect 164570 399218 164806 399454
rect 163930 398898 164166 399134
rect 164250 398898 164486 399134
rect 164570 398898 164806 399134
rect 183930 399218 184166 399454
rect 184250 399218 184486 399454
rect 184570 399218 184806 399454
rect 183930 398898 184166 399134
rect 184250 398898 184486 399134
rect 184570 398898 184806 399134
rect 203930 399218 204166 399454
rect 204250 399218 204486 399454
rect 204570 399218 204806 399454
rect 203930 398898 204166 399134
rect 204250 398898 204486 399134
rect 204570 398898 204806 399134
rect 223930 399218 224166 399454
rect 224250 399218 224486 399454
rect 224570 399218 224806 399454
rect 223930 398898 224166 399134
rect 224250 398898 224486 399134
rect 224570 398898 224806 399134
rect 243930 399218 244166 399454
rect 244250 399218 244486 399454
rect 244570 399218 244806 399454
rect 243930 398898 244166 399134
rect 244250 398898 244486 399134
rect 244570 398898 244806 399134
rect 263930 399218 264166 399454
rect 264250 399218 264486 399454
rect 264570 399218 264806 399454
rect 263930 398898 264166 399134
rect 264250 398898 264486 399134
rect 264570 398898 264806 399134
rect 283930 399218 284166 399454
rect 284250 399218 284486 399454
rect 284570 399218 284806 399454
rect 283930 398898 284166 399134
rect 284250 398898 284486 399134
rect 284570 398898 284806 399134
rect 33930 367718 34166 367954
rect 34250 367718 34486 367954
rect 34570 367718 34806 367954
rect 33930 367398 34166 367634
rect 34250 367398 34486 367634
rect 34570 367398 34806 367634
rect 53930 367718 54166 367954
rect 54250 367718 54486 367954
rect 54570 367718 54806 367954
rect 53930 367398 54166 367634
rect 54250 367398 54486 367634
rect 54570 367398 54806 367634
rect 73930 367718 74166 367954
rect 74250 367718 74486 367954
rect 74570 367718 74806 367954
rect 73930 367398 74166 367634
rect 74250 367398 74486 367634
rect 74570 367398 74806 367634
rect 93930 367718 94166 367954
rect 94250 367718 94486 367954
rect 94570 367718 94806 367954
rect 93930 367398 94166 367634
rect 94250 367398 94486 367634
rect 94570 367398 94806 367634
rect 113930 367718 114166 367954
rect 114250 367718 114486 367954
rect 114570 367718 114806 367954
rect 113930 367398 114166 367634
rect 114250 367398 114486 367634
rect 114570 367398 114806 367634
rect 133930 367718 134166 367954
rect 134250 367718 134486 367954
rect 134570 367718 134806 367954
rect 133930 367398 134166 367634
rect 134250 367398 134486 367634
rect 134570 367398 134806 367634
rect 153930 367718 154166 367954
rect 154250 367718 154486 367954
rect 154570 367718 154806 367954
rect 153930 367398 154166 367634
rect 154250 367398 154486 367634
rect 154570 367398 154806 367634
rect 173930 367718 174166 367954
rect 174250 367718 174486 367954
rect 174570 367718 174806 367954
rect 173930 367398 174166 367634
rect 174250 367398 174486 367634
rect 174570 367398 174806 367634
rect 193930 367718 194166 367954
rect 194250 367718 194486 367954
rect 194570 367718 194806 367954
rect 193930 367398 194166 367634
rect 194250 367398 194486 367634
rect 194570 367398 194806 367634
rect 213930 367718 214166 367954
rect 214250 367718 214486 367954
rect 214570 367718 214806 367954
rect 213930 367398 214166 367634
rect 214250 367398 214486 367634
rect 214570 367398 214806 367634
rect 233930 367718 234166 367954
rect 234250 367718 234486 367954
rect 234570 367718 234806 367954
rect 233930 367398 234166 367634
rect 234250 367398 234486 367634
rect 234570 367398 234806 367634
rect 253930 367718 254166 367954
rect 254250 367718 254486 367954
rect 254570 367718 254806 367954
rect 253930 367398 254166 367634
rect 254250 367398 254486 367634
rect 254570 367398 254806 367634
rect 273930 367718 274166 367954
rect 274250 367718 274486 367954
rect 274570 367718 274806 367954
rect 273930 367398 274166 367634
rect 274250 367398 274486 367634
rect 274570 367398 274806 367634
rect 23930 363218 24166 363454
rect 24250 363218 24486 363454
rect 24570 363218 24806 363454
rect 23930 362898 24166 363134
rect 24250 362898 24486 363134
rect 24570 362898 24806 363134
rect 43930 363218 44166 363454
rect 44250 363218 44486 363454
rect 44570 363218 44806 363454
rect 43930 362898 44166 363134
rect 44250 362898 44486 363134
rect 44570 362898 44806 363134
rect 63930 363218 64166 363454
rect 64250 363218 64486 363454
rect 64570 363218 64806 363454
rect 63930 362898 64166 363134
rect 64250 362898 64486 363134
rect 64570 362898 64806 363134
rect 83930 363218 84166 363454
rect 84250 363218 84486 363454
rect 84570 363218 84806 363454
rect 83930 362898 84166 363134
rect 84250 362898 84486 363134
rect 84570 362898 84806 363134
rect 103930 363218 104166 363454
rect 104250 363218 104486 363454
rect 104570 363218 104806 363454
rect 103930 362898 104166 363134
rect 104250 362898 104486 363134
rect 104570 362898 104806 363134
rect 123930 363218 124166 363454
rect 124250 363218 124486 363454
rect 124570 363218 124806 363454
rect 123930 362898 124166 363134
rect 124250 362898 124486 363134
rect 124570 362898 124806 363134
rect 143930 363218 144166 363454
rect 144250 363218 144486 363454
rect 144570 363218 144806 363454
rect 143930 362898 144166 363134
rect 144250 362898 144486 363134
rect 144570 362898 144806 363134
rect 163930 363218 164166 363454
rect 164250 363218 164486 363454
rect 164570 363218 164806 363454
rect 163930 362898 164166 363134
rect 164250 362898 164486 363134
rect 164570 362898 164806 363134
rect 183930 363218 184166 363454
rect 184250 363218 184486 363454
rect 184570 363218 184806 363454
rect 183930 362898 184166 363134
rect 184250 362898 184486 363134
rect 184570 362898 184806 363134
rect 203930 363218 204166 363454
rect 204250 363218 204486 363454
rect 204570 363218 204806 363454
rect 203930 362898 204166 363134
rect 204250 362898 204486 363134
rect 204570 362898 204806 363134
rect 223930 363218 224166 363454
rect 224250 363218 224486 363454
rect 224570 363218 224806 363454
rect 223930 362898 224166 363134
rect 224250 362898 224486 363134
rect 224570 362898 224806 363134
rect 243930 363218 244166 363454
rect 244250 363218 244486 363454
rect 244570 363218 244806 363454
rect 243930 362898 244166 363134
rect 244250 362898 244486 363134
rect 244570 362898 244806 363134
rect 263930 363218 264166 363454
rect 264250 363218 264486 363454
rect 264570 363218 264806 363454
rect 263930 362898 264166 363134
rect 264250 362898 264486 363134
rect 264570 362898 264806 363134
rect 283930 363218 284166 363454
rect 284250 363218 284486 363454
rect 284570 363218 284806 363454
rect 283930 362898 284166 363134
rect 284250 362898 284486 363134
rect 284570 362898 284806 363134
rect 33930 295718 34166 295954
rect 34250 295718 34486 295954
rect 34570 295718 34806 295954
rect 33930 295398 34166 295634
rect 34250 295398 34486 295634
rect 34570 295398 34806 295634
rect 53930 295718 54166 295954
rect 54250 295718 54486 295954
rect 54570 295718 54806 295954
rect 53930 295398 54166 295634
rect 54250 295398 54486 295634
rect 54570 295398 54806 295634
rect 73930 295718 74166 295954
rect 74250 295718 74486 295954
rect 74570 295718 74806 295954
rect 73930 295398 74166 295634
rect 74250 295398 74486 295634
rect 74570 295398 74806 295634
rect 93930 295718 94166 295954
rect 94250 295718 94486 295954
rect 94570 295718 94806 295954
rect 93930 295398 94166 295634
rect 94250 295398 94486 295634
rect 94570 295398 94806 295634
rect 113930 295718 114166 295954
rect 114250 295718 114486 295954
rect 114570 295718 114806 295954
rect 113930 295398 114166 295634
rect 114250 295398 114486 295634
rect 114570 295398 114806 295634
rect 133930 295718 134166 295954
rect 134250 295718 134486 295954
rect 134570 295718 134806 295954
rect 133930 295398 134166 295634
rect 134250 295398 134486 295634
rect 134570 295398 134806 295634
rect 153930 295718 154166 295954
rect 154250 295718 154486 295954
rect 154570 295718 154806 295954
rect 153930 295398 154166 295634
rect 154250 295398 154486 295634
rect 154570 295398 154806 295634
rect 173930 295718 174166 295954
rect 174250 295718 174486 295954
rect 174570 295718 174806 295954
rect 173930 295398 174166 295634
rect 174250 295398 174486 295634
rect 174570 295398 174806 295634
rect 193930 295718 194166 295954
rect 194250 295718 194486 295954
rect 194570 295718 194806 295954
rect 193930 295398 194166 295634
rect 194250 295398 194486 295634
rect 194570 295398 194806 295634
rect 213930 295718 214166 295954
rect 214250 295718 214486 295954
rect 214570 295718 214806 295954
rect 213930 295398 214166 295634
rect 214250 295398 214486 295634
rect 214570 295398 214806 295634
rect 233930 295718 234166 295954
rect 234250 295718 234486 295954
rect 234570 295718 234806 295954
rect 233930 295398 234166 295634
rect 234250 295398 234486 295634
rect 234570 295398 234806 295634
rect 253930 295718 254166 295954
rect 254250 295718 254486 295954
rect 254570 295718 254806 295954
rect 253930 295398 254166 295634
rect 254250 295398 254486 295634
rect 254570 295398 254806 295634
rect 273930 295718 274166 295954
rect 274250 295718 274486 295954
rect 274570 295718 274806 295954
rect 273930 295398 274166 295634
rect 274250 295398 274486 295634
rect 274570 295398 274806 295634
rect 23930 291218 24166 291454
rect 24250 291218 24486 291454
rect 24570 291218 24806 291454
rect 23930 290898 24166 291134
rect 24250 290898 24486 291134
rect 24570 290898 24806 291134
rect 43930 291218 44166 291454
rect 44250 291218 44486 291454
rect 44570 291218 44806 291454
rect 43930 290898 44166 291134
rect 44250 290898 44486 291134
rect 44570 290898 44806 291134
rect 63930 291218 64166 291454
rect 64250 291218 64486 291454
rect 64570 291218 64806 291454
rect 63930 290898 64166 291134
rect 64250 290898 64486 291134
rect 64570 290898 64806 291134
rect 83930 291218 84166 291454
rect 84250 291218 84486 291454
rect 84570 291218 84806 291454
rect 83930 290898 84166 291134
rect 84250 290898 84486 291134
rect 84570 290898 84806 291134
rect 103930 291218 104166 291454
rect 104250 291218 104486 291454
rect 104570 291218 104806 291454
rect 103930 290898 104166 291134
rect 104250 290898 104486 291134
rect 104570 290898 104806 291134
rect 123930 291218 124166 291454
rect 124250 291218 124486 291454
rect 124570 291218 124806 291454
rect 123930 290898 124166 291134
rect 124250 290898 124486 291134
rect 124570 290898 124806 291134
rect 143930 291218 144166 291454
rect 144250 291218 144486 291454
rect 144570 291218 144806 291454
rect 143930 290898 144166 291134
rect 144250 290898 144486 291134
rect 144570 290898 144806 291134
rect 163930 291218 164166 291454
rect 164250 291218 164486 291454
rect 164570 291218 164806 291454
rect 163930 290898 164166 291134
rect 164250 290898 164486 291134
rect 164570 290898 164806 291134
rect 183930 291218 184166 291454
rect 184250 291218 184486 291454
rect 184570 291218 184806 291454
rect 183930 290898 184166 291134
rect 184250 290898 184486 291134
rect 184570 290898 184806 291134
rect 203930 291218 204166 291454
rect 204250 291218 204486 291454
rect 204570 291218 204806 291454
rect 203930 290898 204166 291134
rect 204250 290898 204486 291134
rect 204570 290898 204806 291134
rect 223930 291218 224166 291454
rect 224250 291218 224486 291454
rect 224570 291218 224806 291454
rect 223930 290898 224166 291134
rect 224250 290898 224486 291134
rect 224570 290898 224806 291134
rect 243930 291218 244166 291454
rect 244250 291218 244486 291454
rect 244570 291218 244806 291454
rect 243930 290898 244166 291134
rect 244250 290898 244486 291134
rect 244570 290898 244806 291134
rect 263930 291218 264166 291454
rect 264250 291218 264486 291454
rect 264570 291218 264806 291454
rect 263930 290898 264166 291134
rect 264250 290898 264486 291134
rect 264570 290898 264806 291134
rect 283930 291218 284166 291454
rect 284250 291218 284486 291454
rect 284570 291218 284806 291454
rect 283930 290898 284166 291134
rect 284250 290898 284486 291134
rect 284570 290898 284806 291134
rect 33930 259718 34166 259954
rect 34250 259718 34486 259954
rect 34570 259718 34806 259954
rect 33930 259398 34166 259634
rect 34250 259398 34486 259634
rect 34570 259398 34806 259634
rect 53930 259718 54166 259954
rect 54250 259718 54486 259954
rect 54570 259718 54806 259954
rect 53930 259398 54166 259634
rect 54250 259398 54486 259634
rect 54570 259398 54806 259634
rect 73930 259718 74166 259954
rect 74250 259718 74486 259954
rect 74570 259718 74806 259954
rect 73930 259398 74166 259634
rect 74250 259398 74486 259634
rect 74570 259398 74806 259634
rect 93930 259718 94166 259954
rect 94250 259718 94486 259954
rect 94570 259718 94806 259954
rect 93930 259398 94166 259634
rect 94250 259398 94486 259634
rect 94570 259398 94806 259634
rect 113930 259718 114166 259954
rect 114250 259718 114486 259954
rect 114570 259718 114806 259954
rect 113930 259398 114166 259634
rect 114250 259398 114486 259634
rect 114570 259398 114806 259634
rect 133930 259718 134166 259954
rect 134250 259718 134486 259954
rect 134570 259718 134806 259954
rect 133930 259398 134166 259634
rect 134250 259398 134486 259634
rect 134570 259398 134806 259634
rect 153930 259718 154166 259954
rect 154250 259718 154486 259954
rect 154570 259718 154806 259954
rect 153930 259398 154166 259634
rect 154250 259398 154486 259634
rect 154570 259398 154806 259634
rect 173930 259718 174166 259954
rect 174250 259718 174486 259954
rect 174570 259718 174806 259954
rect 173930 259398 174166 259634
rect 174250 259398 174486 259634
rect 174570 259398 174806 259634
rect 193930 259718 194166 259954
rect 194250 259718 194486 259954
rect 194570 259718 194806 259954
rect 193930 259398 194166 259634
rect 194250 259398 194486 259634
rect 194570 259398 194806 259634
rect 213930 259718 214166 259954
rect 214250 259718 214486 259954
rect 214570 259718 214806 259954
rect 213930 259398 214166 259634
rect 214250 259398 214486 259634
rect 214570 259398 214806 259634
rect 233930 259718 234166 259954
rect 234250 259718 234486 259954
rect 234570 259718 234806 259954
rect 233930 259398 234166 259634
rect 234250 259398 234486 259634
rect 234570 259398 234806 259634
rect 253930 259718 254166 259954
rect 254250 259718 254486 259954
rect 254570 259718 254806 259954
rect 253930 259398 254166 259634
rect 254250 259398 254486 259634
rect 254570 259398 254806 259634
rect 273930 259718 274166 259954
rect 274250 259718 274486 259954
rect 274570 259718 274806 259954
rect 273930 259398 274166 259634
rect 274250 259398 274486 259634
rect 274570 259398 274806 259634
rect 23930 255218 24166 255454
rect 24250 255218 24486 255454
rect 24570 255218 24806 255454
rect 23930 254898 24166 255134
rect 24250 254898 24486 255134
rect 24570 254898 24806 255134
rect 43930 255218 44166 255454
rect 44250 255218 44486 255454
rect 44570 255218 44806 255454
rect 43930 254898 44166 255134
rect 44250 254898 44486 255134
rect 44570 254898 44806 255134
rect 63930 255218 64166 255454
rect 64250 255218 64486 255454
rect 64570 255218 64806 255454
rect 63930 254898 64166 255134
rect 64250 254898 64486 255134
rect 64570 254898 64806 255134
rect 83930 255218 84166 255454
rect 84250 255218 84486 255454
rect 84570 255218 84806 255454
rect 83930 254898 84166 255134
rect 84250 254898 84486 255134
rect 84570 254898 84806 255134
rect 103930 255218 104166 255454
rect 104250 255218 104486 255454
rect 104570 255218 104806 255454
rect 103930 254898 104166 255134
rect 104250 254898 104486 255134
rect 104570 254898 104806 255134
rect 123930 255218 124166 255454
rect 124250 255218 124486 255454
rect 124570 255218 124806 255454
rect 123930 254898 124166 255134
rect 124250 254898 124486 255134
rect 124570 254898 124806 255134
rect 143930 255218 144166 255454
rect 144250 255218 144486 255454
rect 144570 255218 144806 255454
rect 143930 254898 144166 255134
rect 144250 254898 144486 255134
rect 144570 254898 144806 255134
rect 163930 255218 164166 255454
rect 164250 255218 164486 255454
rect 164570 255218 164806 255454
rect 163930 254898 164166 255134
rect 164250 254898 164486 255134
rect 164570 254898 164806 255134
rect 183930 255218 184166 255454
rect 184250 255218 184486 255454
rect 184570 255218 184806 255454
rect 183930 254898 184166 255134
rect 184250 254898 184486 255134
rect 184570 254898 184806 255134
rect 203930 255218 204166 255454
rect 204250 255218 204486 255454
rect 204570 255218 204806 255454
rect 203930 254898 204166 255134
rect 204250 254898 204486 255134
rect 204570 254898 204806 255134
rect 223930 255218 224166 255454
rect 224250 255218 224486 255454
rect 224570 255218 224806 255454
rect 223930 254898 224166 255134
rect 224250 254898 224486 255134
rect 224570 254898 224806 255134
rect 243930 255218 244166 255454
rect 244250 255218 244486 255454
rect 244570 255218 244806 255454
rect 243930 254898 244166 255134
rect 244250 254898 244486 255134
rect 244570 254898 244806 255134
rect 263930 255218 264166 255454
rect 264250 255218 264486 255454
rect 264570 255218 264806 255454
rect 263930 254898 264166 255134
rect 264250 254898 264486 255134
rect 264570 254898 264806 255134
rect 283930 255218 284166 255454
rect 284250 255218 284486 255454
rect 284570 255218 284806 255454
rect 283930 254898 284166 255134
rect 284250 254898 284486 255134
rect 284570 254898 284806 255134
rect 33930 223718 34166 223954
rect 34250 223718 34486 223954
rect 34570 223718 34806 223954
rect 33930 223398 34166 223634
rect 34250 223398 34486 223634
rect 34570 223398 34806 223634
rect 53930 223718 54166 223954
rect 54250 223718 54486 223954
rect 54570 223718 54806 223954
rect 53930 223398 54166 223634
rect 54250 223398 54486 223634
rect 54570 223398 54806 223634
rect 73930 223718 74166 223954
rect 74250 223718 74486 223954
rect 74570 223718 74806 223954
rect 73930 223398 74166 223634
rect 74250 223398 74486 223634
rect 74570 223398 74806 223634
rect 93930 223718 94166 223954
rect 94250 223718 94486 223954
rect 94570 223718 94806 223954
rect 93930 223398 94166 223634
rect 94250 223398 94486 223634
rect 94570 223398 94806 223634
rect 113930 223718 114166 223954
rect 114250 223718 114486 223954
rect 114570 223718 114806 223954
rect 113930 223398 114166 223634
rect 114250 223398 114486 223634
rect 114570 223398 114806 223634
rect 133930 223718 134166 223954
rect 134250 223718 134486 223954
rect 134570 223718 134806 223954
rect 133930 223398 134166 223634
rect 134250 223398 134486 223634
rect 134570 223398 134806 223634
rect 153930 223718 154166 223954
rect 154250 223718 154486 223954
rect 154570 223718 154806 223954
rect 153930 223398 154166 223634
rect 154250 223398 154486 223634
rect 154570 223398 154806 223634
rect 173930 223718 174166 223954
rect 174250 223718 174486 223954
rect 174570 223718 174806 223954
rect 173930 223398 174166 223634
rect 174250 223398 174486 223634
rect 174570 223398 174806 223634
rect 193930 223718 194166 223954
rect 194250 223718 194486 223954
rect 194570 223718 194806 223954
rect 193930 223398 194166 223634
rect 194250 223398 194486 223634
rect 194570 223398 194806 223634
rect 213930 223718 214166 223954
rect 214250 223718 214486 223954
rect 214570 223718 214806 223954
rect 213930 223398 214166 223634
rect 214250 223398 214486 223634
rect 214570 223398 214806 223634
rect 233930 223718 234166 223954
rect 234250 223718 234486 223954
rect 234570 223718 234806 223954
rect 233930 223398 234166 223634
rect 234250 223398 234486 223634
rect 234570 223398 234806 223634
rect 253930 223718 254166 223954
rect 254250 223718 254486 223954
rect 254570 223718 254806 223954
rect 253930 223398 254166 223634
rect 254250 223398 254486 223634
rect 254570 223398 254806 223634
rect 273930 223718 274166 223954
rect 274250 223718 274486 223954
rect 274570 223718 274806 223954
rect 273930 223398 274166 223634
rect 274250 223398 274486 223634
rect 274570 223398 274806 223634
rect 23930 219218 24166 219454
rect 24250 219218 24486 219454
rect 24570 219218 24806 219454
rect 23930 218898 24166 219134
rect 24250 218898 24486 219134
rect 24570 218898 24806 219134
rect 43930 219218 44166 219454
rect 44250 219218 44486 219454
rect 44570 219218 44806 219454
rect 43930 218898 44166 219134
rect 44250 218898 44486 219134
rect 44570 218898 44806 219134
rect 63930 219218 64166 219454
rect 64250 219218 64486 219454
rect 64570 219218 64806 219454
rect 63930 218898 64166 219134
rect 64250 218898 64486 219134
rect 64570 218898 64806 219134
rect 83930 219218 84166 219454
rect 84250 219218 84486 219454
rect 84570 219218 84806 219454
rect 83930 218898 84166 219134
rect 84250 218898 84486 219134
rect 84570 218898 84806 219134
rect 103930 219218 104166 219454
rect 104250 219218 104486 219454
rect 104570 219218 104806 219454
rect 103930 218898 104166 219134
rect 104250 218898 104486 219134
rect 104570 218898 104806 219134
rect 123930 219218 124166 219454
rect 124250 219218 124486 219454
rect 124570 219218 124806 219454
rect 123930 218898 124166 219134
rect 124250 218898 124486 219134
rect 124570 218898 124806 219134
rect 143930 219218 144166 219454
rect 144250 219218 144486 219454
rect 144570 219218 144806 219454
rect 143930 218898 144166 219134
rect 144250 218898 144486 219134
rect 144570 218898 144806 219134
rect 163930 219218 164166 219454
rect 164250 219218 164486 219454
rect 164570 219218 164806 219454
rect 163930 218898 164166 219134
rect 164250 218898 164486 219134
rect 164570 218898 164806 219134
rect 183930 219218 184166 219454
rect 184250 219218 184486 219454
rect 184570 219218 184806 219454
rect 183930 218898 184166 219134
rect 184250 218898 184486 219134
rect 184570 218898 184806 219134
rect 203930 219218 204166 219454
rect 204250 219218 204486 219454
rect 204570 219218 204806 219454
rect 203930 218898 204166 219134
rect 204250 218898 204486 219134
rect 204570 218898 204806 219134
rect 223930 219218 224166 219454
rect 224250 219218 224486 219454
rect 224570 219218 224806 219454
rect 223930 218898 224166 219134
rect 224250 218898 224486 219134
rect 224570 218898 224806 219134
rect 243930 219218 244166 219454
rect 244250 219218 244486 219454
rect 244570 219218 244806 219454
rect 243930 218898 244166 219134
rect 244250 218898 244486 219134
rect 244570 218898 244806 219134
rect 263930 219218 264166 219454
rect 264250 219218 264486 219454
rect 264570 219218 264806 219454
rect 263930 218898 264166 219134
rect 264250 218898 264486 219134
rect 264570 218898 264806 219134
rect 283930 219218 284166 219454
rect 284250 219218 284486 219454
rect 284570 219218 284806 219454
rect 283930 218898 284166 219134
rect 284250 218898 284486 219134
rect 284570 218898 284806 219134
rect 23930 183218 24166 183454
rect 24250 183218 24486 183454
rect 24570 183218 24806 183454
rect 23930 182898 24166 183134
rect 24250 182898 24486 183134
rect 24570 182898 24806 183134
rect 43930 183218 44166 183454
rect 44250 183218 44486 183454
rect 44570 183218 44806 183454
rect 43930 182898 44166 183134
rect 44250 182898 44486 183134
rect 44570 182898 44806 183134
rect 63930 183218 64166 183454
rect 64250 183218 64486 183454
rect 64570 183218 64806 183454
rect 63930 182898 64166 183134
rect 64250 182898 64486 183134
rect 64570 182898 64806 183134
rect 83930 183218 84166 183454
rect 84250 183218 84486 183454
rect 84570 183218 84806 183454
rect 83930 182898 84166 183134
rect 84250 182898 84486 183134
rect 84570 182898 84806 183134
rect 103930 183218 104166 183454
rect 104250 183218 104486 183454
rect 104570 183218 104806 183454
rect 103930 182898 104166 183134
rect 104250 182898 104486 183134
rect 104570 182898 104806 183134
rect 123930 183218 124166 183454
rect 124250 183218 124486 183454
rect 124570 183218 124806 183454
rect 123930 182898 124166 183134
rect 124250 182898 124486 183134
rect 124570 182898 124806 183134
rect 143930 183218 144166 183454
rect 144250 183218 144486 183454
rect 144570 183218 144806 183454
rect 143930 182898 144166 183134
rect 144250 182898 144486 183134
rect 144570 182898 144806 183134
rect 163930 183218 164166 183454
rect 164250 183218 164486 183454
rect 164570 183218 164806 183454
rect 163930 182898 164166 183134
rect 164250 182898 164486 183134
rect 164570 182898 164806 183134
rect 183930 183218 184166 183454
rect 184250 183218 184486 183454
rect 184570 183218 184806 183454
rect 183930 182898 184166 183134
rect 184250 182898 184486 183134
rect 184570 182898 184806 183134
rect 203930 183218 204166 183454
rect 204250 183218 204486 183454
rect 204570 183218 204806 183454
rect 203930 182898 204166 183134
rect 204250 182898 204486 183134
rect 204570 182898 204806 183134
rect 223930 183218 224166 183454
rect 224250 183218 224486 183454
rect 224570 183218 224806 183454
rect 223930 182898 224166 183134
rect 224250 182898 224486 183134
rect 224570 182898 224806 183134
rect 243930 183218 244166 183454
rect 244250 183218 244486 183454
rect 244570 183218 244806 183454
rect 243930 182898 244166 183134
rect 244250 182898 244486 183134
rect 244570 182898 244806 183134
rect 263930 183218 264166 183454
rect 264250 183218 264486 183454
rect 264570 183218 264806 183454
rect 263930 182898 264166 183134
rect 264250 182898 264486 183134
rect 264570 182898 264806 183134
rect 283930 183218 284166 183454
rect 284250 183218 284486 183454
rect 284570 183218 284806 183454
rect 283930 182898 284166 183134
rect 284250 182898 284486 183134
rect 284570 182898 284806 183134
rect 33930 151718 34166 151954
rect 34250 151718 34486 151954
rect 34570 151718 34806 151954
rect 33930 151398 34166 151634
rect 34250 151398 34486 151634
rect 34570 151398 34806 151634
rect 53930 151718 54166 151954
rect 54250 151718 54486 151954
rect 54570 151718 54806 151954
rect 53930 151398 54166 151634
rect 54250 151398 54486 151634
rect 54570 151398 54806 151634
rect 73930 151718 74166 151954
rect 74250 151718 74486 151954
rect 74570 151718 74806 151954
rect 73930 151398 74166 151634
rect 74250 151398 74486 151634
rect 74570 151398 74806 151634
rect 93930 151718 94166 151954
rect 94250 151718 94486 151954
rect 94570 151718 94806 151954
rect 93930 151398 94166 151634
rect 94250 151398 94486 151634
rect 94570 151398 94806 151634
rect 113930 151718 114166 151954
rect 114250 151718 114486 151954
rect 114570 151718 114806 151954
rect 113930 151398 114166 151634
rect 114250 151398 114486 151634
rect 114570 151398 114806 151634
rect 133930 151718 134166 151954
rect 134250 151718 134486 151954
rect 134570 151718 134806 151954
rect 133930 151398 134166 151634
rect 134250 151398 134486 151634
rect 134570 151398 134806 151634
rect 153930 151718 154166 151954
rect 154250 151718 154486 151954
rect 154570 151718 154806 151954
rect 153930 151398 154166 151634
rect 154250 151398 154486 151634
rect 154570 151398 154806 151634
rect 173930 151718 174166 151954
rect 174250 151718 174486 151954
rect 174570 151718 174806 151954
rect 173930 151398 174166 151634
rect 174250 151398 174486 151634
rect 174570 151398 174806 151634
rect 193930 151718 194166 151954
rect 194250 151718 194486 151954
rect 194570 151718 194806 151954
rect 193930 151398 194166 151634
rect 194250 151398 194486 151634
rect 194570 151398 194806 151634
rect 213930 151718 214166 151954
rect 214250 151718 214486 151954
rect 214570 151718 214806 151954
rect 213930 151398 214166 151634
rect 214250 151398 214486 151634
rect 214570 151398 214806 151634
rect 233930 151718 234166 151954
rect 234250 151718 234486 151954
rect 234570 151718 234806 151954
rect 233930 151398 234166 151634
rect 234250 151398 234486 151634
rect 234570 151398 234806 151634
rect 253930 151718 254166 151954
rect 254250 151718 254486 151954
rect 254570 151718 254806 151954
rect 253930 151398 254166 151634
rect 254250 151398 254486 151634
rect 254570 151398 254806 151634
rect 273930 151718 274166 151954
rect 274250 151718 274486 151954
rect 274570 151718 274806 151954
rect 273930 151398 274166 151634
rect 274250 151398 274486 151634
rect 274570 151398 274806 151634
rect 23930 147218 24166 147454
rect 24250 147218 24486 147454
rect 24570 147218 24806 147454
rect 23930 146898 24166 147134
rect 24250 146898 24486 147134
rect 24570 146898 24806 147134
rect 43930 147218 44166 147454
rect 44250 147218 44486 147454
rect 44570 147218 44806 147454
rect 43930 146898 44166 147134
rect 44250 146898 44486 147134
rect 44570 146898 44806 147134
rect 63930 147218 64166 147454
rect 64250 147218 64486 147454
rect 64570 147218 64806 147454
rect 63930 146898 64166 147134
rect 64250 146898 64486 147134
rect 64570 146898 64806 147134
rect 83930 147218 84166 147454
rect 84250 147218 84486 147454
rect 84570 147218 84806 147454
rect 83930 146898 84166 147134
rect 84250 146898 84486 147134
rect 84570 146898 84806 147134
rect 103930 147218 104166 147454
rect 104250 147218 104486 147454
rect 104570 147218 104806 147454
rect 103930 146898 104166 147134
rect 104250 146898 104486 147134
rect 104570 146898 104806 147134
rect 123930 147218 124166 147454
rect 124250 147218 124486 147454
rect 124570 147218 124806 147454
rect 123930 146898 124166 147134
rect 124250 146898 124486 147134
rect 124570 146898 124806 147134
rect 143930 147218 144166 147454
rect 144250 147218 144486 147454
rect 144570 147218 144806 147454
rect 143930 146898 144166 147134
rect 144250 146898 144486 147134
rect 144570 146898 144806 147134
rect 163930 147218 164166 147454
rect 164250 147218 164486 147454
rect 164570 147218 164806 147454
rect 163930 146898 164166 147134
rect 164250 146898 164486 147134
rect 164570 146898 164806 147134
rect 183930 147218 184166 147454
rect 184250 147218 184486 147454
rect 184570 147218 184806 147454
rect 183930 146898 184166 147134
rect 184250 146898 184486 147134
rect 184570 146898 184806 147134
rect 203930 147218 204166 147454
rect 204250 147218 204486 147454
rect 204570 147218 204806 147454
rect 203930 146898 204166 147134
rect 204250 146898 204486 147134
rect 204570 146898 204806 147134
rect 223930 147218 224166 147454
rect 224250 147218 224486 147454
rect 224570 147218 224806 147454
rect 223930 146898 224166 147134
rect 224250 146898 224486 147134
rect 224570 146898 224806 147134
rect 243930 147218 244166 147454
rect 244250 147218 244486 147454
rect 244570 147218 244806 147454
rect 243930 146898 244166 147134
rect 244250 146898 244486 147134
rect 244570 146898 244806 147134
rect 263930 147218 264166 147454
rect 264250 147218 264486 147454
rect 264570 147218 264806 147454
rect 263930 146898 264166 147134
rect 264250 146898 264486 147134
rect 264570 146898 264806 147134
rect 283930 147218 284166 147454
rect 284250 147218 284486 147454
rect 284570 147218 284806 147454
rect 283930 146898 284166 147134
rect 284250 146898 284486 147134
rect 284570 146898 284806 147134
rect 33930 115718 34166 115954
rect 34250 115718 34486 115954
rect 34570 115718 34806 115954
rect 33930 115398 34166 115634
rect 34250 115398 34486 115634
rect 34570 115398 34806 115634
rect 53930 115718 54166 115954
rect 54250 115718 54486 115954
rect 54570 115718 54806 115954
rect 53930 115398 54166 115634
rect 54250 115398 54486 115634
rect 54570 115398 54806 115634
rect 73930 115718 74166 115954
rect 74250 115718 74486 115954
rect 74570 115718 74806 115954
rect 73930 115398 74166 115634
rect 74250 115398 74486 115634
rect 74570 115398 74806 115634
rect 93930 115718 94166 115954
rect 94250 115718 94486 115954
rect 94570 115718 94806 115954
rect 93930 115398 94166 115634
rect 94250 115398 94486 115634
rect 94570 115398 94806 115634
rect 113930 115718 114166 115954
rect 114250 115718 114486 115954
rect 114570 115718 114806 115954
rect 113930 115398 114166 115634
rect 114250 115398 114486 115634
rect 114570 115398 114806 115634
rect 133930 115718 134166 115954
rect 134250 115718 134486 115954
rect 134570 115718 134806 115954
rect 133930 115398 134166 115634
rect 134250 115398 134486 115634
rect 134570 115398 134806 115634
rect 153930 115718 154166 115954
rect 154250 115718 154486 115954
rect 154570 115718 154806 115954
rect 153930 115398 154166 115634
rect 154250 115398 154486 115634
rect 154570 115398 154806 115634
rect 173930 115718 174166 115954
rect 174250 115718 174486 115954
rect 174570 115718 174806 115954
rect 173930 115398 174166 115634
rect 174250 115398 174486 115634
rect 174570 115398 174806 115634
rect 193930 115718 194166 115954
rect 194250 115718 194486 115954
rect 194570 115718 194806 115954
rect 193930 115398 194166 115634
rect 194250 115398 194486 115634
rect 194570 115398 194806 115634
rect 213930 115718 214166 115954
rect 214250 115718 214486 115954
rect 214570 115718 214806 115954
rect 213930 115398 214166 115634
rect 214250 115398 214486 115634
rect 214570 115398 214806 115634
rect 233930 115718 234166 115954
rect 234250 115718 234486 115954
rect 234570 115718 234806 115954
rect 233930 115398 234166 115634
rect 234250 115398 234486 115634
rect 234570 115398 234806 115634
rect 253930 115718 254166 115954
rect 254250 115718 254486 115954
rect 254570 115718 254806 115954
rect 253930 115398 254166 115634
rect 254250 115398 254486 115634
rect 254570 115398 254806 115634
rect 273930 115718 274166 115954
rect 274250 115718 274486 115954
rect 274570 115718 274806 115954
rect 273930 115398 274166 115634
rect 274250 115398 274486 115634
rect 274570 115398 274806 115634
rect 23930 111218 24166 111454
rect 24250 111218 24486 111454
rect 24570 111218 24806 111454
rect 23930 110898 24166 111134
rect 24250 110898 24486 111134
rect 24570 110898 24806 111134
rect 43930 111218 44166 111454
rect 44250 111218 44486 111454
rect 44570 111218 44806 111454
rect 43930 110898 44166 111134
rect 44250 110898 44486 111134
rect 44570 110898 44806 111134
rect 63930 111218 64166 111454
rect 64250 111218 64486 111454
rect 64570 111218 64806 111454
rect 63930 110898 64166 111134
rect 64250 110898 64486 111134
rect 64570 110898 64806 111134
rect 83930 111218 84166 111454
rect 84250 111218 84486 111454
rect 84570 111218 84806 111454
rect 83930 110898 84166 111134
rect 84250 110898 84486 111134
rect 84570 110898 84806 111134
rect 103930 111218 104166 111454
rect 104250 111218 104486 111454
rect 104570 111218 104806 111454
rect 103930 110898 104166 111134
rect 104250 110898 104486 111134
rect 104570 110898 104806 111134
rect 123930 111218 124166 111454
rect 124250 111218 124486 111454
rect 124570 111218 124806 111454
rect 123930 110898 124166 111134
rect 124250 110898 124486 111134
rect 124570 110898 124806 111134
rect 143930 111218 144166 111454
rect 144250 111218 144486 111454
rect 144570 111218 144806 111454
rect 143930 110898 144166 111134
rect 144250 110898 144486 111134
rect 144570 110898 144806 111134
rect 163930 111218 164166 111454
rect 164250 111218 164486 111454
rect 164570 111218 164806 111454
rect 163930 110898 164166 111134
rect 164250 110898 164486 111134
rect 164570 110898 164806 111134
rect 183930 111218 184166 111454
rect 184250 111218 184486 111454
rect 184570 111218 184806 111454
rect 183930 110898 184166 111134
rect 184250 110898 184486 111134
rect 184570 110898 184806 111134
rect 203930 111218 204166 111454
rect 204250 111218 204486 111454
rect 204570 111218 204806 111454
rect 203930 110898 204166 111134
rect 204250 110898 204486 111134
rect 204570 110898 204806 111134
rect 223930 111218 224166 111454
rect 224250 111218 224486 111454
rect 224570 111218 224806 111454
rect 223930 110898 224166 111134
rect 224250 110898 224486 111134
rect 224570 110898 224806 111134
rect 243930 111218 244166 111454
rect 244250 111218 244486 111454
rect 244570 111218 244806 111454
rect 243930 110898 244166 111134
rect 244250 110898 244486 111134
rect 244570 110898 244806 111134
rect 263930 111218 264166 111454
rect 264250 111218 264486 111454
rect 264570 111218 264806 111454
rect 263930 110898 264166 111134
rect 264250 110898 264486 111134
rect 264570 110898 264806 111134
rect 283930 111218 284166 111454
rect 284250 111218 284486 111454
rect 284570 111218 284806 111454
rect 283930 110898 284166 111134
rect 284250 110898 284486 111134
rect 284570 110898 284806 111134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 313930 691718 314166 691954
rect 314250 691718 314486 691954
rect 314570 691718 314806 691954
rect 313930 691398 314166 691634
rect 314250 691398 314486 691634
rect 314570 691398 314806 691634
rect 333930 691718 334166 691954
rect 334250 691718 334486 691954
rect 334570 691718 334806 691954
rect 333930 691398 334166 691634
rect 334250 691398 334486 691634
rect 334570 691398 334806 691634
rect 353930 691718 354166 691954
rect 354250 691718 354486 691954
rect 354570 691718 354806 691954
rect 353930 691398 354166 691634
rect 354250 691398 354486 691634
rect 354570 691398 354806 691634
rect 373930 691718 374166 691954
rect 374250 691718 374486 691954
rect 374570 691718 374806 691954
rect 373930 691398 374166 691634
rect 374250 691398 374486 691634
rect 374570 691398 374806 691634
rect 393930 691718 394166 691954
rect 394250 691718 394486 691954
rect 394570 691718 394806 691954
rect 393930 691398 394166 691634
rect 394250 691398 394486 691634
rect 394570 691398 394806 691634
rect 413930 691718 414166 691954
rect 414250 691718 414486 691954
rect 414570 691718 414806 691954
rect 413930 691398 414166 691634
rect 414250 691398 414486 691634
rect 414570 691398 414806 691634
rect 433930 691718 434166 691954
rect 434250 691718 434486 691954
rect 434570 691718 434806 691954
rect 433930 691398 434166 691634
rect 434250 691398 434486 691634
rect 434570 691398 434806 691634
rect 453930 691718 454166 691954
rect 454250 691718 454486 691954
rect 454570 691718 454806 691954
rect 453930 691398 454166 691634
rect 454250 691398 454486 691634
rect 454570 691398 454806 691634
rect 473930 691718 474166 691954
rect 474250 691718 474486 691954
rect 474570 691718 474806 691954
rect 473930 691398 474166 691634
rect 474250 691398 474486 691634
rect 474570 691398 474806 691634
rect 493930 691718 494166 691954
rect 494250 691718 494486 691954
rect 494570 691718 494806 691954
rect 493930 691398 494166 691634
rect 494250 691398 494486 691634
rect 494570 691398 494806 691634
rect 513930 691718 514166 691954
rect 514250 691718 514486 691954
rect 514570 691718 514806 691954
rect 513930 691398 514166 691634
rect 514250 691398 514486 691634
rect 514570 691398 514806 691634
rect 533930 691718 534166 691954
rect 534250 691718 534486 691954
rect 534570 691718 534806 691954
rect 533930 691398 534166 691634
rect 534250 691398 534486 691634
rect 534570 691398 534806 691634
rect 553930 691718 554166 691954
rect 554250 691718 554486 691954
rect 554570 691718 554806 691954
rect 553930 691398 554166 691634
rect 554250 691398 554486 691634
rect 554570 691398 554806 691634
rect 303930 687218 304166 687454
rect 304250 687218 304486 687454
rect 304570 687218 304806 687454
rect 303930 686898 304166 687134
rect 304250 686898 304486 687134
rect 304570 686898 304806 687134
rect 323930 687218 324166 687454
rect 324250 687218 324486 687454
rect 324570 687218 324806 687454
rect 323930 686898 324166 687134
rect 324250 686898 324486 687134
rect 324570 686898 324806 687134
rect 343930 687218 344166 687454
rect 344250 687218 344486 687454
rect 344570 687218 344806 687454
rect 343930 686898 344166 687134
rect 344250 686898 344486 687134
rect 344570 686898 344806 687134
rect 363930 687218 364166 687454
rect 364250 687218 364486 687454
rect 364570 687218 364806 687454
rect 363930 686898 364166 687134
rect 364250 686898 364486 687134
rect 364570 686898 364806 687134
rect 383930 687218 384166 687454
rect 384250 687218 384486 687454
rect 384570 687218 384806 687454
rect 383930 686898 384166 687134
rect 384250 686898 384486 687134
rect 384570 686898 384806 687134
rect 403930 687218 404166 687454
rect 404250 687218 404486 687454
rect 404570 687218 404806 687454
rect 403930 686898 404166 687134
rect 404250 686898 404486 687134
rect 404570 686898 404806 687134
rect 423930 687218 424166 687454
rect 424250 687218 424486 687454
rect 424570 687218 424806 687454
rect 423930 686898 424166 687134
rect 424250 686898 424486 687134
rect 424570 686898 424806 687134
rect 443930 687218 444166 687454
rect 444250 687218 444486 687454
rect 444570 687218 444806 687454
rect 443930 686898 444166 687134
rect 444250 686898 444486 687134
rect 444570 686898 444806 687134
rect 463930 687218 464166 687454
rect 464250 687218 464486 687454
rect 464570 687218 464806 687454
rect 463930 686898 464166 687134
rect 464250 686898 464486 687134
rect 464570 686898 464806 687134
rect 483930 687218 484166 687454
rect 484250 687218 484486 687454
rect 484570 687218 484806 687454
rect 483930 686898 484166 687134
rect 484250 686898 484486 687134
rect 484570 686898 484806 687134
rect 503930 687218 504166 687454
rect 504250 687218 504486 687454
rect 504570 687218 504806 687454
rect 503930 686898 504166 687134
rect 504250 686898 504486 687134
rect 504570 686898 504806 687134
rect 523930 687218 524166 687454
rect 524250 687218 524486 687454
rect 524570 687218 524806 687454
rect 523930 686898 524166 687134
rect 524250 686898 524486 687134
rect 524570 686898 524806 687134
rect 543930 687218 544166 687454
rect 544250 687218 544486 687454
rect 544570 687218 544806 687454
rect 543930 686898 544166 687134
rect 544250 686898 544486 687134
rect 544570 686898 544806 687134
rect 563930 687218 564166 687454
rect 564250 687218 564486 687454
rect 564570 687218 564806 687454
rect 563930 686898 564166 687134
rect 564250 686898 564486 687134
rect 564570 686898 564806 687134
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 313930 655718 314166 655954
rect 314250 655718 314486 655954
rect 314570 655718 314806 655954
rect 313930 655398 314166 655634
rect 314250 655398 314486 655634
rect 314570 655398 314806 655634
rect 333930 655718 334166 655954
rect 334250 655718 334486 655954
rect 334570 655718 334806 655954
rect 333930 655398 334166 655634
rect 334250 655398 334486 655634
rect 334570 655398 334806 655634
rect 353930 655718 354166 655954
rect 354250 655718 354486 655954
rect 354570 655718 354806 655954
rect 353930 655398 354166 655634
rect 354250 655398 354486 655634
rect 354570 655398 354806 655634
rect 373930 655718 374166 655954
rect 374250 655718 374486 655954
rect 374570 655718 374806 655954
rect 373930 655398 374166 655634
rect 374250 655398 374486 655634
rect 374570 655398 374806 655634
rect 393930 655718 394166 655954
rect 394250 655718 394486 655954
rect 394570 655718 394806 655954
rect 393930 655398 394166 655634
rect 394250 655398 394486 655634
rect 394570 655398 394806 655634
rect 413930 655718 414166 655954
rect 414250 655718 414486 655954
rect 414570 655718 414806 655954
rect 413930 655398 414166 655634
rect 414250 655398 414486 655634
rect 414570 655398 414806 655634
rect 433930 655718 434166 655954
rect 434250 655718 434486 655954
rect 434570 655718 434806 655954
rect 433930 655398 434166 655634
rect 434250 655398 434486 655634
rect 434570 655398 434806 655634
rect 453930 655718 454166 655954
rect 454250 655718 454486 655954
rect 454570 655718 454806 655954
rect 453930 655398 454166 655634
rect 454250 655398 454486 655634
rect 454570 655398 454806 655634
rect 473930 655718 474166 655954
rect 474250 655718 474486 655954
rect 474570 655718 474806 655954
rect 473930 655398 474166 655634
rect 474250 655398 474486 655634
rect 474570 655398 474806 655634
rect 493930 655718 494166 655954
rect 494250 655718 494486 655954
rect 494570 655718 494806 655954
rect 493930 655398 494166 655634
rect 494250 655398 494486 655634
rect 494570 655398 494806 655634
rect 513930 655718 514166 655954
rect 514250 655718 514486 655954
rect 514570 655718 514806 655954
rect 513930 655398 514166 655634
rect 514250 655398 514486 655634
rect 514570 655398 514806 655634
rect 533930 655718 534166 655954
rect 534250 655718 534486 655954
rect 534570 655718 534806 655954
rect 533930 655398 534166 655634
rect 534250 655398 534486 655634
rect 534570 655398 534806 655634
rect 553930 655718 554166 655954
rect 554250 655718 554486 655954
rect 554570 655718 554806 655954
rect 553930 655398 554166 655634
rect 554250 655398 554486 655634
rect 554570 655398 554806 655634
rect 303930 651218 304166 651454
rect 304250 651218 304486 651454
rect 304570 651218 304806 651454
rect 303930 650898 304166 651134
rect 304250 650898 304486 651134
rect 304570 650898 304806 651134
rect 323930 651218 324166 651454
rect 324250 651218 324486 651454
rect 324570 651218 324806 651454
rect 323930 650898 324166 651134
rect 324250 650898 324486 651134
rect 324570 650898 324806 651134
rect 343930 651218 344166 651454
rect 344250 651218 344486 651454
rect 344570 651218 344806 651454
rect 343930 650898 344166 651134
rect 344250 650898 344486 651134
rect 344570 650898 344806 651134
rect 363930 651218 364166 651454
rect 364250 651218 364486 651454
rect 364570 651218 364806 651454
rect 363930 650898 364166 651134
rect 364250 650898 364486 651134
rect 364570 650898 364806 651134
rect 383930 651218 384166 651454
rect 384250 651218 384486 651454
rect 384570 651218 384806 651454
rect 383930 650898 384166 651134
rect 384250 650898 384486 651134
rect 384570 650898 384806 651134
rect 403930 651218 404166 651454
rect 404250 651218 404486 651454
rect 404570 651218 404806 651454
rect 403930 650898 404166 651134
rect 404250 650898 404486 651134
rect 404570 650898 404806 651134
rect 423930 651218 424166 651454
rect 424250 651218 424486 651454
rect 424570 651218 424806 651454
rect 423930 650898 424166 651134
rect 424250 650898 424486 651134
rect 424570 650898 424806 651134
rect 443930 651218 444166 651454
rect 444250 651218 444486 651454
rect 444570 651218 444806 651454
rect 443930 650898 444166 651134
rect 444250 650898 444486 651134
rect 444570 650898 444806 651134
rect 463930 651218 464166 651454
rect 464250 651218 464486 651454
rect 464570 651218 464806 651454
rect 463930 650898 464166 651134
rect 464250 650898 464486 651134
rect 464570 650898 464806 651134
rect 483930 651218 484166 651454
rect 484250 651218 484486 651454
rect 484570 651218 484806 651454
rect 483930 650898 484166 651134
rect 484250 650898 484486 651134
rect 484570 650898 484806 651134
rect 503930 651218 504166 651454
rect 504250 651218 504486 651454
rect 504570 651218 504806 651454
rect 503930 650898 504166 651134
rect 504250 650898 504486 651134
rect 504570 650898 504806 651134
rect 523930 651218 524166 651454
rect 524250 651218 524486 651454
rect 524570 651218 524806 651454
rect 523930 650898 524166 651134
rect 524250 650898 524486 651134
rect 524570 650898 524806 651134
rect 543930 651218 544166 651454
rect 544250 651218 544486 651454
rect 544570 651218 544806 651454
rect 543930 650898 544166 651134
rect 544250 650898 544486 651134
rect 544570 650898 544806 651134
rect 563930 651218 564166 651454
rect 564250 651218 564486 651454
rect 564570 651218 564806 651454
rect 563930 650898 564166 651134
rect 564250 650898 564486 651134
rect 564570 650898 564806 651134
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 313930 619718 314166 619954
rect 314250 619718 314486 619954
rect 314570 619718 314806 619954
rect 313930 619398 314166 619634
rect 314250 619398 314486 619634
rect 314570 619398 314806 619634
rect 333930 619718 334166 619954
rect 334250 619718 334486 619954
rect 334570 619718 334806 619954
rect 333930 619398 334166 619634
rect 334250 619398 334486 619634
rect 334570 619398 334806 619634
rect 353930 619718 354166 619954
rect 354250 619718 354486 619954
rect 354570 619718 354806 619954
rect 353930 619398 354166 619634
rect 354250 619398 354486 619634
rect 354570 619398 354806 619634
rect 373930 619718 374166 619954
rect 374250 619718 374486 619954
rect 374570 619718 374806 619954
rect 373930 619398 374166 619634
rect 374250 619398 374486 619634
rect 374570 619398 374806 619634
rect 393930 619718 394166 619954
rect 394250 619718 394486 619954
rect 394570 619718 394806 619954
rect 393930 619398 394166 619634
rect 394250 619398 394486 619634
rect 394570 619398 394806 619634
rect 413930 619718 414166 619954
rect 414250 619718 414486 619954
rect 414570 619718 414806 619954
rect 413930 619398 414166 619634
rect 414250 619398 414486 619634
rect 414570 619398 414806 619634
rect 433930 619718 434166 619954
rect 434250 619718 434486 619954
rect 434570 619718 434806 619954
rect 433930 619398 434166 619634
rect 434250 619398 434486 619634
rect 434570 619398 434806 619634
rect 453930 619718 454166 619954
rect 454250 619718 454486 619954
rect 454570 619718 454806 619954
rect 453930 619398 454166 619634
rect 454250 619398 454486 619634
rect 454570 619398 454806 619634
rect 473930 619718 474166 619954
rect 474250 619718 474486 619954
rect 474570 619718 474806 619954
rect 473930 619398 474166 619634
rect 474250 619398 474486 619634
rect 474570 619398 474806 619634
rect 493930 619718 494166 619954
rect 494250 619718 494486 619954
rect 494570 619718 494806 619954
rect 493930 619398 494166 619634
rect 494250 619398 494486 619634
rect 494570 619398 494806 619634
rect 513930 619718 514166 619954
rect 514250 619718 514486 619954
rect 514570 619718 514806 619954
rect 513930 619398 514166 619634
rect 514250 619398 514486 619634
rect 514570 619398 514806 619634
rect 533930 619718 534166 619954
rect 534250 619718 534486 619954
rect 534570 619718 534806 619954
rect 533930 619398 534166 619634
rect 534250 619398 534486 619634
rect 534570 619398 534806 619634
rect 553930 619718 554166 619954
rect 554250 619718 554486 619954
rect 554570 619718 554806 619954
rect 553930 619398 554166 619634
rect 554250 619398 554486 619634
rect 554570 619398 554806 619634
rect 303930 615218 304166 615454
rect 304250 615218 304486 615454
rect 304570 615218 304806 615454
rect 303930 614898 304166 615134
rect 304250 614898 304486 615134
rect 304570 614898 304806 615134
rect 323930 615218 324166 615454
rect 324250 615218 324486 615454
rect 324570 615218 324806 615454
rect 323930 614898 324166 615134
rect 324250 614898 324486 615134
rect 324570 614898 324806 615134
rect 343930 615218 344166 615454
rect 344250 615218 344486 615454
rect 344570 615218 344806 615454
rect 343930 614898 344166 615134
rect 344250 614898 344486 615134
rect 344570 614898 344806 615134
rect 363930 615218 364166 615454
rect 364250 615218 364486 615454
rect 364570 615218 364806 615454
rect 363930 614898 364166 615134
rect 364250 614898 364486 615134
rect 364570 614898 364806 615134
rect 383930 615218 384166 615454
rect 384250 615218 384486 615454
rect 384570 615218 384806 615454
rect 383930 614898 384166 615134
rect 384250 614898 384486 615134
rect 384570 614898 384806 615134
rect 403930 615218 404166 615454
rect 404250 615218 404486 615454
rect 404570 615218 404806 615454
rect 403930 614898 404166 615134
rect 404250 614898 404486 615134
rect 404570 614898 404806 615134
rect 423930 615218 424166 615454
rect 424250 615218 424486 615454
rect 424570 615218 424806 615454
rect 423930 614898 424166 615134
rect 424250 614898 424486 615134
rect 424570 614898 424806 615134
rect 443930 615218 444166 615454
rect 444250 615218 444486 615454
rect 444570 615218 444806 615454
rect 443930 614898 444166 615134
rect 444250 614898 444486 615134
rect 444570 614898 444806 615134
rect 463930 615218 464166 615454
rect 464250 615218 464486 615454
rect 464570 615218 464806 615454
rect 463930 614898 464166 615134
rect 464250 614898 464486 615134
rect 464570 614898 464806 615134
rect 483930 615218 484166 615454
rect 484250 615218 484486 615454
rect 484570 615218 484806 615454
rect 483930 614898 484166 615134
rect 484250 614898 484486 615134
rect 484570 614898 484806 615134
rect 503930 615218 504166 615454
rect 504250 615218 504486 615454
rect 504570 615218 504806 615454
rect 503930 614898 504166 615134
rect 504250 614898 504486 615134
rect 504570 614898 504806 615134
rect 523930 615218 524166 615454
rect 524250 615218 524486 615454
rect 524570 615218 524806 615454
rect 523930 614898 524166 615134
rect 524250 614898 524486 615134
rect 524570 614898 524806 615134
rect 543930 615218 544166 615454
rect 544250 615218 544486 615454
rect 544570 615218 544806 615454
rect 543930 614898 544166 615134
rect 544250 614898 544486 615134
rect 544570 614898 544806 615134
rect 563930 615218 564166 615454
rect 564250 615218 564486 615454
rect 564570 615218 564806 615454
rect 563930 614898 564166 615134
rect 564250 614898 564486 615134
rect 564570 614898 564806 615134
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 313930 547718 314166 547954
rect 314250 547718 314486 547954
rect 314570 547718 314806 547954
rect 313930 547398 314166 547634
rect 314250 547398 314486 547634
rect 314570 547398 314806 547634
rect 333930 547718 334166 547954
rect 334250 547718 334486 547954
rect 334570 547718 334806 547954
rect 333930 547398 334166 547634
rect 334250 547398 334486 547634
rect 334570 547398 334806 547634
rect 353930 547718 354166 547954
rect 354250 547718 354486 547954
rect 354570 547718 354806 547954
rect 353930 547398 354166 547634
rect 354250 547398 354486 547634
rect 354570 547398 354806 547634
rect 373930 547718 374166 547954
rect 374250 547718 374486 547954
rect 374570 547718 374806 547954
rect 373930 547398 374166 547634
rect 374250 547398 374486 547634
rect 374570 547398 374806 547634
rect 393930 547718 394166 547954
rect 394250 547718 394486 547954
rect 394570 547718 394806 547954
rect 393930 547398 394166 547634
rect 394250 547398 394486 547634
rect 394570 547398 394806 547634
rect 413930 547718 414166 547954
rect 414250 547718 414486 547954
rect 414570 547718 414806 547954
rect 413930 547398 414166 547634
rect 414250 547398 414486 547634
rect 414570 547398 414806 547634
rect 433930 547718 434166 547954
rect 434250 547718 434486 547954
rect 434570 547718 434806 547954
rect 433930 547398 434166 547634
rect 434250 547398 434486 547634
rect 434570 547398 434806 547634
rect 453930 547718 454166 547954
rect 454250 547718 454486 547954
rect 454570 547718 454806 547954
rect 453930 547398 454166 547634
rect 454250 547398 454486 547634
rect 454570 547398 454806 547634
rect 473930 547718 474166 547954
rect 474250 547718 474486 547954
rect 474570 547718 474806 547954
rect 473930 547398 474166 547634
rect 474250 547398 474486 547634
rect 474570 547398 474806 547634
rect 493930 547718 494166 547954
rect 494250 547718 494486 547954
rect 494570 547718 494806 547954
rect 493930 547398 494166 547634
rect 494250 547398 494486 547634
rect 494570 547398 494806 547634
rect 513930 547718 514166 547954
rect 514250 547718 514486 547954
rect 514570 547718 514806 547954
rect 513930 547398 514166 547634
rect 514250 547398 514486 547634
rect 514570 547398 514806 547634
rect 533930 547718 534166 547954
rect 534250 547718 534486 547954
rect 534570 547718 534806 547954
rect 533930 547398 534166 547634
rect 534250 547398 534486 547634
rect 534570 547398 534806 547634
rect 553930 547718 554166 547954
rect 554250 547718 554486 547954
rect 554570 547718 554806 547954
rect 553930 547398 554166 547634
rect 554250 547398 554486 547634
rect 554570 547398 554806 547634
rect 303930 543218 304166 543454
rect 304250 543218 304486 543454
rect 304570 543218 304806 543454
rect 303930 542898 304166 543134
rect 304250 542898 304486 543134
rect 304570 542898 304806 543134
rect 323930 543218 324166 543454
rect 324250 543218 324486 543454
rect 324570 543218 324806 543454
rect 323930 542898 324166 543134
rect 324250 542898 324486 543134
rect 324570 542898 324806 543134
rect 343930 543218 344166 543454
rect 344250 543218 344486 543454
rect 344570 543218 344806 543454
rect 343930 542898 344166 543134
rect 344250 542898 344486 543134
rect 344570 542898 344806 543134
rect 363930 543218 364166 543454
rect 364250 543218 364486 543454
rect 364570 543218 364806 543454
rect 363930 542898 364166 543134
rect 364250 542898 364486 543134
rect 364570 542898 364806 543134
rect 383930 543218 384166 543454
rect 384250 543218 384486 543454
rect 384570 543218 384806 543454
rect 383930 542898 384166 543134
rect 384250 542898 384486 543134
rect 384570 542898 384806 543134
rect 403930 543218 404166 543454
rect 404250 543218 404486 543454
rect 404570 543218 404806 543454
rect 403930 542898 404166 543134
rect 404250 542898 404486 543134
rect 404570 542898 404806 543134
rect 423930 543218 424166 543454
rect 424250 543218 424486 543454
rect 424570 543218 424806 543454
rect 423930 542898 424166 543134
rect 424250 542898 424486 543134
rect 424570 542898 424806 543134
rect 443930 543218 444166 543454
rect 444250 543218 444486 543454
rect 444570 543218 444806 543454
rect 443930 542898 444166 543134
rect 444250 542898 444486 543134
rect 444570 542898 444806 543134
rect 463930 543218 464166 543454
rect 464250 543218 464486 543454
rect 464570 543218 464806 543454
rect 463930 542898 464166 543134
rect 464250 542898 464486 543134
rect 464570 542898 464806 543134
rect 483930 543218 484166 543454
rect 484250 543218 484486 543454
rect 484570 543218 484806 543454
rect 483930 542898 484166 543134
rect 484250 542898 484486 543134
rect 484570 542898 484806 543134
rect 503930 543218 504166 543454
rect 504250 543218 504486 543454
rect 504570 543218 504806 543454
rect 503930 542898 504166 543134
rect 504250 542898 504486 543134
rect 504570 542898 504806 543134
rect 523930 543218 524166 543454
rect 524250 543218 524486 543454
rect 524570 543218 524806 543454
rect 523930 542898 524166 543134
rect 524250 542898 524486 543134
rect 524570 542898 524806 543134
rect 543930 543218 544166 543454
rect 544250 543218 544486 543454
rect 544570 543218 544806 543454
rect 543930 542898 544166 543134
rect 544250 542898 544486 543134
rect 544570 542898 544806 543134
rect 563930 543218 564166 543454
rect 564250 543218 564486 543454
rect 564570 543218 564806 543454
rect 563930 542898 564166 543134
rect 564250 542898 564486 543134
rect 564570 542898 564806 543134
rect 313930 511718 314166 511954
rect 314250 511718 314486 511954
rect 314570 511718 314806 511954
rect 313930 511398 314166 511634
rect 314250 511398 314486 511634
rect 314570 511398 314806 511634
rect 333930 511718 334166 511954
rect 334250 511718 334486 511954
rect 334570 511718 334806 511954
rect 333930 511398 334166 511634
rect 334250 511398 334486 511634
rect 334570 511398 334806 511634
rect 353930 511718 354166 511954
rect 354250 511718 354486 511954
rect 354570 511718 354806 511954
rect 353930 511398 354166 511634
rect 354250 511398 354486 511634
rect 354570 511398 354806 511634
rect 373930 511718 374166 511954
rect 374250 511718 374486 511954
rect 374570 511718 374806 511954
rect 373930 511398 374166 511634
rect 374250 511398 374486 511634
rect 374570 511398 374806 511634
rect 393930 511718 394166 511954
rect 394250 511718 394486 511954
rect 394570 511718 394806 511954
rect 393930 511398 394166 511634
rect 394250 511398 394486 511634
rect 394570 511398 394806 511634
rect 413930 511718 414166 511954
rect 414250 511718 414486 511954
rect 414570 511718 414806 511954
rect 413930 511398 414166 511634
rect 414250 511398 414486 511634
rect 414570 511398 414806 511634
rect 433930 511718 434166 511954
rect 434250 511718 434486 511954
rect 434570 511718 434806 511954
rect 433930 511398 434166 511634
rect 434250 511398 434486 511634
rect 434570 511398 434806 511634
rect 453930 511718 454166 511954
rect 454250 511718 454486 511954
rect 454570 511718 454806 511954
rect 453930 511398 454166 511634
rect 454250 511398 454486 511634
rect 454570 511398 454806 511634
rect 473930 511718 474166 511954
rect 474250 511718 474486 511954
rect 474570 511718 474806 511954
rect 473930 511398 474166 511634
rect 474250 511398 474486 511634
rect 474570 511398 474806 511634
rect 493930 511718 494166 511954
rect 494250 511718 494486 511954
rect 494570 511718 494806 511954
rect 493930 511398 494166 511634
rect 494250 511398 494486 511634
rect 494570 511398 494806 511634
rect 513930 511718 514166 511954
rect 514250 511718 514486 511954
rect 514570 511718 514806 511954
rect 513930 511398 514166 511634
rect 514250 511398 514486 511634
rect 514570 511398 514806 511634
rect 533930 511718 534166 511954
rect 534250 511718 534486 511954
rect 534570 511718 534806 511954
rect 533930 511398 534166 511634
rect 534250 511398 534486 511634
rect 534570 511398 534806 511634
rect 553930 511718 554166 511954
rect 554250 511718 554486 511954
rect 554570 511718 554806 511954
rect 553930 511398 554166 511634
rect 554250 511398 554486 511634
rect 554570 511398 554806 511634
rect 303930 507218 304166 507454
rect 304250 507218 304486 507454
rect 304570 507218 304806 507454
rect 303930 506898 304166 507134
rect 304250 506898 304486 507134
rect 304570 506898 304806 507134
rect 323930 507218 324166 507454
rect 324250 507218 324486 507454
rect 324570 507218 324806 507454
rect 323930 506898 324166 507134
rect 324250 506898 324486 507134
rect 324570 506898 324806 507134
rect 343930 507218 344166 507454
rect 344250 507218 344486 507454
rect 344570 507218 344806 507454
rect 343930 506898 344166 507134
rect 344250 506898 344486 507134
rect 344570 506898 344806 507134
rect 363930 507218 364166 507454
rect 364250 507218 364486 507454
rect 364570 507218 364806 507454
rect 363930 506898 364166 507134
rect 364250 506898 364486 507134
rect 364570 506898 364806 507134
rect 383930 507218 384166 507454
rect 384250 507218 384486 507454
rect 384570 507218 384806 507454
rect 383930 506898 384166 507134
rect 384250 506898 384486 507134
rect 384570 506898 384806 507134
rect 403930 507218 404166 507454
rect 404250 507218 404486 507454
rect 404570 507218 404806 507454
rect 403930 506898 404166 507134
rect 404250 506898 404486 507134
rect 404570 506898 404806 507134
rect 423930 507218 424166 507454
rect 424250 507218 424486 507454
rect 424570 507218 424806 507454
rect 423930 506898 424166 507134
rect 424250 506898 424486 507134
rect 424570 506898 424806 507134
rect 443930 507218 444166 507454
rect 444250 507218 444486 507454
rect 444570 507218 444806 507454
rect 443930 506898 444166 507134
rect 444250 506898 444486 507134
rect 444570 506898 444806 507134
rect 463930 507218 464166 507454
rect 464250 507218 464486 507454
rect 464570 507218 464806 507454
rect 463930 506898 464166 507134
rect 464250 506898 464486 507134
rect 464570 506898 464806 507134
rect 483930 507218 484166 507454
rect 484250 507218 484486 507454
rect 484570 507218 484806 507454
rect 483930 506898 484166 507134
rect 484250 506898 484486 507134
rect 484570 506898 484806 507134
rect 503930 507218 504166 507454
rect 504250 507218 504486 507454
rect 504570 507218 504806 507454
rect 503930 506898 504166 507134
rect 504250 506898 504486 507134
rect 504570 506898 504806 507134
rect 523930 507218 524166 507454
rect 524250 507218 524486 507454
rect 524570 507218 524806 507454
rect 523930 506898 524166 507134
rect 524250 506898 524486 507134
rect 524570 506898 524806 507134
rect 543930 507218 544166 507454
rect 544250 507218 544486 507454
rect 544570 507218 544806 507454
rect 543930 506898 544166 507134
rect 544250 506898 544486 507134
rect 544570 506898 544806 507134
rect 563930 507218 564166 507454
rect 564250 507218 564486 507454
rect 564570 507218 564806 507454
rect 563930 506898 564166 507134
rect 564250 506898 564486 507134
rect 564570 506898 564806 507134
rect 313930 475718 314166 475954
rect 314250 475718 314486 475954
rect 314570 475718 314806 475954
rect 313930 475398 314166 475634
rect 314250 475398 314486 475634
rect 314570 475398 314806 475634
rect 333930 475718 334166 475954
rect 334250 475718 334486 475954
rect 334570 475718 334806 475954
rect 333930 475398 334166 475634
rect 334250 475398 334486 475634
rect 334570 475398 334806 475634
rect 353930 475718 354166 475954
rect 354250 475718 354486 475954
rect 354570 475718 354806 475954
rect 353930 475398 354166 475634
rect 354250 475398 354486 475634
rect 354570 475398 354806 475634
rect 373930 475718 374166 475954
rect 374250 475718 374486 475954
rect 374570 475718 374806 475954
rect 373930 475398 374166 475634
rect 374250 475398 374486 475634
rect 374570 475398 374806 475634
rect 393930 475718 394166 475954
rect 394250 475718 394486 475954
rect 394570 475718 394806 475954
rect 393930 475398 394166 475634
rect 394250 475398 394486 475634
rect 394570 475398 394806 475634
rect 413930 475718 414166 475954
rect 414250 475718 414486 475954
rect 414570 475718 414806 475954
rect 413930 475398 414166 475634
rect 414250 475398 414486 475634
rect 414570 475398 414806 475634
rect 433930 475718 434166 475954
rect 434250 475718 434486 475954
rect 434570 475718 434806 475954
rect 433930 475398 434166 475634
rect 434250 475398 434486 475634
rect 434570 475398 434806 475634
rect 453930 475718 454166 475954
rect 454250 475718 454486 475954
rect 454570 475718 454806 475954
rect 453930 475398 454166 475634
rect 454250 475398 454486 475634
rect 454570 475398 454806 475634
rect 473930 475718 474166 475954
rect 474250 475718 474486 475954
rect 474570 475718 474806 475954
rect 473930 475398 474166 475634
rect 474250 475398 474486 475634
rect 474570 475398 474806 475634
rect 493930 475718 494166 475954
rect 494250 475718 494486 475954
rect 494570 475718 494806 475954
rect 493930 475398 494166 475634
rect 494250 475398 494486 475634
rect 494570 475398 494806 475634
rect 513930 475718 514166 475954
rect 514250 475718 514486 475954
rect 514570 475718 514806 475954
rect 513930 475398 514166 475634
rect 514250 475398 514486 475634
rect 514570 475398 514806 475634
rect 533930 475718 534166 475954
rect 534250 475718 534486 475954
rect 534570 475718 534806 475954
rect 533930 475398 534166 475634
rect 534250 475398 534486 475634
rect 534570 475398 534806 475634
rect 553930 475718 554166 475954
rect 554250 475718 554486 475954
rect 554570 475718 554806 475954
rect 553930 475398 554166 475634
rect 554250 475398 554486 475634
rect 554570 475398 554806 475634
rect 303930 471218 304166 471454
rect 304250 471218 304486 471454
rect 304570 471218 304806 471454
rect 303930 470898 304166 471134
rect 304250 470898 304486 471134
rect 304570 470898 304806 471134
rect 323930 471218 324166 471454
rect 324250 471218 324486 471454
rect 324570 471218 324806 471454
rect 323930 470898 324166 471134
rect 324250 470898 324486 471134
rect 324570 470898 324806 471134
rect 343930 471218 344166 471454
rect 344250 471218 344486 471454
rect 344570 471218 344806 471454
rect 343930 470898 344166 471134
rect 344250 470898 344486 471134
rect 344570 470898 344806 471134
rect 363930 471218 364166 471454
rect 364250 471218 364486 471454
rect 364570 471218 364806 471454
rect 363930 470898 364166 471134
rect 364250 470898 364486 471134
rect 364570 470898 364806 471134
rect 383930 471218 384166 471454
rect 384250 471218 384486 471454
rect 384570 471218 384806 471454
rect 383930 470898 384166 471134
rect 384250 470898 384486 471134
rect 384570 470898 384806 471134
rect 403930 471218 404166 471454
rect 404250 471218 404486 471454
rect 404570 471218 404806 471454
rect 403930 470898 404166 471134
rect 404250 470898 404486 471134
rect 404570 470898 404806 471134
rect 423930 471218 424166 471454
rect 424250 471218 424486 471454
rect 424570 471218 424806 471454
rect 423930 470898 424166 471134
rect 424250 470898 424486 471134
rect 424570 470898 424806 471134
rect 443930 471218 444166 471454
rect 444250 471218 444486 471454
rect 444570 471218 444806 471454
rect 443930 470898 444166 471134
rect 444250 470898 444486 471134
rect 444570 470898 444806 471134
rect 463930 471218 464166 471454
rect 464250 471218 464486 471454
rect 464570 471218 464806 471454
rect 463930 470898 464166 471134
rect 464250 470898 464486 471134
rect 464570 470898 464806 471134
rect 483930 471218 484166 471454
rect 484250 471218 484486 471454
rect 484570 471218 484806 471454
rect 483930 470898 484166 471134
rect 484250 470898 484486 471134
rect 484570 470898 484806 471134
rect 503930 471218 504166 471454
rect 504250 471218 504486 471454
rect 504570 471218 504806 471454
rect 503930 470898 504166 471134
rect 504250 470898 504486 471134
rect 504570 470898 504806 471134
rect 523930 471218 524166 471454
rect 524250 471218 524486 471454
rect 524570 471218 524806 471454
rect 523930 470898 524166 471134
rect 524250 470898 524486 471134
rect 524570 470898 524806 471134
rect 543930 471218 544166 471454
rect 544250 471218 544486 471454
rect 544570 471218 544806 471454
rect 543930 470898 544166 471134
rect 544250 470898 544486 471134
rect 544570 470898 544806 471134
rect 563930 471218 564166 471454
rect 564250 471218 564486 471454
rect 564570 471218 564806 471454
rect 563930 470898 564166 471134
rect 564250 470898 564486 471134
rect 564570 470898 564806 471134
rect 313930 439718 314166 439954
rect 314250 439718 314486 439954
rect 314570 439718 314806 439954
rect 313930 439398 314166 439634
rect 314250 439398 314486 439634
rect 314570 439398 314806 439634
rect 333930 439718 334166 439954
rect 334250 439718 334486 439954
rect 334570 439718 334806 439954
rect 333930 439398 334166 439634
rect 334250 439398 334486 439634
rect 334570 439398 334806 439634
rect 353930 439718 354166 439954
rect 354250 439718 354486 439954
rect 354570 439718 354806 439954
rect 353930 439398 354166 439634
rect 354250 439398 354486 439634
rect 354570 439398 354806 439634
rect 373930 439718 374166 439954
rect 374250 439718 374486 439954
rect 374570 439718 374806 439954
rect 373930 439398 374166 439634
rect 374250 439398 374486 439634
rect 374570 439398 374806 439634
rect 393930 439718 394166 439954
rect 394250 439718 394486 439954
rect 394570 439718 394806 439954
rect 393930 439398 394166 439634
rect 394250 439398 394486 439634
rect 394570 439398 394806 439634
rect 413930 439718 414166 439954
rect 414250 439718 414486 439954
rect 414570 439718 414806 439954
rect 413930 439398 414166 439634
rect 414250 439398 414486 439634
rect 414570 439398 414806 439634
rect 433930 439718 434166 439954
rect 434250 439718 434486 439954
rect 434570 439718 434806 439954
rect 433930 439398 434166 439634
rect 434250 439398 434486 439634
rect 434570 439398 434806 439634
rect 453930 439718 454166 439954
rect 454250 439718 454486 439954
rect 454570 439718 454806 439954
rect 453930 439398 454166 439634
rect 454250 439398 454486 439634
rect 454570 439398 454806 439634
rect 473930 439718 474166 439954
rect 474250 439718 474486 439954
rect 474570 439718 474806 439954
rect 473930 439398 474166 439634
rect 474250 439398 474486 439634
rect 474570 439398 474806 439634
rect 493930 439718 494166 439954
rect 494250 439718 494486 439954
rect 494570 439718 494806 439954
rect 493930 439398 494166 439634
rect 494250 439398 494486 439634
rect 494570 439398 494806 439634
rect 513930 439718 514166 439954
rect 514250 439718 514486 439954
rect 514570 439718 514806 439954
rect 513930 439398 514166 439634
rect 514250 439398 514486 439634
rect 514570 439398 514806 439634
rect 533930 439718 534166 439954
rect 534250 439718 534486 439954
rect 534570 439718 534806 439954
rect 533930 439398 534166 439634
rect 534250 439398 534486 439634
rect 534570 439398 534806 439634
rect 553930 439718 554166 439954
rect 554250 439718 554486 439954
rect 554570 439718 554806 439954
rect 553930 439398 554166 439634
rect 554250 439398 554486 439634
rect 554570 439398 554806 439634
rect 303930 435218 304166 435454
rect 304250 435218 304486 435454
rect 304570 435218 304806 435454
rect 303930 434898 304166 435134
rect 304250 434898 304486 435134
rect 304570 434898 304806 435134
rect 323930 435218 324166 435454
rect 324250 435218 324486 435454
rect 324570 435218 324806 435454
rect 323930 434898 324166 435134
rect 324250 434898 324486 435134
rect 324570 434898 324806 435134
rect 343930 435218 344166 435454
rect 344250 435218 344486 435454
rect 344570 435218 344806 435454
rect 343930 434898 344166 435134
rect 344250 434898 344486 435134
rect 344570 434898 344806 435134
rect 363930 435218 364166 435454
rect 364250 435218 364486 435454
rect 364570 435218 364806 435454
rect 363930 434898 364166 435134
rect 364250 434898 364486 435134
rect 364570 434898 364806 435134
rect 383930 435218 384166 435454
rect 384250 435218 384486 435454
rect 384570 435218 384806 435454
rect 383930 434898 384166 435134
rect 384250 434898 384486 435134
rect 384570 434898 384806 435134
rect 403930 435218 404166 435454
rect 404250 435218 404486 435454
rect 404570 435218 404806 435454
rect 403930 434898 404166 435134
rect 404250 434898 404486 435134
rect 404570 434898 404806 435134
rect 423930 435218 424166 435454
rect 424250 435218 424486 435454
rect 424570 435218 424806 435454
rect 423930 434898 424166 435134
rect 424250 434898 424486 435134
rect 424570 434898 424806 435134
rect 443930 435218 444166 435454
rect 444250 435218 444486 435454
rect 444570 435218 444806 435454
rect 443930 434898 444166 435134
rect 444250 434898 444486 435134
rect 444570 434898 444806 435134
rect 463930 435218 464166 435454
rect 464250 435218 464486 435454
rect 464570 435218 464806 435454
rect 463930 434898 464166 435134
rect 464250 434898 464486 435134
rect 464570 434898 464806 435134
rect 483930 435218 484166 435454
rect 484250 435218 484486 435454
rect 484570 435218 484806 435454
rect 483930 434898 484166 435134
rect 484250 434898 484486 435134
rect 484570 434898 484806 435134
rect 503930 435218 504166 435454
rect 504250 435218 504486 435454
rect 504570 435218 504806 435454
rect 503930 434898 504166 435134
rect 504250 434898 504486 435134
rect 504570 434898 504806 435134
rect 523930 435218 524166 435454
rect 524250 435218 524486 435454
rect 524570 435218 524806 435454
rect 523930 434898 524166 435134
rect 524250 434898 524486 435134
rect 524570 434898 524806 435134
rect 543930 435218 544166 435454
rect 544250 435218 544486 435454
rect 544570 435218 544806 435454
rect 543930 434898 544166 435134
rect 544250 434898 544486 435134
rect 544570 434898 544806 435134
rect 563930 435218 564166 435454
rect 564250 435218 564486 435454
rect 564570 435218 564806 435454
rect 563930 434898 564166 435134
rect 564250 434898 564486 435134
rect 564570 434898 564806 435134
rect 313930 403718 314166 403954
rect 314250 403718 314486 403954
rect 314570 403718 314806 403954
rect 313930 403398 314166 403634
rect 314250 403398 314486 403634
rect 314570 403398 314806 403634
rect 333930 403718 334166 403954
rect 334250 403718 334486 403954
rect 334570 403718 334806 403954
rect 333930 403398 334166 403634
rect 334250 403398 334486 403634
rect 334570 403398 334806 403634
rect 353930 403718 354166 403954
rect 354250 403718 354486 403954
rect 354570 403718 354806 403954
rect 353930 403398 354166 403634
rect 354250 403398 354486 403634
rect 354570 403398 354806 403634
rect 373930 403718 374166 403954
rect 374250 403718 374486 403954
rect 374570 403718 374806 403954
rect 373930 403398 374166 403634
rect 374250 403398 374486 403634
rect 374570 403398 374806 403634
rect 393930 403718 394166 403954
rect 394250 403718 394486 403954
rect 394570 403718 394806 403954
rect 393930 403398 394166 403634
rect 394250 403398 394486 403634
rect 394570 403398 394806 403634
rect 413930 403718 414166 403954
rect 414250 403718 414486 403954
rect 414570 403718 414806 403954
rect 413930 403398 414166 403634
rect 414250 403398 414486 403634
rect 414570 403398 414806 403634
rect 433930 403718 434166 403954
rect 434250 403718 434486 403954
rect 434570 403718 434806 403954
rect 433930 403398 434166 403634
rect 434250 403398 434486 403634
rect 434570 403398 434806 403634
rect 453930 403718 454166 403954
rect 454250 403718 454486 403954
rect 454570 403718 454806 403954
rect 453930 403398 454166 403634
rect 454250 403398 454486 403634
rect 454570 403398 454806 403634
rect 473930 403718 474166 403954
rect 474250 403718 474486 403954
rect 474570 403718 474806 403954
rect 473930 403398 474166 403634
rect 474250 403398 474486 403634
rect 474570 403398 474806 403634
rect 493930 403718 494166 403954
rect 494250 403718 494486 403954
rect 494570 403718 494806 403954
rect 493930 403398 494166 403634
rect 494250 403398 494486 403634
rect 494570 403398 494806 403634
rect 513930 403718 514166 403954
rect 514250 403718 514486 403954
rect 514570 403718 514806 403954
rect 513930 403398 514166 403634
rect 514250 403398 514486 403634
rect 514570 403398 514806 403634
rect 533930 403718 534166 403954
rect 534250 403718 534486 403954
rect 534570 403718 534806 403954
rect 533930 403398 534166 403634
rect 534250 403398 534486 403634
rect 534570 403398 534806 403634
rect 553930 403718 554166 403954
rect 554250 403718 554486 403954
rect 554570 403718 554806 403954
rect 553930 403398 554166 403634
rect 554250 403398 554486 403634
rect 554570 403398 554806 403634
rect 303930 399218 304166 399454
rect 304250 399218 304486 399454
rect 304570 399218 304806 399454
rect 303930 398898 304166 399134
rect 304250 398898 304486 399134
rect 304570 398898 304806 399134
rect 323930 399218 324166 399454
rect 324250 399218 324486 399454
rect 324570 399218 324806 399454
rect 323930 398898 324166 399134
rect 324250 398898 324486 399134
rect 324570 398898 324806 399134
rect 343930 399218 344166 399454
rect 344250 399218 344486 399454
rect 344570 399218 344806 399454
rect 343930 398898 344166 399134
rect 344250 398898 344486 399134
rect 344570 398898 344806 399134
rect 363930 399218 364166 399454
rect 364250 399218 364486 399454
rect 364570 399218 364806 399454
rect 363930 398898 364166 399134
rect 364250 398898 364486 399134
rect 364570 398898 364806 399134
rect 383930 399218 384166 399454
rect 384250 399218 384486 399454
rect 384570 399218 384806 399454
rect 383930 398898 384166 399134
rect 384250 398898 384486 399134
rect 384570 398898 384806 399134
rect 403930 399218 404166 399454
rect 404250 399218 404486 399454
rect 404570 399218 404806 399454
rect 403930 398898 404166 399134
rect 404250 398898 404486 399134
rect 404570 398898 404806 399134
rect 423930 399218 424166 399454
rect 424250 399218 424486 399454
rect 424570 399218 424806 399454
rect 423930 398898 424166 399134
rect 424250 398898 424486 399134
rect 424570 398898 424806 399134
rect 443930 399218 444166 399454
rect 444250 399218 444486 399454
rect 444570 399218 444806 399454
rect 443930 398898 444166 399134
rect 444250 398898 444486 399134
rect 444570 398898 444806 399134
rect 463930 399218 464166 399454
rect 464250 399218 464486 399454
rect 464570 399218 464806 399454
rect 463930 398898 464166 399134
rect 464250 398898 464486 399134
rect 464570 398898 464806 399134
rect 483930 399218 484166 399454
rect 484250 399218 484486 399454
rect 484570 399218 484806 399454
rect 483930 398898 484166 399134
rect 484250 398898 484486 399134
rect 484570 398898 484806 399134
rect 503930 399218 504166 399454
rect 504250 399218 504486 399454
rect 504570 399218 504806 399454
rect 503930 398898 504166 399134
rect 504250 398898 504486 399134
rect 504570 398898 504806 399134
rect 523930 399218 524166 399454
rect 524250 399218 524486 399454
rect 524570 399218 524806 399454
rect 523930 398898 524166 399134
rect 524250 398898 524486 399134
rect 524570 398898 524806 399134
rect 543930 399218 544166 399454
rect 544250 399218 544486 399454
rect 544570 399218 544806 399454
rect 543930 398898 544166 399134
rect 544250 398898 544486 399134
rect 544570 398898 544806 399134
rect 563930 399218 564166 399454
rect 564250 399218 564486 399454
rect 564570 399218 564806 399454
rect 563930 398898 564166 399134
rect 564250 398898 564486 399134
rect 564570 398898 564806 399134
rect 313930 367718 314166 367954
rect 314250 367718 314486 367954
rect 314570 367718 314806 367954
rect 313930 367398 314166 367634
rect 314250 367398 314486 367634
rect 314570 367398 314806 367634
rect 333930 367718 334166 367954
rect 334250 367718 334486 367954
rect 334570 367718 334806 367954
rect 333930 367398 334166 367634
rect 334250 367398 334486 367634
rect 334570 367398 334806 367634
rect 353930 367718 354166 367954
rect 354250 367718 354486 367954
rect 354570 367718 354806 367954
rect 353930 367398 354166 367634
rect 354250 367398 354486 367634
rect 354570 367398 354806 367634
rect 373930 367718 374166 367954
rect 374250 367718 374486 367954
rect 374570 367718 374806 367954
rect 373930 367398 374166 367634
rect 374250 367398 374486 367634
rect 374570 367398 374806 367634
rect 393930 367718 394166 367954
rect 394250 367718 394486 367954
rect 394570 367718 394806 367954
rect 393930 367398 394166 367634
rect 394250 367398 394486 367634
rect 394570 367398 394806 367634
rect 413930 367718 414166 367954
rect 414250 367718 414486 367954
rect 414570 367718 414806 367954
rect 413930 367398 414166 367634
rect 414250 367398 414486 367634
rect 414570 367398 414806 367634
rect 433930 367718 434166 367954
rect 434250 367718 434486 367954
rect 434570 367718 434806 367954
rect 433930 367398 434166 367634
rect 434250 367398 434486 367634
rect 434570 367398 434806 367634
rect 453930 367718 454166 367954
rect 454250 367718 454486 367954
rect 454570 367718 454806 367954
rect 453930 367398 454166 367634
rect 454250 367398 454486 367634
rect 454570 367398 454806 367634
rect 473930 367718 474166 367954
rect 474250 367718 474486 367954
rect 474570 367718 474806 367954
rect 473930 367398 474166 367634
rect 474250 367398 474486 367634
rect 474570 367398 474806 367634
rect 493930 367718 494166 367954
rect 494250 367718 494486 367954
rect 494570 367718 494806 367954
rect 493930 367398 494166 367634
rect 494250 367398 494486 367634
rect 494570 367398 494806 367634
rect 513930 367718 514166 367954
rect 514250 367718 514486 367954
rect 514570 367718 514806 367954
rect 513930 367398 514166 367634
rect 514250 367398 514486 367634
rect 514570 367398 514806 367634
rect 533930 367718 534166 367954
rect 534250 367718 534486 367954
rect 534570 367718 534806 367954
rect 533930 367398 534166 367634
rect 534250 367398 534486 367634
rect 534570 367398 534806 367634
rect 553930 367718 554166 367954
rect 554250 367718 554486 367954
rect 554570 367718 554806 367954
rect 553930 367398 554166 367634
rect 554250 367398 554486 367634
rect 554570 367398 554806 367634
rect 303930 363218 304166 363454
rect 304250 363218 304486 363454
rect 304570 363218 304806 363454
rect 303930 362898 304166 363134
rect 304250 362898 304486 363134
rect 304570 362898 304806 363134
rect 323930 363218 324166 363454
rect 324250 363218 324486 363454
rect 324570 363218 324806 363454
rect 323930 362898 324166 363134
rect 324250 362898 324486 363134
rect 324570 362898 324806 363134
rect 343930 363218 344166 363454
rect 344250 363218 344486 363454
rect 344570 363218 344806 363454
rect 343930 362898 344166 363134
rect 344250 362898 344486 363134
rect 344570 362898 344806 363134
rect 363930 363218 364166 363454
rect 364250 363218 364486 363454
rect 364570 363218 364806 363454
rect 363930 362898 364166 363134
rect 364250 362898 364486 363134
rect 364570 362898 364806 363134
rect 383930 363218 384166 363454
rect 384250 363218 384486 363454
rect 384570 363218 384806 363454
rect 383930 362898 384166 363134
rect 384250 362898 384486 363134
rect 384570 362898 384806 363134
rect 403930 363218 404166 363454
rect 404250 363218 404486 363454
rect 404570 363218 404806 363454
rect 403930 362898 404166 363134
rect 404250 362898 404486 363134
rect 404570 362898 404806 363134
rect 423930 363218 424166 363454
rect 424250 363218 424486 363454
rect 424570 363218 424806 363454
rect 423930 362898 424166 363134
rect 424250 362898 424486 363134
rect 424570 362898 424806 363134
rect 443930 363218 444166 363454
rect 444250 363218 444486 363454
rect 444570 363218 444806 363454
rect 443930 362898 444166 363134
rect 444250 362898 444486 363134
rect 444570 362898 444806 363134
rect 463930 363218 464166 363454
rect 464250 363218 464486 363454
rect 464570 363218 464806 363454
rect 463930 362898 464166 363134
rect 464250 362898 464486 363134
rect 464570 362898 464806 363134
rect 483930 363218 484166 363454
rect 484250 363218 484486 363454
rect 484570 363218 484806 363454
rect 483930 362898 484166 363134
rect 484250 362898 484486 363134
rect 484570 362898 484806 363134
rect 503930 363218 504166 363454
rect 504250 363218 504486 363454
rect 504570 363218 504806 363454
rect 503930 362898 504166 363134
rect 504250 362898 504486 363134
rect 504570 362898 504806 363134
rect 523930 363218 524166 363454
rect 524250 363218 524486 363454
rect 524570 363218 524806 363454
rect 523930 362898 524166 363134
rect 524250 362898 524486 363134
rect 524570 362898 524806 363134
rect 543930 363218 544166 363454
rect 544250 363218 544486 363454
rect 544570 363218 544806 363454
rect 543930 362898 544166 363134
rect 544250 362898 544486 363134
rect 544570 362898 544806 363134
rect 563930 363218 564166 363454
rect 564250 363218 564486 363454
rect 564570 363218 564806 363454
rect 563930 362898 564166 363134
rect 564250 362898 564486 363134
rect 564570 362898 564806 363134
rect 313930 295718 314166 295954
rect 314250 295718 314486 295954
rect 314570 295718 314806 295954
rect 313930 295398 314166 295634
rect 314250 295398 314486 295634
rect 314570 295398 314806 295634
rect 333930 295718 334166 295954
rect 334250 295718 334486 295954
rect 334570 295718 334806 295954
rect 333930 295398 334166 295634
rect 334250 295398 334486 295634
rect 334570 295398 334806 295634
rect 353930 295718 354166 295954
rect 354250 295718 354486 295954
rect 354570 295718 354806 295954
rect 353930 295398 354166 295634
rect 354250 295398 354486 295634
rect 354570 295398 354806 295634
rect 373930 295718 374166 295954
rect 374250 295718 374486 295954
rect 374570 295718 374806 295954
rect 373930 295398 374166 295634
rect 374250 295398 374486 295634
rect 374570 295398 374806 295634
rect 393930 295718 394166 295954
rect 394250 295718 394486 295954
rect 394570 295718 394806 295954
rect 393930 295398 394166 295634
rect 394250 295398 394486 295634
rect 394570 295398 394806 295634
rect 413930 295718 414166 295954
rect 414250 295718 414486 295954
rect 414570 295718 414806 295954
rect 413930 295398 414166 295634
rect 414250 295398 414486 295634
rect 414570 295398 414806 295634
rect 433930 295718 434166 295954
rect 434250 295718 434486 295954
rect 434570 295718 434806 295954
rect 433930 295398 434166 295634
rect 434250 295398 434486 295634
rect 434570 295398 434806 295634
rect 453930 295718 454166 295954
rect 454250 295718 454486 295954
rect 454570 295718 454806 295954
rect 453930 295398 454166 295634
rect 454250 295398 454486 295634
rect 454570 295398 454806 295634
rect 473930 295718 474166 295954
rect 474250 295718 474486 295954
rect 474570 295718 474806 295954
rect 473930 295398 474166 295634
rect 474250 295398 474486 295634
rect 474570 295398 474806 295634
rect 493930 295718 494166 295954
rect 494250 295718 494486 295954
rect 494570 295718 494806 295954
rect 493930 295398 494166 295634
rect 494250 295398 494486 295634
rect 494570 295398 494806 295634
rect 513930 295718 514166 295954
rect 514250 295718 514486 295954
rect 514570 295718 514806 295954
rect 513930 295398 514166 295634
rect 514250 295398 514486 295634
rect 514570 295398 514806 295634
rect 533930 295718 534166 295954
rect 534250 295718 534486 295954
rect 534570 295718 534806 295954
rect 533930 295398 534166 295634
rect 534250 295398 534486 295634
rect 534570 295398 534806 295634
rect 553930 295718 554166 295954
rect 554250 295718 554486 295954
rect 554570 295718 554806 295954
rect 553930 295398 554166 295634
rect 554250 295398 554486 295634
rect 554570 295398 554806 295634
rect 303930 291218 304166 291454
rect 304250 291218 304486 291454
rect 304570 291218 304806 291454
rect 303930 290898 304166 291134
rect 304250 290898 304486 291134
rect 304570 290898 304806 291134
rect 323930 291218 324166 291454
rect 324250 291218 324486 291454
rect 324570 291218 324806 291454
rect 323930 290898 324166 291134
rect 324250 290898 324486 291134
rect 324570 290898 324806 291134
rect 343930 291218 344166 291454
rect 344250 291218 344486 291454
rect 344570 291218 344806 291454
rect 343930 290898 344166 291134
rect 344250 290898 344486 291134
rect 344570 290898 344806 291134
rect 363930 291218 364166 291454
rect 364250 291218 364486 291454
rect 364570 291218 364806 291454
rect 363930 290898 364166 291134
rect 364250 290898 364486 291134
rect 364570 290898 364806 291134
rect 383930 291218 384166 291454
rect 384250 291218 384486 291454
rect 384570 291218 384806 291454
rect 383930 290898 384166 291134
rect 384250 290898 384486 291134
rect 384570 290898 384806 291134
rect 403930 291218 404166 291454
rect 404250 291218 404486 291454
rect 404570 291218 404806 291454
rect 403930 290898 404166 291134
rect 404250 290898 404486 291134
rect 404570 290898 404806 291134
rect 423930 291218 424166 291454
rect 424250 291218 424486 291454
rect 424570 291218 424806 291454
rect 423930 290898 424166 291134
rect 424250 290898 424486 291134
rect 424570 290898 424806 291134
rect 443930 291218 444166 291454
rect 444250 291218 444486 291454
rect 444570 291218 444806 291454
rect 443930 290898 444166 291134
rect 444250 290898 444486 291134
rect 444570 290898 444806 291134
rect 463930 291218 464166 291454
rect 464250 291218 464486 291454
rect 464570 291218 464806 291454
rect 463930 290898 464166 291134
rect 464250 290898 464486 291134
rect 464570 290898 464806 291134
rect 483930 291218 484166 291454
rect 484250 291218 484486 291454
rect 484570 291218 484806 291454
rect 483930 290898 484166 291134
rect 484250 290898 484486 291134
rect 484570 290898 484806 291134
rect 503930 291218 504166 291454
rect 504250 291218 504486 291454
rect 504570 291218 504806 291454
rect 503930 290898 504166 291134
rect 504250 290898 504486 291134
rect 504570 290898 504806 291134
rect 523930 291218 524166 291454
rect 524250 291218 524486 291454
rect 524570 291218 524806 291454
rect 523930 290898 524166 291134
rect 524250 290898 524486 291134
rect 524570 290898 524806 291134
rect 543930 291218 544166 291454
rect 544250 291218 544486 291454
rect 544570 291218 544806 291454
rect 543930 290898 544166 291134
rect 544250 290898 544486 291134
rect 544570 290898 544806 291134
rect 563930 291218 564166 291454
rect 564250 291218 564486 291454
rect 564570 291218 564806 291454
rect 563930 290898 564166 291134
rect 564250 290898 564486 291134
rect 564570 290898 564806 291134
rect 313930 259718 314166 259954
rect 314250 259718 314486 259954
rect 314570 259718 314806 259954
rect 313930 259398 314166 259634
rect 314250 259398 314486 259634
rect 314570 259398 314806 259634
rect 333930 259718 334166 259954
rect 334250 259718 334486 259954
rect 334570 259718 334806 259954
rect 333930 259398 334166 259634
rect 334250 259398 334486 259634
rect 334570 259398 334806 259634
rect 353930 259718 354166 259954
rect 354250 259718 354486 259954
rect 354570 259718 354806 259954
rect 353930 259398 354166 259634
rect 354250 259398 354486 259634
rect 354570 259398 354806 259634
rect 373930 259718 374166 259954
rect 374250 259718 374486 259954
rect 374570 259718 374806 259954
rect 373930 259398 374166 259634
rect 374250 259398 374486 259634
rect 374570 259398 374806 259634
rect 393930 259718 394166 259954
rect 394250 259718 394486 259954
rect 394570 259718 394806 259954
rect 393930 259398 394166 259634
rect 394250 259398 394486 259634
rect 394570 259398 394806 259634
rect 413930 259718 414166 259954
rect 414250 259718 414486 259954
rect 414570 259718 414806 259954
rect 413930 259398 414166 259634
rect 414250 259398 414486 259634
rect 414570 259398 414806 259634
rect 433930 259718 434166 259954
rect 434250 259718 434486 259954
rect 434570 259718 434806 259954
rect 433930 259398 434166 259634
rect 434250 259398 434486 259634
rect 434570 259398 434806 259634
rect 453930 259718 454166 259954
rect 454250 259718 454486 259954
rect 454570 259718 454806 259954
rect 453930 259398 454166 259634
rect 454250 259398 454486 259634
rect 454570 259398 454806 259634
rect 473930 259718 474166 259954
rect 474250 259718 474486 259954
rect 474570 259718 474806 259954
rect 473930 259398 474166 259634
rect 474250 259398 474486 259634
rect 474570 259398 474806 259634
rect 493930 259718 494166 259954
rect 494250 259718 494486 259954
rect 494570 259718 494806 259954
rect 493930 259398 494166 259634
rect 494250 259398 494486 259634
rect 494570 259398 494806 259634
rect 513930 259718 514166 259954
rect 514250 259718 514486 259954
rect 514570 259718 514806 259954
rect 513930 259398 514166 259634
rect 514250 259398 514486 259634
rect 514570 259398 514806 259634
rect 533930 259718 534166 259954
rect 534250 259718 534486 259954
rect 534570 259718 534806 259954
rect 533930 259398 534166 259634
rect 534250 259398 534486 259634
rect 534570 259398 534806 259634
rect 553930 259718 554166 259954
rect 554250 259718 554486 259954
rect 554570 259718 554806 259954
rect 553930 259398 554166 259634
rect 554250 259398 554486 259634
rect 554570 259398 554806 259634
rect 303930 255218 304166 255454
rect 304250 255218 304486 255454
rect 304570 255218 304806 255454
rect 303930 254898 304166 255134
rect 304250 254898 304486 255134
rect 304570 254898 304806 255134
rect 323930 255218 324166 255454
rect 324250 255218 324486 255454
rect 324570 255218 324806 255454
rect 323930 254898 324166 255134
rect 324250 254898 324486 255134
rect 324570 254898 324806 255134
rect 343930 255218 344166 255454
rect 344250 255218 344486 255454
rect 344570 255218 344806 255454
rect 343930 254898 344166 255134
rect 344250 254898 344486 255134
rect 344570 254898 344806 255134
rect 363930 255218 364166 255454
rect 364250 255218 364486 255454
rect 364570 255218 364806 255454
rect 363930 254898 364166 255134
rect 364250 254898 364486 255134
rect 364570 254898 364806 255134
rect 383930 255218 384166 255454
rect 384250 255218 384486 255454
rect 384570 255218 384806 255454
rect 383930 254898 384166 255134
rect 384250 254898 384486 255134
rect 384570 254898 384806 255134
rect 403930 255218 404166 255454
rect 404250 255218 404486 255454
rect 404570 255218 404806 255454
rect 403930 254898 404166 255134
rect 404250 254898 404486 255134
rect 404570 254898 404806 255134
rect 423930 255218 424166 255454
rect 424250 255218 424486 255454
rect 424570 255218 424806 255454
rect 423930 254898 424166 255134
rect 424250 254898 424486 255134
rect 424570 254898 424806 255134
rect 443930 255218 444166 255454
rect 444250 255218 444486 255454
rect 444570 255218 444806 255454
rect 443930 254898 444166 255134
rect 444250 254898 444486 255134
rect 444570 254898 444806 255134
rect 463930 255218 464166 255454
rect 464250 255218 464486 255454
rect 464570 255218 464806 255454
rect 463930 254898 464166 255134
rect 464250 254898 464486 255134
rect 464570 254898 464806 255134
rect 483930 255218 484166 255454
rect 484250 255218 484486 255454
rect 484570 255218 484806 255454
rect 483930 254898 484166 255134
rect 484250 254898 484486 255134
rect 484570 254898 484806 255134
rect 503930 255218 504166 255454
rect 504250 255218 504486 255454
rect 504570 255218 504806 255454
rect 503930 254898 504166 255134
rect 504250 254898 504486 255134
rect 504570 254898 504806 255134
rect 523930 255218 524166 255454
rect 524250 255218 524486 255454
rect 524570 255218 524806 255454
rect 523930 254898 524166 255134
rect 524250 254898 524486 255134
rect 524570 254898 524806 255134
rect 543930 255218 544166 255454
rect 544250 255218 544486 255454
rect 544570 255218 544806 255454
rect 543930 254898 544166 255134
rect 544250 254898 544486 255134
rect 544570 254898 544806 255134
rect 563930 255218 564166 255454
rect 564250 255218 564486 255454
rect 564570 255218 564806 255454
rect 563930 254898 564166 255134
rect 564250 254898 564486 255134
rect 564570 254898 564806 255134
rect 313930 223718 314166 223954
rect 314250 223718 314486 223954
rect 314570 223718 314806 223954
rect 313930 223398 314166 223634
rect 314250 223398 314486 223634
rect 314570 223398 314806 223634
rect 333930 223718 334166 223954
rect 334250 223718 334486 223954
rect 334570 223718 334806 223954
rect 333930 223398 334166 223634
rect 334250 223398 334486 223634
rect 334570 223398 334806 223634
rect 353930 223718 354166 223954
rect 354250 223718 354486 223954
rect 354570 223718 354806 223954
rect 353930 223398 354166 223634
rect 354250 223398 354486 223634
rect 354570 223398 354806 223634
rect 373930 223718 374166 223954
rect 374250 223718 374486 223954
rect 374570 223718 374806 223954
rect 373930 223398 374166 223634
rect 374250 223398 374486 223634
rect 374570 223398 374806 223634
rect 393930 223718 394166 223954
rect 394250 223718 394486 223954
rect 394570 223718 394806 223954
rect 393930 223398 394166 223634
rect 394250 223398 394486 223634
rect 394570 223398 394806 223634
rect 413930 223718 414166 223954
rect 414250 223718 414486 223954
rect 414570 223718 414806 223954
rect 413930 223398 414166 223634
rect 414250 223398 414486 223634
rect 414570 223398 414806 223634
rect 433930 223718 434166 223954
rect 434250 223718 434486 223954
rect 434570 223718 434806 223954
rect 433930 223398 434166 223634
rect 434250 223398 434486 223634
rect 434570 223398 434806 223634
rect 453930 223718 454166 223954
rect 454250 223718 454486 223954
rect 454570 223718 454806 223954
rect 453930 223398 454166 223634
rect 454250 223398 454486 223634
rect 454570 223398 454806 223634
rect 473930 223718 474166 223954
rect 474250 223718 474486 223954
rect 474570 223718 474806 223954
rect 473930 223398 474166 223634
rect 474250 223398 474486 223634
rect 474570 223398 474806 223634
rect 493930 223718 494166 223954
rect 494250 223718 494486 223954
rect 494570 223718 494806 223954
rect 493930 223398 494166 223634
rect 494250 223398 494486 223634
rect 494570 223398 494806 223634
rect 513930 223718 514166 223954
rect 514250 223718 514486 223954
rect 514570 223718 514806 223954
rect 513930 223398 514166 223634
rect 514250 223398 514486 223634
rect 514570 223398 514806 223634
rect 533930 223718 534166 223954
rect 534250 223718 534486 223954
rect 534570 223718 534806 223954
rect 533930 223398 534166 223634
rect 534250 223398 534486 223634
rect 534570 223398 534806 223634
rect 553930 223718 554166 223954
rect 554250 223718 554486 223954
rect 554570 223718 554806 223954
rect 553930 223398 554166 223634
rect 554250 223398 554486 223634
rect 554570 223398 554806 223634
rect 303930 219218 304166 219454
rect 304250 219218 304486 219454
rect 304570 219218 304806 219454
rect 303930 218898 304166 219134
rect 304250 218898 304486 219134
rect 304570 218898 304806 219134
rect 323930 219218 324166 219454
rect 324250 219218 324486 219454
rect 324570 219218 324806 219454
rect 323930 218898 324166 219134
rect 324250 218898 324486 219134
rect 324570 218898 324806 219134
rect 343930 219218 344166 219454
rect 344250 219218 344486 219454
rect 344570 219218 344806 219454
rect 343930 218898 344166 219134
rect 344250 218898 344486 219134
rect 344570 218898 344806 219134
rect 363930 219218 364166 219454
rect 364250 219218 364486 219454
rect 364570 219218 364806 219454
rect 363930 218898 364166 219134
rect 364250 218898 364486 219134
rect 364570 218898 364806 219134
rect 383930 219218 384166 219454
rect 384250 219218 384486 219454
rect 384570 219218 384806 219454
rect 383930 218898 384166 219134
rect 384250 218898 384486 219134
rect 384570 218898 384806 219134
rect 403930 219218 404166 219454
rect 404250 219218 404486 219454
rect 404570 219218 404806 219454
rect 403930 218898 404166 219134
rect 404250 218898 404486 219134
rect 404570 218898 404806 219134
rect 423930 219218 424166 219454
rect 424250 219218 424486 219454
rect 424570 219218 424806 219454
rect 423930 218898 424166 219134
rect 424250 218898 424486 219134
rect 424570 218898 424806 219134
rect 443930 219218 444166 219454
rect 444250 219218 444486 219454
rect 444570 219218 444806 219454
rect 443930 218898 444166 219134
rect 444250 218898 444486 219134
rect 444570 218898 444806 219134
rect 463930 219218 464166 219454
rect 464250 219218 464486 219454
rect 464570 219218 464806 219454
rect 463930 218898 464166 219134
rect 464250 218898 464486 219134
rect 464570 218898 464806 219134
rect 483930 219218 484166 219454
rect 484250 219218 484486 219454
rect 484570 219218 484806 219454
rect 483930 218898 484166 219134
rect 484250 218898 484486 219134
rect 484570 218898 484806 219134
rect 503930 219218 504166 219454
rect 504250 219218 504486 219454
rect 504570 219218 504806 219454
rect 503930 218898 504166 219134
rect 504250 218898 504486 219134
rect 504570 218898 504806 219134
rect 523930 219218 524166 219454
rect 524250 219218 524486 219454
rect 524570 219218 524806 219454
rect 523930 218898 524166 219134
rect 524250 218898 524486 219134
rect 524570 218898 524806 219134
rect 543930 219218 544166 219454
rect 544250 219218 544486 219454
rect 544570 219218 544806 219454
rect 543930 218898 544166 219134
rect 544250 218898 544486 219134
rect 544570 218898 544806 219134
rect 563930 219218 564166 219454
rect 564250 219218 564486 219454
rect 564570 219218 564806 219454
rect 563930 218898 564166 219134
rect 564250 218898 564486 219134
rect 564570 218898 564806 219134
rect 303930 183218 304166 183454
rect 304250 183218 304486 183454
rect 304570 183218 304806 183454
rect 303930 182898 304166 183134
rect 304250 182898 304486 183134
rect 304570 182898 304806 183134
rect 323930 183218 324166 183454
rect 324250 183218 324486 183454
rect 324570 183218 324806 183454
rect 323930 182898 324166 183134
rect 324250 182898 324486 183134
rect 324570 182898 324806 183134
rect 343930 183218 344166 183454
rect 344250 183218 344486 183454
rect 344570 183218 344806 183454
rect 343930 182898 344166 183134
rect 344250 182898 344486 183134
rect 344570 182898 344806 183134
rect 363930 183218 364166 183454
rect 364250 183218 364486 183454
rect 364570 183218 364806 183454
rect 363930 182898 364166 183134
rect 364250 182898 364486 183134
rect 364570 182898 364806 183134
rect 383930 183218 384166 183454
rect 384250 183218 384486 183454
rect 384570 183218 384806 183454
rect 383930 182898 384166 183134
rect 384250 182898 384486 183134
rect 384570 182898 384806 183134
rect 403930 183218 404166 183454
rect 404250 183218 404486 183454
rect 404570 183218 404806 183454
rect 403930 182898 404166 183134
rect 404250 182898 404486 183134
rect 404570 182898 404806 183134
rect 423930 183218 424166 183454
rect 424250 183218 424486 183454
rect 424570 183218 424806 183454
rect 423930 182898 424166 183134
rect 424250 182898 424486 183134
rect 424570 182898 424806 183134
rect 443930 183218 444166 183454
rect 444250 183218 444486 183454
rect 444570 183218 444806 183454
rect 443930 182898 444166 183134
rect 444250 182898 444486 183134
rect 444570 182898 444806 183134
rect 463930 183218 464166 183454
rect 464250 183218 464486 183454
rect 464570 183218 464806 183454
rect 463930 182898 464166 183134
rect 464250 182898 464486 183134
rect 464570 182898 464806 183134
rect 483930 183218 484166 183454
rect 484250 183218 484486 183454
rect 484570 183218 484806 183454
rect 483930 182898 484166 183134
rect 484250 182898 484486 183134
rect 484570 182898 484806 183134
rect 503930 183218 504166 183454
rect 504250 183218 504486 183454
rect 504570 183218 504806 183454
rect 503930 182898 504166 183134
rect 504250 182898 504486 183134
rect 504570 182898 504806 183134
rect 523930 183218 524166 183454
rect 524250 183218 524486 183454
rect 524570 183218 524806 183454
rect 523930 182898 524166 183134
rect 524250 182898 524486 183134
rect 524570 182898 524806 183134
rect 543930 183218 544166 183454
rect 544250 183218 544486 183454
rect 544570 183218 544806 183454
rect 543930 182898 544166 183134
rect 544250 182898 544486 183134
rect 544570 182898 544806 183134
rect 563930 183218 564166 183454
rect 564250 183218 564486 183454
rect 564570 183218 564806 183454
rect 563930 182898 564166 183134
rect 564250 182898 564486 183134
rect 564570 182898 564806 183134
rect 313930 151718 314166 151954
rect 314250 151718 314486 151954
rect 314570 151718 314806 151954
rect 313930 151398 314166 151634
rect 314250 151398 314486 151634
rect 314570 151398 314806 151634
rect 333930 151718 334166 151954
rect 334250 151718 334486 151954
rect 334570 151718 334806 151954
rect 333930 151398 334166 151634
rect 334250 151398 334486 151634
rect 334570 151398 334806 151634
rect 353930 151718 354166 151954
rect 354250 151718 354486 151954
rect 354570 151718 354806 151954
rect 353930 151398 354166 151634
rect 354250 151398 354486 151634
rect 354570 151398 354806 151634
rect 373930 151718 374166 151954
rect 374250 151718 374486 151954
rect 374570 151718 374806 151954
rect 373930 151398 374166 151634
rect 374250 151398 374486 151634
rect 374570 151398 374806 151634
rect 393930 151718 394166 151954
rect 394250 151718 394486 151954
rect 394570 151718 394806 151954
rect 393930 151398 394166 151634
rect 394250 151398 394486 151634
rect 394570 151398 394806 151634
rect 413930 151718 414166 151954
rect 414250 151718 414486 151954
rect 414570 151718 414806 151954
rect 413930 151398 414166 151634
rect 414250 151398 414486 151634
rect 414570 151398 414806 151634
rect 433930 151718 434166 151954
rect 434250 151718 434486 151954
rect 434570 151718 434806 151954
rect 433930 151398 434166 151634
rect 434250 151398 434486 151634
rect 434570 151398 434806 151634
rect 453930 151718 454166 151954
rect 454250 151718 454486 151954
rect 454570 151718 454806 151954
rect 453930 151398 454166 151634
rect 454250 151398 454486 151634
rect 454570 151398 454806 151634
rect 473930 151718 474166 151954
rect 474250 151718 474486 151954
rect 474570 151718 474806 151954
rect 473930 151398 474166 151634
rect 474250 151398 474486 151634
rect 474570 151398 474806 151634
rect 493930 151718 494166 151954
rect 494250 151718 494486 151954
rect 494570 151718 494806 151954
rect 493930 151398 494166 151634
rect 494250 151398 494486 151634
rect 494570 151398 494806 151634
rect 513930 151718 514166 151954
rect 514250 151718 514486 151954
rect 514570 151718 514806 151954
rect 513930 151398 514166 151634
rect 514250 151398 514486 151634
rect 514570 151398 514806 151634
rect 533930 151718 534166 151954
rect 534250 151718 534486 151954
rect 534570 151718 534806 151954
rect 533930 151398 534166 151634
rect 534250 151398 534486 151634
rect 534570 151398 534806 151634
rect 553930 151718 554166 151954
rect 554250 151718 554486 151954
rect 554570 151718 554806 151954
rect 553930 151398 554166 151634
rect 554250 151398 554486 151634
rect 554570 151398 554806 151634
rect 303930 147218 304166 147454
rect 304250 147218 304486 147454
rect 304570 147218 304806 147454
rect 303930 146898 304166 147134
rect 304250 146898 304486 147134
rect 304570 146898 304806 147134
rect 323930 147218 324166 147454
rect 324250 147218 324486 147454
rect 324570 147218 324806 147454
rect 323930 146898 324166 147134
rect 324250 146898 324486 147134
rect 324570 146898 324806 147134
rect 343930 147218 344166 147454
rect 344250 147218 344486 147454
rect 344570 147218 344806 147454
rect 343930 146898 344166 147134
rect 344250 146898 344486 147134
rect 344570 146898 344806 147134
rect 363930 147218 364166 147454
rect 364250 147218 364486 147454
rect 364570 147218 364806 147454
rect 363930 146898 364166 147134
rect 364250 146898 364486 147134
rect 364570 146898 364806 147134
rect 383930 147218 384166 147454
rect 384250 147218 384486 147454
rect 384570 147218 384806 147454
rect 383930 146898 384166 147134
rect 384250 146898 384486 147134
rect 384570 146898 384806 147134
rect 403930 147218 404166 147454
rect 404250 147218 404486 147454
rect 404570 147218 404806 147454
rect 403930 146898 404166 147134
rect 404250 146898 404486 147134
rect 404570 146898 404806 147134
rect 423930 147218 424166 147454
rect 424250 147218 424486 147454
rect 424570 147218 424806 147454
rect 423930 146898 424166 147134
rect 424250 146898 424486 147134
rect 424570 146898 424806 147134
rect 443930 147218 444166 147454
rect 444250 147218 444486 147454
rect 444570 147218 444806 147454
rect 443930 146898 444166 147134
rect 444250 146898 444486 147134
rect 444570 146898 444806 147134
rect 463930 147218 464166 147454
rect 464250 147218 464486 147454
rect 464570 147218 464806 147454
rect 463930 146898 464166 147134
rect 464250 146898 464486 147134
rect 464570 146898 464806 147134
rect 483930 147218 484166 147454
rect 484250 147218 484486 147454
rect 484570 147218 484806 147454
rect 483930 146898 484166 147134
rect 484250 146898 484486 147134
rect 484570 146898 484806 147134
rect 503930 147218 504166 147454
rect 504250 147218 504486 147454
rect 504570 147218 504806 147454
rect 503930 146898 504166 147134
rect 504250 146898 504486 147134
rect 504570 146898 504806 147134
rect 523930 147218 524166 147454
rect 524250 147218 524486 147454
rect 524570 147218 524806 147454
rect 523930 146898 524166 147134
rect 524250 146898 524486 147134
rect 524570 146898 524806 147134
rect 543930 147218 544166 147454
rect 544250 147218 544486 147454
rect 544570 147218 544806 147454
rect 543930 146898 544166 147134
rect 544250 146898 544486 147134
rect 544570 146898 544806 147134
rect 563930 147218 564166 147454
rect 564250 147218 564486 147454
rect 564570 147218 564806 147454
rect 563930 146898 564166 147134
rect 564250 146898 564486 147134
rect 564570 146898 564806 147134
rect 313930 115718 314166 115954
rect 314250 115718 314486 115954
rect 314570 115718 314806 115954
rect 313930 115398 314166 115634
rect 314250 115398 314486 115634
rect 314570 115398 314806 115634
rect 333930 115718 334166 115954
rect 334250 115718 334486 115954
rect 334570 115718 334806 115954
rect 333930 115398 334166 115634
rect 334250 115398 334486 115634
rect 334570 115398 334806 115634
rect 353930 115718 354166 115954
rect 354250 115718 354486 115954
rect 354570 115718 354806 115954
rect 353930 115398 354166 115634
rect 354250 115398 354486 115634
rect 354570 115398 354806 115634
rect 373930 115718 374166 115954
rect 374250 115718 374486 115954
rect 374570 115718 374806 115954
rect 373930 115398 374166 115634
rect 374250 115398 374486 115634
rect 374570 115398 374806 115634
rect 393930 115718 394166 115954
rect 394250 115718 394486 115954
rect 394570 115718 394806 115954
rect 393930 115398 394166 115634
rect 394250 115398 394486 115634
rect 394570 115398 394806 115634
rect 413930 115718 414166 115954
rect 414250 115718 414486 115954
rect 414570 115718 414806 115954
rect 413930 115398 414166 115634
rect 414250 115398 414486 115634
rect 414570 115398 414806 115634
rect 433930 115718 434166 115954
rect 434250 115718 434486 115954
rect 434570 115718 434806 115954
rect 433930 115398 434166 115634
rect 434250 115398 434486 115634
rect 434570 115398 434806 115634
rect 453930 115718 454166 115954
rect 454250 115718 454486 115954
rect 454570 115718 454806 115954
rect 453930 115398 454166 115634
rect 454250 115398 454486 115634
rect 454570 115398 454806 115634
rect 473930 115718 474166 115954
rect 474250 115718 474486 115954
rect 474570 115718 474806 115954
rect 473930 115398 474166 115634
rect 474250 115398 474486 115634
rect 474570 115398 474806 115634
rect 493930 115718 494166 115954
rect 494250 115718 494486 115954
rect 494570 115718 494806 115954
rect 493930 115398 494166 115634
rect 494250 115398 494486 115634
rect 494570 115398 494806 115634
rect 513930 115718 514166 115954
rect 514250 115718 514486 115954
rect 514570 115718 514806 115954
rect 513930 115398 514166 115634
rect 514250 115398 514486 115634
rect 514570 115398 514806 115634
rect 533930 115718 534166 115954
rect 534250 115718 534486 115954
rect 534570 115718 534806 115954
rect 533930 115398 534166 115634
rect 534250 115398 534486 115634
rect 534570 115398 534806 115634
rect 553930 115718 554166 115954
rect 554250 115718 554486 115954
rect 554570 115718 554806 115954
rect 553930 115398 554166 115634
rect 554250 115398 554486 115634
rect 554570 115398 554806 115634
rect 303930 111218 304166 111454
rect 304250 111218 304486 111454
rect 304570 111218 304806 111454
rect 303930 110898 304166 111134
rect 304250 110898 304486 111134
rect 304570 110898 304806 111134
rect 323930 111218 324166 111454
rect 324250 111218 324486 111454
rect 324570 111218 324806 111454
rect 323930 110898 324166 111134
rect 324250 110898 324486 111134
rect 324570 110898 324806 111134
rect 343930 111218 344166 111454
rect 344250 111218 344486 111454
rect 344570 111218 344806 111454
rect 343930 110898 344166 111134
rect 344250 110898 344486 111134
rect 344570 110898 344806 111134
rect 363930 111218 364166 111454
rect 364250 111218 364486 111454
rect 364570 111218 364806 111454
rect 363930 110898 364166 111134
rect 364250 110898 364486 111134
rect 364570 110898 364806 111134
rect 383930 111218 384166 111454
rect 384250 111218 384486 111454
rect 384570 111218 384806 111454
rect 383930 110898 384166 111134
rect 384250 110898 384486 111134
rect 384570 110898 384806 111134
rect 403930 111218 404166 111454
rect 404250 111218 404486 111454
rect 404570 111218 404806 111454
rect 403930 110898 404166 111134
rect 404250 110898 404486 111134
rect 404570 110898 404806 111134
rect 423930 111218 424166 111454
rect 424250 111218 424486 111454
rect 424570 111218 424806 111454
rect 423930 110898 424166 111134
rect 424250 110898 424486 111134
rect 424570 110898 424806 111134
rect 443930 111218 444166 111454
rect 444250 111218 444486 111454
rect 444570 111218 444806 111454
rect 443930 110898 444166 111134
rect 444250 110898 444486 111134
rect 444570 110898 444806 111134
rect 463930 111218 464166 111454
rect 464250 111218 464486 111454
rect 464570 111218 464806 111454
rect 463930 110898 464166 111134
rect 464250 110898 464486 111134
rect 464570 110898 464806 111134
rect 483930 111218 484166 111454
rect 484250 111218 484486 111454
rect 484570 111218 484806 111454
rect 483930 110898 484166 111134
rect 484250 110898 484486 111134
rect 484570 110898 484806 111134
rect 503930 111218 504166 111454
rect 504250 111218 504486 111454
rect 504570 111218 504806 111454
rect 503930 110898 504166 111134
rect 504250 110898 504486 111134
rect 504570 110898 504806 111134
rect 523930 111218 524166 111454
rect 524250 111218 524486 111454
rect 524570 111218 524806 111454
rect 523930 110898 524166 111134
rect 524250 110898 524486 111134
rect 524570 110898 524806 111134
rect 543930 111218 544166 111454
rect 544250 111218 544486 111454
rect 544570 111218 544806 111454
rect 543930 110898 544166 111134
rect 544250 110898 544486 111134
rect 544570 110898 544806 111134
rect 563930 111218 564166 111454
rect 564250 111218 564486 111454
rect 564570 111218 564806 111454
rect 563930 110898 564166 111134
rect 564250 110898 564486 111134
rect 564570 110898 564806 111134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 167930 43718 168166 43954
rect 168250 43718 168486 43954
rect 168570 43718 168806 43954
rect 167930 43398 168166 43634
rect 168250 43398 168486 43634
rect 168570 43398 168806 43634
rect 187930 43718 188166 43954
rect 188250 43718 188486 43954
rect 188570 43718 188806 43954
rect 187930 43398 188166 43634
rect 188250 43398 188486 43634
rect 188570 43398 188806 43634
rect 207930 43718 208166 43954
rect 208250 43718 208486 43954
rect 208570 43718 208806 43954
rect 207930 43398 208166 43634
rect 208250 43398 208486 43634
rect 208570 43398 208806 43634
rect 227930 43718 228166 43954
rect 228250 43718 228486 43954
rect 228570 43718 228806 43954
rect 227930 43398 228166 43634
rect 228250 43398 228486 43634
rect 228570 43398 228806 43634
rect 247930 43718 248166 43954
rect 248250 43718 248486 43954
rect 248570 43718 248806 43954
rect 247930 43398 248166 43634
rect 248250 43398 248486 43634
rect 248570 43398 248806 43634
rect 267930 43718 268166 43954
rect 268250 43718 268486 43954
rect 268570 43718 268806 43954
rect 267930 43398 268166 43634
rect 268250 43398 268486 43634
rect 268570 43398 268806 43634
rect 287930 43718 288166 43954
rect 288250 43718 288486 43954
rect 288570 43718 288806 43954
rect 287930 43398 288166 43634
rect 288250 43398 288486 43634
rect 288570 43398 288806 43634
rect 307930 43718 308166 43954
rect 308250 43718 308486 43954
rect 308570 43718 308806 43954
rect 307930 43398 308166 43634
rect 308250 43398 308486 43634
rect 308570 43398 308806 43634
rect 327930 43718 328166 43954
rect 328250 43718 328486 43954
rect 328570 43718 328806 43954
rect 327930 43398 328166 43634
rect 328250 43398 328486 43634
rect 328570 43398 328806 43634
rect 347930 43718 348166 43954
rect 348250 43718 348486 43954
rect 348570 43718 348806 43954
rect 347930 43398 348166 43634
rect 348250 43398 348486 43634
rect 348570 43398 348806 43634
rect 367930 43718 368166 43954
rect 368250 43718 368486 43954
rect 368570 43718 368806 43954
rect 367930 43398 368166 43634
rect 368250 43398 368486 43634
rect 368570 43398 368806 43634
rect 387930 43718 388166 43954
rect 388250 43718 388486 43954
rect 388570 43718 388806 43954
rect 387930 43398 388166 43634
rect 388250 43398 388486 43634
rect 388570 43398 388806 43634
rect 407930 43718 408166 43954
rect 408250 43718 408486 43954
rect 408570 43718 408806 43954
rect 407930 43398 408166 43634
rect 408250 43398 408486 43634
rect 408570 43398 408806 43634
rect 427930 43718 428166 43954
rect 428250 43718 428486 43954
rect 428570 43718 428806 43954
rect 427930 43398 428166 43634
rect 428250 43398 428486 43634
rect 428570 43398 428806 43634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 157930 39218 158166 39454
rect 158250 39218 158486 39454
rect 158570 39218 158806 39454
rect 157930 38898 158166 39134
rect 158250 38898 158486 39134
rect 158570 38898 158806 39134
rect 177930 39218 178166 39454
rect 178250 39218 178486 39454
rect 178570 39218 178806 39454
rect 177930 38898 178166 39134
rect 178250 38898 178486 39134
rect 178570 38898 178806 39134
rect 197930 39218 198166 39454
rect 198250 39218 198486 39454
rect 198570 39218 198806 39454
rect 197930 38898 198166 39134
rect 198250 38898 198486 39134
rect 198570 38898 198806 39134
rect 217930 39218 218166 39454
rect 218250 39218 218486 39454
rect 218570 39218 218806 39454
rect 217930 38898 218166 39134
rect 218250 38898 218486 39134
rect 218570 38898 218806 39134
rect 237930 39218 238166 39454
rect 238250 39218 238486 39454
rect 238570 39218 238806 39454
rect 237930 38898 238166 39134
rect 238250 38898 238486 39134
rect 238570 38898 238806 39134
rect 257930 39218 258166 39454
rect 258250 39218 258486 39454
rect 258570 39218 258806 39454
rect 257930 38898 258166 39134
rect 258250 38898 258486 39134
rect 258570 38898 258806 39134
rect 277930 39218 278166 39454
rect 278250 39218 278486 39454
rect 278570 39218 278806 39454
rect 277930 38898 278166 39134
rect 278250 38898 278486 39134
rect 278570 38898 278806 39134
rect 297930 39218 298166 39454
rect 298250 39218 298486 39454
rect 298570 39218 298806 39454
rect 297930 38898 298166 39134
rect 298250 38898 298486 39134
rect 298570 38898 298806 39134
rect 317930 39218 318166 39454
rect 318250 39218 318486 39454
rect 318570 39218 318806 39454
rect 317930 38898 318166 39134
rect 318250 38898 318486 39134
rect 318570 38898 318806 39134
rect 337930 39218 338166 39454
rect 338250 39218 338486 39454
rect 338570 39218 338806 39454
rect 337930 38898 338166 39134
rect 338250 38898 338486 39134
rect 338570 38898 338806 39134
rect 357930 39218 358166 39454
rect 358250 39218 358486 39454
rect 358570 39218 358806 39454
rect 357930 38898 358166 39134
rect 358250 38898 358486 39134
rect 358570 38898 358806 39134
rect 377930 39218 378166 39454
rect 378250 39218 378486 39454
rect 378570 39218 378806 39454
rect 377930 38898 378166 39134
rect 378250 38898 378486 39134
rect 378570 38898 378806 39134
rect 397930 39218 398166 39454
rect 398250 39218 398486 39454
rect 398570 39218 398806 39454
rect 397930 38898 398166 39134
rect 398250 38898 398486 39134
rect 398570 38898 398806 39134
rect 417930 39218 418166 39454
rect 418250 39218 418486 39454
rect 418570 39218 418806 39454
rect 417930 38898 418166 39134
rect 418250 38898 418486 39134
rect 418570 38898 418806 39134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 213930 691954
rect 214166 691718 214250 691954
rect 214486 691718 214570 691954
rect 214806 691718 233930 691954
rect 234166 691718 234250 691954
rect 234486 691718 234570 691954
rect 234806 691718 253930 691954
rect 254166 691718 254250 691954
rect 254486 691718 254570 691954
rect 254806 691718 273930 691954
rect 274166 691718 274250 691954
rect 274486 691718 274570 691954
rect 274806 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 493930 691954
rect 494166 691718 494250 691954
rect 494486 691718 494570 691954
rect 494806 691718 513930 691954
rect 514166 691718 514250 691954
rect 514486 691718 514570 691954
rect 514806 691718 533930 691954
rect 534166 691718 534250 691954
rect 534486 691718 534570 691954
rect 534806 691718 553930 691954
rect 554166 691718 554250 691954
rect 554486 691718 554570 691954
rect 554806 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 213930 691634
rect 214166 691398 214250 691634
rect 214486 691398 214570 691634
rect 214806 691398 233930 691634
rect 234166 691398 234250 691634
rect 234486 691398 234570 691634
rect 234806 691398 253930 691634
rect 254166 691398 254250 691634
rect 254486 691398 254570 691634
rect 254806 691398 273930 691634
rect 274166 691398 274250 691634
rect 274486 691398 274570 691634
rect 274806 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 493930 691634
rect 494166 691398 494250 691634
rect 494486 691398 494570 691634
rect 494806 691398 513930 691634
rect 514166 691398 514250 691634
rect 514486 691398 514570 691634
rect 514806 691398 533930 691634
rect 534166 691398 534250 691634
rect 534486 691398 534570 691634
rect 534806 691398 553930 691634
rect 554166 691398 554250 691634
rect 554486 691398 554570 691634
rect 554806 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 203930 687454
rect 204166 687218 204250 687454
rect 204486 687218 204570 687454
rect 204806 687218 223930 687454
rect 224166 687218 224250 687454
rect 224486 687218 224570 687454
rect 224806 687218 243930 687454
rect 244166 687218 244250 687454
rect 244486 687218 244570 687454
rect 244806 687218 263930 687454
rect 264166 687218 264250 687454
rect 264486 687218 264570 687454
rect 264806 687218 283930 687454
rect 284166 687218 284250 687454
rect 284486 687218 284570 687454
rect 284806 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 483930 687454
rect 484166 687218 484250 687454
rect 484486 687218 484570 687454
rect 484806 687218 503930 687454
rect 504166 687218 504250 687454
rect 504486 687218 504570 687454
rect 504806 687218 523930 687454
rect 524166 687218 524250 687454
rect 524486 687218 524570 687454
rect 524806 687218 543930 687454
rect 544166 687218 544250 687454
rect 544486 687218 544570 687454
rect 544806 687218 563930 687454
rect 564166 687218 564250 687454
rect 564486 687218 564570 687454
rect 564806 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 203930 687134
rect 204166 686898 204250 687134
rect 204486 686898 204570 687134
rect 204806 686898 223930 687134
rect 224166 686898 224250 687134
rect 224486 686898 224570 687134
rect 224806 686898 243930 687134
rect 244166 686898 244250 687134
rect 244486 686898 244570 687134
rect 244806 686898 263930 687134
rect 264166 686898 264250 687134
rect 264486 686898 264570 687134
rect 264806 686898 283930 687134
rect 284166 686898 284250 687134
rect 284486 686898 284570 687134
rect 284806 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 483930 687134
rect 484166 686898 484250 687134
rect 484486 686898 484570 687134
rect 484806 686898 503930 687134
rect 504166 686898 504250 687134
rect 504486 686898 504570 687134
rect 504806 686898 523930 687134
rect 524166 686898 524250 687134
rect 524486 686898 524570 687134
rect 524806 686898 543930 687134
rect 544166 686898 544250 687134
rect 544486 686898 544570 687134
rect 544806 686898 563930 687134
rect 564166 686898 564250 687134
rect 564486 686898 564570 687134
rect 564806 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 213930 655954
rect 214166 655718 214250 655954
rect 214486 655718 214570 655954
rect 214806 655718 233930 655954
rect 234166 655718 234250 655954
rect 234486 655718 234570 655954
rect 234806 655718 253930 655954
rect 254166 655718 254250 655954
rect 254486 655718 254570 655954
rect 254806 655718 273930 655954
rect 274166 655718 274250 655954
rect 274486 655718 274570 655954
rect 274806 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 493930 655954
rect 494166 655718 494250 655954
rect 494486 655718 494570 655954
rect 494806 655718 513930 655954
rect 514166 655718 514250 655954
rect 514486 655718 514570 655954
rect 514806 655718 533930 655954
rect 534166 655718 534250 655954
rect 534486 655718 534570 655954
rect 534806 655718 553930 655954
rect 554166 655718 554250 655954
rect 554486 655718 554570 655954
rect 554806 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 213930 655634
rect 214166 655398 214250 655634
rect 214486 655398 214570 655634
rect 214806 655398 233930 655634
rect 234166 655398 234250 655634
rect 234486 655398 234570 655634
rect 234806 655398 253930 655634
rect 254166 655398 254250 655634
rect 254486 655398 254570 655634
rect 254806 655398 273930 655634
rect 274166 655398 274250 655634
rect 274486 655398 274570 655634
rect 274806 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 493930 655634
rect 494166 655398 494250 655634
rect 494486 655398 494570 655634
rect 494806 655398 513930 655634
rect 514166 655398 514250 655634
rect 514486 655398 514570 655634
rect 514806 655398 533930 655634
rect 534166 655398 534250 655634
rect 534486 655398 534570 655634
rect 534806 655398 553930 655634
rect 554166 655398 554250 655634
rect 554486 655398 554570 655634
rect 554806 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 203930 651454
rect 204166 651218 204250 651454
rect 204486 651218 204570 651454
rect 204806 651218 223930 651454
rect 224166 651218 224250 651454
rect 224486 651218 224570 651454
rect 224806 651218 243930 651454
rect 244166 651218 244250 651454
rect 244486 651218 244570 651454
rect 244806 651218 263930 651454
rect 264166 651218 264250 651454
rect 264486 651218 264570 651454
rect 264806 651218 283930 651454
rect 284166 651218 284250 651454
rect 284486 651218 284570 651454
rect 284806 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 483930 651454
rect 484166 651218 484250 651454
rect 484486 651218 484570 651454
rect 484806 651218 503930 651454
rect 504166 651218 504250 651454
rect 504486 651218 504570 651454
rect 504806 651218 523930 651454
rect 524166 651218 524250 651454
rect 524486 651218 524570 651454
rect 524806 651218 543930 651454
rect 544166 651218 544250 651454
rect 544486 651218 544570 651454
rect 544806 651218 563930 651454
rect 564166 651218 564250 651454
rect 564486 651218 564570 651454
rect 564806 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 203930 651134
rect 204166 650898 204250 651134
rect 204486 650898 204570 651134
rect 204806 650898 223930 651134
rect 224166 650898 224250 651134
rect 224486 650898 224570 651134
rect 224806 650898 243930 651134
rect 244166 650898 244250 651134
rect 244486 650898 244570 651134
rect 244806 650898 263930 651134
rect 264166 650898 264250 651134
rect 264486 650898 264570 651134
rect 264806 650898 283930 651134
rect 284166 650898 284250 651134
rect 284486 650898 284570 651134
rect 284806 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 483930 651134
rect 484166 650898 484250 651134
rect 484486 650898 484570 651134
rect 484806 650898 503930 651134
rect 504166 650898 504250 651134
rect 504486 650898 504570 651134
rect 504806 650898 523930 651134
rect 524166 650898 524250 651134
rect 524486 650898 524570 651134
rect 524806 650898 543930 651134
rect 544166 650898 544250 651134
rect 544486 650898 544570 651134
rect 544806 650898 563930 651134
rect 564166 650898 564250 651134
rect 564486 650898 564570 651134
rect 564806 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 213930 619954
rect 214166 619718 214250 619954
rect 214486 619718 214570 619954
rect 214806 619718 233930 619954
rect 234166 619718 234250 619954
rect 234486 619718 234570 619954
rect 234806 619718 253930 619954
rect 254166 619718 254250 619954
rect 254486 619718 254570 619954
rect 254806 619718 273930 619954
rect 274166 619718 274250 619954
rect 274486 619718 274570 619954
rect 274806 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 493930 619954
rect 494166 619718 494250 619954
rect 494486 619718 494570 619954
rect 494806 619718 513930 619954
rect 514166 619718 514250 619954
rect 514486 619718 514570 619954
rect 514806 619718 533930 619954
rect 534166 619718 534250 619954
rect 534486 619718 534570 619954
rect 534806 619718 553930 619954
rect 554166 619718 554250 619954
rect 554486 619718 554570 619954
rect 554806 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 213930 619634
rect 214166 619398 214250 619634
rect 214486 619398 214570 619634
rect 214806 619398 233930 619634
rect 234166 619398 234250 619634
rect 234486 619398 234570 619634
rect 234806 619398 253930 619634
rect 254166 619398 254250 619634
rect 254486 619398 254570 619634
rect 254806 619398 273930 619634
rect 274166 619398 274250 619634
rect 274486 619398 274570 619634
rect 274806 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 493930 619634
rect 494166 619398 494250 619634
rect 494486 619398 494570 619634
rect 494806 619398 513930 619634
rect 514166 619398 514250 619634
rect 514486 619398 514570 619634
rect 514806 619398 533930 619634
rect 534166 619398 534250 619634
rect 534486 619398 534570 619634
rect 534806 619398 553930 619634
rect 554166 619398 554250 619634
rect 554486 619398 554570 619634
rect 554806 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 203930 615454
rect 204166 615218 204250 615454
rect 204486 615218 204570 615454
rect 204806 615218 223930 615454
rect 224166 615218 224250 615454
rect 224486 615218 224570 615454
rect 224806 615218 243930 615454
rect 244166 615218 244250 615454
rect 244486 615218 244570 615454
rect 244806 615218 263930 615454
rect 264166 615218 264250 615454
rect 264486 615218 264570 615454
rect 264806 615218 283930 615454
rect 284166 615218 284250 615454
rect 284486 615218 284570 615454
rect 284806 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 483930 615454
rect 484166 615218 484250 615454
rect 484486 615218 484570 615454
rect 484806 615218 503930 615454
rect 504166 615218 504250 615454
rect 504486 615218 504570 615454
rect 504806 615218 523930 615454
rect 524166 615218 524250 615454
rect 524486 615218 524570 615454
rect 524806 615218 543930 615454
rect 544166 615218 544250 615454
rect 544486 615218 544570 615454
rect 544806 615218 563930 615454
rect 564166 615218 564250 615454
rect 564486 615218 564570 615454
rect 564806 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 203930 615134
rect 204166 614898 204250 615134
rect 204486 614898 204570 615134
rect 204806 614898 223930 615134
rect 224166 614898 224250 615134
rect 224486 614898 224570 615134
rect 224806 614898 243930 615134
rect 244166 614898 244250 615134
rect 244486 614898 244570 615134
rect 244806 614898 263930 615134
rect 264166 614898 264250 615134
rect 264486 614898 264570 615134
rect 264806 614898 283930 615134
rect 284166 614898 284250 615134
rect 284486 614898 284570 615134
rect 284806 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 483930 615134
rect 484166 614898 484250 615134
rect 484486 614898 484570 615134
rect 484806 614898 503930 615134
rect 504166 614898 504250 615134
rect 504486 614898 504570 615134
rect 504806 614898 523930 615134
rect 524166 614898 524250 615134
rect 524486 614898 524570 615134
rect 524806 614898 543930 615134
rect 544166 614898 544250 615134
rect 544486 614898 544570 615134
rect 544806 614898 563930 615134
rect 564166 614898 564250 615134
rect 564486 614898 564570 615134
rect 564806 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 213930 547954
rect 214166 547718 214250 547954
rect 214486 547718 214570 547954
rect 214806 547718 233930 547954
rect 234166 547718 234250 547954
rect 234486 547718 234570 547954
rect 234806 547718 253930 547954
rect 254166 547718 254250 547954
rect 254486 547718 254570 547954
rect 254806 547718 273930 547954
rect 274166 547718 274250 547954
rect 274486 547718 274570 547954
rect 274806 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 493930 547954
rect 494166 547718 494250 547954
rect 494486 547718 494570 547954
rect 494806 547718 513930 547954
rect 514166 547718 514250 547954
rect 514486 547718 514570 547954
rect 514806 547718 533930 547954
rect 534166 547718 534250 547954
rect 534486 547718 534570 547954
rect 534806 547718 553930 547954
rect 554166 547718 554250 547954
rect 554486 547718 554570 547954
rect 554806 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 213930 547634
rect 214166 547398 214250 547634
rect 214486 547398 214570 547634
rect 214806 547398 233930 547634
rect 234166 547398 234250 547634
rect 234486 547398 234570 547634
rect 234806 547398 253930 547634
rect 254166 547398 254250 547634
rect 254486 547398 254570 547634
rect 254806 547398 273930 547634
rect 274166 547398 274250 547634
rect 274486 547398 274570 547634
rect 274806 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 493930 547634
rect 494166 547398 494250 547634
rect 494486 547398 494570 547634
rect 494806 547398 513930 547634
rect 514166 547398 514250 547634
rect 514486 547398 514570 547634
rect 514806 547398 533930 547634
rect 534166 547398 534250 547634
rect 534486 547398 534570 547634
rect 534806 547398 553930 547634
rect 554166 547398 554250 547634
rect 554486 547398 554570 547634
rect 554806 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 203930 543454
rect 204166 543218 204250 543454
rect 204486 543218 204570 543454
rect 204806 543218 223930 543454
rect 224166 543218 224250 543454
rect 224486 543218 224570 543454
rect 224806 543218 243930 543454
rect 244166 543218 244250 543454
rect 244486 543218 244570 543454
rect 244806 543218 263930 543454
rect 264166 543218 264250 543454
rect 264486 543218 264570 543454
rect 264806 543218 283930 543454
rect 284166 543218 284250 543454
rect 284486 543218 284570 543454
rect 284806 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 483930 543454
rect 484166 543218 484250 543454
rect 484486 543218 484570 543454
rect 484806 543218 503930 543454
rect 504166 543218 504250 543454
rect 504486 543218 504570 543454
rect 504806 543218 523930 543454
rect 524166 543218 524250 543454
rect 524486 543218 524570 543454
rect 524806 543218 543930 543454
rect 544166 543218 544250 543454
rect 544486 543218 544570 543454
rect 544806 543218 563930 543454
rect 564166 543218 564250 543454
rect 564486 543218 564570 543454
rect 564806 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 203930 543134
rect 204166 542898 204250 543134
rect 204486 542898 204570 543134
rect 204806 542898 223930 543134
rect 224166 542898 224250 543134
rect 224486 542898 224570 543134
rect 224806 542898 243930 543134
rect 244166 542898 244250 543134
rect 244486 542898 244570 543134
rect 244806 542898 263930 543134
rect 264166 542898 264250 543134
rect 264486 542898 264570 543134
rect 264806 542898 283930 543134
rect 284166 542898 284250 543134
rect 284486 542898 284570 543134
rect 284806 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 483930 543134
rect 484166 542898 484250 543134
rect 484486 542898 484570 543134
rect 484806 542898 503930 543134
rect 504166 542898 504250 543134
rect 504486 542898 504570 543134
rect 504806 542898 523930 543134
rect 524166 542898 524250 543134
rect 524486 542898 524570 543134
rect 524806 542898 543930 543134
rect 544166 542898 544250 543134
rect 544486 542898 544570 543134
rect 544806 542898 563930 543134
rect 564166 542898 564250 543134
rect 564486 542898 564570 543134
rect 564806 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 213930 511954
rect 214166 511718 214250 511954
rect 214486 511718 214570 511954
rect 214806 511718 233930 511954
rect 234166 511718 234250 511954
rect 234486 511718 234570 511954
rect 234806 511718 253930 511954
rect 254166 511718 254250 511954
rect 254486 511718 254570 511954
rect 254806 511718 273930 511954
rect 274166 511718 274250 511954
rect 274486 511718 274570 511954
rect 274806 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 493930 511954
rect 494166 511718 494250 511954
rect 494486 511718 494570 511954
rect 494806 511718 513930 511954
rect 514166 511718 514250 511954
rect 514486 511718 514570 511954
rect 514806 511718 533930 511954
rect 534166 511718 534250 511954
rect 534486 511718 534570 511954
rect 534806 511718 553930 511954
rect 554166 511718 554250 511954
rect 554486 511718 554570 511954
rect 554806 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 213930 511634
rect 214166 511398 214250 511634
rect 214486 511398 214570 511634
rect 214806 511398 233930 511634
rect 234166 511398 234250 511634
rect 234486 511398 234570 511634
rect 234806 511398 253930 511634
rect 254166 511398 254250 511634
rect 254486 511398 254570 511634
rect 254806 511398 273930 511634
rect 274166 511398 274250 511634
rect 274486 511398 274570 511634
rect 274806 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 493930 511634
rect 494166 511398 494250 511634
rect 494486 511398 494570 511634
rect 494806 511398 513930 511634
rect 514166 511398 514250 511634
rect 514486 511398 514570 511634
rect 514806 511398 533930 511634
rect 534166 511398 534250 511634
rect 534486 511398 534570 511634
rect 534806 511398 553930 511634
rect 554166 511398 554250 511634
rect 554486 511398 554570 511634
rect 554806 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 203930 507454
rect 204166 507218 204250 507454
rect 204486 507218 204570 507454
rect 204806 507218 223930 507454
rect 224166 507218 224250 507454
rect 224486 507218 224570 507454
rect 224806 507218 243930 507454
rect 244166 507218 244250 507454
rect 244486 507218 244570 507454
rect 244806 507218 263930 507454
rect 264166 507218 264250 507454
rect 264486 507218 264570 507454
rect 264806 507218 283930 507454
rect 284166 507218 284250 507454
rect 284486 507218 284570 507454
rect 284806 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 483930 507454
rect 484166 507218 484250 507454
rect 484486 507218 484570 507454
rect 484806 507218 503930 507454
rect 504166 507218 504250 507454
rect 504486 507218 504570 507454
rect 504806 507218 523930 507454
rect 524166 507218 524250 507454
rect 524486 507218 524570 507454
rect 524806 507218 543930 507454
rect 544166 507218 544250 507454
rect 544486 507218 544570 507454
rect 544806 507218 563930 507454
rect 564166 507218 564250 507454
rect 564486 507218 564570 507454
rect 564806 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 203930 507134
rect 204166 506898 204250 507134
rect 204486 506898 204570 507134
rect 204806 506898 223930 507134
rect 224166 506898 224250 507134
rect 224486 506898 224570 507134
rect 224806 506898 243930 507134
rect 244166 506898 244250 507134
rect 244486 506898 244570 507134
rect 244806 506898 263930 507134
rect 264166 506898 264250 507134
rect 264486 506898 264570 507134
rect 264806 506898 283930 507134
rect 284166 506898 284250 507134
rect 284486 506898 284570 507134
rect 284806 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 483930 507134
rect 484166 506898 484250 507134
rect 484486 506898 484570 507134
rect 484806 506898 503930 507134
rect 504166 506898 504250 507134
rect 504486 506898 504570 507134
rect 504806 506898 523930 507134
rect 524166 506898 524250 507134
rect 524486 506898 524570 507134
rect 524806 506898 543930 507134
rect 544166 506898 544250 507134
rect 544486 506898 544570 507134
rect 544806 506898 563930 507134
rect 564166 506898 564250 507134
rect 564486 506898 564570 507134
rect 564806 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 213930 475954
rect 214166 475718 214250 475954
rect 214486 475718 214570 475954
rect 214806 475718 233930 475954
rect 234166 475718 234250 475954
rect 234486 475718 234570 475954
rect 234806 475718 253930 475954
rect 254166 475718 254250 475954
rect 254486 475718 254570 475954
rect 254806 475718 273930 475954
rect 274166 475718 274250 475954
rect 274486 475718 274570 475954
rect 274806 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 493930 475954
rect 494166 475718 494250 475954
rect 494486 475718 494570 475954
rect 494806 475718 513930 475954
rect 514166 475718 514250 475954
rect 514486 475718 514570 475954
rect 514806 475718 533930 475954
rect 534166 475718 534250 475954
rect 534486 475718 534570 475954
rect 534806 475718 553930 475954
rect 554166 475718 554250 475954
rect 554486 475718 554570 475954
rect 554806 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 213930 475634
rect 214166 475398 214250 475634
rect 214486 475398 214570 475634
rect 214806 475398 233930 475634
rect 234166 475398 234250 475634
rect 234486 475398 234570 475634
rect 234806 475398 253930 475634
rect 254166 475398 254250 475634
rect 254486 475398 254570 475634
rect 254806 475398 273930 475634
rect 274166 475398 274250 475634
rect 274486 475398 274570 475634
rect 274806 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 493930 475634
rect 494166 475398 494250 475634
rect 494486 475398 494570 475634
rect 494806 475398 513930 475634
rect 514166 475398 514250 475634
rect 514486 475398 514570 475634
rect 514806 475398 533930 475634
rect 534166 475398 534250 475634
rect 534486 475398 534570 475634
rect 534806 475398 553930 475634
rect 554166 475398 554250 475634
rect 554486 475398 554570 475634
rect 554806 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 203930 471454
rect 204166 471218 204250 471454
rect 204486 471218 204570 471454
rect 204806 471218 223930 471454
rect 224166 471218 224250 471454
rect 224486 471218 224570 471454
rect 224806 471218 243930 471454
rect 244166 471218 244250 471454
rect 244486 471218 244570 471454
rect 244806 471218 263930 471454
rect 264166 471218 264250 471454
rect 264486 471218 264570 471454
rect 264806 471218 283930 471454
rect 284166 471218 284250 471454
rect 284486 471218 284570 471454
rect 284806 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 483930 471454
rect 484166 471218 484250 471454
rect 484486 471218 484570 471454
rect 484806 471218 503930 471454
rect 504166 471218 504250 471454
rect 504486 471218 504570 471454
rect 504806 471218 523930 471454
rect 524166 471218 524250 471454
rect 524486 471218 524570 471454
rect 524806 471218 543930 471454
rect 544166 471218 544250 471454
rect 544486 471218 544570 471454
rect 544806 471218 563930 471454
rect 564166 471218 564250 471454
rect 564486 471218 564570 471454
rect 564806 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 203930 471134
rect 204166 470898 204250 471134
rect 204486 470898 204570 471134
rect 204806 470898 223930 471134
rect 224166 470898 224250 471134
rect 224486 470898 224570 471134
rect 224806 470898 243930 471134
rect 244166 470898 244250 471134
rect 244486 470898 244570 471134
rect 244806 470898 263930 471134
rect 264166 470898 264250 471134
rect 264486 470898 264570 471134
rect 264806 470898 283930 471134
rect 284166 470898 284250 471134
rect 284486 470898 284570 471134
rect 284806 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 483930 471134
rect 484166 470898 484250 471134
rect 484486 470898 484570 471134
rect 484806 470898 503930 471134
rect 504166 470898 504250 471134
rect 504486 470898 504570 471134
rect 504806 470898 523930 471134
rect 524166 470898 524250 471134
rect 524486 470898 524570 471134
rect 524806 470898 543930 471134
rect 544166 470898 544250 471134
rect 544486 470898 544570 471134
rect 544806 470898 563930 471134
rect 564166 470898 564250 471134
rect 564486 470898 564570 471134
rect 564806 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 213930 439954
rect 214166 439718 214250 439954
rect 214486 439718 214570 439954
rect 214806 439718 233930 439954
rect 234166 439718 234250 439954
rect 234486 439718 234570 439954
rect 234806 439718 253930 439954
rect 254166 439718 254250 439954
rect 254486 439718 254570 439954
rect 254806 439718 273930 439954
rect 274166 439718 274250 439954
rect 274486 439718 274570 439954
rect 274806 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 493930 439954
rect 494166 439718 494250 439954
rect 494486 439718 494570 439954
rect 494806 439718 513930 439954
rect 514166 439718 514250 439954
rect 514486 439718 514570 439954
rect 514806 439718 533930 439954
rect 534166 439718 534250 439954
rect 534486 439718 534570 439954
rect 534806 439718 553930 439954
rect 554166 439718 554250 439954
rect 554486 439718 554570 439954
rect 554806 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 213930 439634
rect 214166 439398 214250 439634
rect 214486 439398 214570 439634
rect 214806 439398 233930 439634
rect 234166 439398 234250 439634
rect 234486 439398 234570 439634
rect 234806 439398 253930 439634
rect 254166 439398 254250 439634
rect 254486 439398 254570 439634
rect 254806 439398 273930 439634
rect 274166 439398 274250 439634
rect 274486 439398 274570 439634
rect 274806 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 493930 439634
rect 494166 439398 494250 439634
rect 494486 439398 494570 439634
rect 494806 439398 513930 439634
rect 514166 439398 514250 439634
rect 514486 439398 514570 439634
rect 514806 439398 533930 439634
rect 534166 439398 534250 439634
rect 534486 439398 534570 439634
rect 534806 439398 553930 439634
rect 554166 439398 554250 439634
rect 554486 439398 554570 439634
rect 554806 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 203930 435454
rect 204166 435218 204250 435454
rect 204486 435218 204570 435454
rect 204806 435218 223930 435454
rect 224166 435218 224250 435454
rect 224486 435218 224570 435454
rect 224806 435218 243930 435454
rect 244166 435218 244250 435454
rect 244486 435218 244570 435454
rect 244806 435218 263930 435454
rect 264166 435218 264250 435454
rect 264486 435218 264570 435454
rect 264806 435218 283930 435454
rect 284166 435218 284250 435454
rect 284486 435218 284570 435454
rect 284806 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 483930 435454
rect 484166 435218 484250 435454
rect 484486 435218 484570 435454
rect 484806 435218 503930 435454
rect 504166 435218 504250 435454
rect 504486 435218 504570 435454
rect 504806 435218 523930 435454
rect 524166 435218 524250 435454
rect 524486 435218 524570 435454
rect 524806 435218 543930 435454
rect 544166 435218 544250 435454
rect 544486 435218 544570 435454
rect 544806 435218 563930 435454
rect 564166 435218 564250 435454
rect 564486 435218 564570 435454
rect 564806 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 203930 435134
rect 204166 434898 204250 435134
rect 204486 434898 204570 435134
rect 204806 434898 223930 435134
rect 224166 434898 224250 435134
rect 224486 434898 224570 435134
rect 224806 434898 243930 435134
rect 244166 434898 244250 435134
rect 244486 434898 244570 435134
rect 244806 434898 263930 435134
rect 264166 434898 264250 435134
rect 264486 434898 264570 435134
rect 264806 434898 283930 435134
rect 284166 434898 284250 435134
rect 284486 434898 284570 435134
rect 284806 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 483930 435134
rect 484166 434898 484250 435134
rect 484486 434898 484570 435134
rect 484806 434898 503930 435134
rect 504166 434898 504250 435134
rect 504486 434898 504570 435134
rect 504806 434898 523930 435134
rect 524166 434898 524250 435134
rect 524486 434898 524570 435134
rect 524806 434898 543930 435134
rect 544166 434898 544250 435134
rect 544486 434898 544570 435134
rect 544806 434898 563930 435134
rect 564166 434898 564250 435134
rect 564486 434898 564570 435134
rect 564806 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 213930 403954
rect 214166 403718 214250 403954
rect 214486 403718 214570 403954
rect 214806 403718 233930 403954
rect 234166 403718 234250 403954
rect 234486 403718 234570 403954
rect 234806 403718 253930 403954
rect 254166 403718 254250 403954
rect 254486 403718 254570 403954
rect 254806 403718 273930 403954
rect 274166 403718 274250 403954
rect 274486 403718 274570 403954
rect 274806 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 493930 403954
rect 494166 403718 494250 403954
rect 494486 403718 494570 403954
rect 494806 403718 513930 403954
rect 514166 403718 514250 403954
rect 514486 403718 514570 403954
rect 514806 403718 533930 403954
rect 534166 403718 534250 403954
rect 534486 403718 534570 403954
rect 534806 403718 553930 403954
rect 554166 403718 554250 403954
rect 554486 403718 554570 403954
rect 554806 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 213930 403634
rect 214166 403398 214250 403634
rect 214486 403398 214570 403634
rect 214806 403398 233930 403634
rect 234166 403398 234250 403634
rect 234486 403398 234570 403634
rect 234806 403398 253930 403634
rect 254166 403398 254250 403634
rect 254486 403398 254570 403634
rect 254806 403398 273930 403634
rect 274166 403398 274250 403634
rect 274486 403398 274570 403634
rect 274806 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 493930 403634
rect 494166 403398 494250 403634
rect 494486 403398 494570 403634
rect 494806 403398 513930 403634
rect 514166 403398 514250 403634
rect 514486 403398 514570 403634
rect 514806 403398 533930 403634
rect 534166 403398 534250 403634
rect 534486 403398 534570 403634
rect 534806 403398 553930 403634
rect 554166 403398 554250 403634
rect 554486 403398 554570 403634
rect 554806 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 203930 399454
rect 204166 399218 204250 399454
rect 204486 399218 204570 399454
rect 204806 399218 223930 399454
rect 224166 399218 224250 399454
rect 224486 399218 224570 399454
rect 224806 399218 243930 399454
rect 244166 399218 244250 399454
rect 244486 399218 244570 399454
rect 244806 399218 263930 399454
rect 264166 399218 264250 399454
rect 264486 399218 264570 399454
rect 264806 399218 283930 399454
rect 284166 399218 284250 399454
rect 284486 399218 284570 399454
rect 284806 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 483930 399454
rect 484166 399218 484250 399454
rect 484486 399218 484570 399454
rect 484806 399218 503930 399454
rect 504166 399218 504250 399454
rect 504486 399218 504570 399454
rect 504806 399218 523930 399454
rect 524166 399218 524250 399454
rect 524486 399218 524570 399454
rect 524806 399218 543930 399454
rect 544166 399218 544250 399454
rect 544486 399218 544570 399454
rect 544806 399218 563930 399454
rect 564166 399218 564250 399454
rect 564486 399218 564570 399454
rect 564806 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 203930 399134
rect 204166 398898 204250 399134
rect 204486 398898 204570 399134
rect 204806 398898 223930 399134
rect 224166 398898 224250 399134
rect 224486 398898 224570 399134
rect 224806 398898 243930 399134
rect 244166 398898 244250 399134
rect 244486 398898 244570 399134
rect 244806 398898 263930 399134
rect 264166 398898 264250 399134
rect 264486 398898 264570 399134
rect 264806 398898 283930 399134
rect 284166 398898 284250 399134
rect 284486 398898 284570 399134
rect 284806 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 483930 399134
rect 484166 398898 484250 399134
rect 484486 398898 484570 399134
rect 484806 398898 503930 399134
rect 504166 398898 504250 399134
rect 504486 398898 504570 399134
rect 504806 398898 523930 399134
rect 524166 398898 524250 399134
rect 524486 398898 524570 399134
rect 524806 398898 543930 399134
rect 544166 398898 544250 399134
rect 544486 398898 544570 399134
rect 544806 398898 563930 399134
rect 564166 398898 564250 399134
rect 564486 398898 564570 399134
rect 564806 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 213930 367954
rect 214166 367718 214250 367954
rect 214486 367718 214570 367954
rect 214806 367718 233930 367954
rect 234166 367718 234250 367954
rect 234486 367718 234570 367954
rect 234806 367718 253930 367954
rect 254166 367718 254250 367954
rect 254486 367718 254570 367954
rect 254806 367718 273930 367954
rect 274166 367718 274250 367954
rect 274486 367718 274570 367954
rect 274806 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 493930 367954
rect 494166 367718 494250 367954
rect 494486 367718 494570 367954
rect 494806 367718 513930 367954
rect 514166 367718 514250 367954
rect 514486 367718 514570 367954
rect 514806 367718 533930 367954
rect 534166 367718 534250 367954
rect 534486 367718 534570 367954
rect 534806 367718 553930 367954
rect 554166 367718 554250 367954
rect 554486 367718 554570 367954
rect 554806 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 213930 367634
rect 214166 367398 214250 367634
rect 214486 367398 214570 367634
rect 214806 367398 233930 367634
rect 234166 367398 234250 367634
rect 234486 367398 234570 367634
rect 234806 367398 253930 367634
rect 254166 367398 254250 367634
rect 254486 367398 254570 367634
rect 254806 367398 273930 367634
rect 274166 367398 274250 367634
rect 274486 367398 274570 367634
rect 274806 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 493930 367634
rect 494166 367398 494250 367634
rect 494486 367398 494570 367634
rect 494806 367398 513930 367634
rect 514166 367398 514250 367634
rect 514486 367398 514570 367634
rect 514806 367398 533930 367634
rect 534166 367398 534250 367634
rect 534486 367398 534570 367634
rect 534806 367398 553930 367634
rect 554166 367398 554250 367634
rect 554486 367398 554570 367634
rect 554806 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 203930 363454
rect 204166 363218 204250 363454
rect 204486 363218 204570 363454
rect 204806 363218 223930 363454
rect 224166 363218 224250 363454
rect 224486 363218 224570 363454
rect 224806 363218 243930 363454
rect 244166 363218 244250 363454
rect 244486 363218 244570 363454
rect 244806 363218 263930 363454
rect 264166 363218 264250 363454
rect 264486 363218 264570 363454
rect 264806 363218 283930 363454
rect 284166 363218 284250 363454
rect 284486 363218 284570 363454
rect 284806 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 483930 363454
rect 484166 363218 484250 363454
rect 484486 363218 484570 363454
rect 484806 363218 503930 363454
rect 504166 363218 504250 363454
rect 504486 363218 504570 363454
rect 504806 363218 523930 363454
rect 524166 363218 524250 363454
rect 524486 363218 524570 363454
rect 524806 363218 543930 363454
rect 544166 363218 544250 363454
rect 544486 363218 544570 363454
rect 544806 363218 563930 363454
rect 564166 363218 564250 363454
rect 564486 363218 564570 363454
rect 564806 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 203930 363134
rect 204166 362898 204250 363134
rect 204486 362898 204570 363134
rect 204806 362898 223930 363134
rect 224166 362898 224250 363134
rect 224486 362898 224570 363134
rect 224806 362898 243930 363134
rect 244166 362898 244250 363134
rect 244486 362898 244570 363134
rect 244806 362898 263930 363134
rect 264166 362898 264250 363134
rect 264486 362898 264570 363134
rect 264806 362898 283930 363134
rect 284166 362898 284250 363134
rect 284486 362898 284570 363134
rect 284806 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 483930 363134
rect 484166 362898 484250 363134
rect 484486 362898 484570 363134
rect 484806 362898 503930 363134
rect 504166 362898 504250 363134
rect 504486 362898 504570 363134
rect 504806 362898 523930 363134
rect 524166 362898 524250 363134
rect 524486 362898 524570 363134
rect 524806 362898 543930 363134
rect 544166 362898 544250 363134
rect 544486 362898 544570 363134
rect 544806 362898 563930 363134
rect 564166 362898 564250 363134
rect 564486 362898 564570 363134
rect 564806 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 213930 295954
rect 214166 295718 214250 295954
rect 214486 295718 214570 295954
rect 214806 295718 233930 295954
rect 234166 295718 234250 295954
rect 234486 295718 234570 295954
rect 234806 295718 253930 295954
rect 254166 295718 254250 295954
rect 254486 295718 254570 295954
rect 254806 295718 273930 295954
rect 274166 295718 274250 295954
rect 274486 295718 274570 295954
rect 274806 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 493930 295954
rect 494166 295718 494250 295954
rect 494486 295718 494570 295954
rect 494806 295718 513930 295954
rect 514166 295718 514250 295954
rect 514486 295718 514570 295954
rect 514806 295718 533930 295954
rect 534166 295718 534250 295954
rect 534486 295718 534570 295954
rect 534806 295718 553930 295954
rect 554166 295718 554250 295954
rect 554486 295718 554570 295954
rect 554806 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 213930 295634
rect 214166 295398 214250 295634
rect 214486 295398 214570 295634
rect 214806 295398 233930 295634
rect 234166 295398 234250 295634
rect 234486 295398 234570 295634
rect 234806 295398 253930 295634
rect 254166 295398 254250 295634
rect 254486 295398 254570 295634
rect 254806 295398 273930 295634
rect 274166 295398 274250 295634
rect 274486 295398 274570 295634
rect 274806 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 493930 295634
rect 494166 295398 494250 295634
rect 494486 295398 494570 295634
rect 494806 295398 513930 295634
rect 514166 295398 514250 295634
rect 514486 295398 514570 295634
rect 514806 295398 533930 295634
rect 534166 295398 534250 295634
rect 534486 295398 534570 295634
rect 534806 295398 553930 295634
rect 554166 295398 554250 295634
rect 554486 295398 554570 295634
rect 554806 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 203930 291454
rect 204166 291218 204250 291454
rect 204486 291218 204570 291454
rect 204806 291218 223930 291454
rect 224166 291218 224250 291454
rect 224486 291218 224570 291454
rect 224806 291218 243930 291454
rect 244166 291218 244250 291454
rect 244486 291218 244570 291454
rect 244806 291218 263930 291454
rect 264166 291218 264250 291454
rect 264486 291218 264570 291454
rect 264806 291218 283930 291454
rect 284166 291218 284250 291454
rect 284486 291218 284570 291454
rect 284806 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 483930 291454
rect 484166 291218 484250 291454
rect 484486 291218 484570 291454
rect 484806 291218 503930 291454
rect 504166 291218 504250 291454
rect 504486 291218 504570 291454
rect 504806 291218 523930 291454
rect 524166 291218 524250 291454
rect 524486 291218 524570 291454
rect 524806 291218 543930 291454
rect 544166 291218 544250 291454
rect 544486 291218 544570 291454
rect 544806 291218 563930 291454
rect 564166 291218 564250 291454
rect 564486 291218 564570 291454
rect 564806 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 203930 291134
rect 204166 290898 204250 291134
rect 204486 290898 204570 291134
rect 204806 290898 223930 291134
rect 224166 290898 224250 291134
rect 224486 290898 224570 291134
rect 224806 290898 243930 291134
rect 244166 290898 244250 291134
rect 244486 290898 244570 291134
rect 244806 290898 263930 291134
rect 264166 290898 264250 291134
rect 264486 290898 264570 291134
rect 264806 290898 283930 291134
rect 284166 290898 284250 291134
rect 284486 290898 284570 291134
rect 284806 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 483930 291134
rect 484166 290898 484250 291134
rect 484486 290898 484570 291134
rect 484806 290898 503930 291134
rect 504166 290898 504250 291134
rect 504486 290898 504570 291134
rect 504806 290898 523930 291134
rect 524166 290898 524250 291134
rect 524486 290898 524570 291134
rect 524806 290898 543930 291134
rect 544166 290898 544250 291134
rect 544486 290898 544570 291134
rect 544806 290898 563930 291134
rect 564166 290898 564250 291134
rect 564486 290898 564570 291134
rect 564806 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 213930 259954
rect 214166 259718 214250 259954
rect 214486 259718 214570 259954
rect 214806 259718 233930 259954
rect 234166 259718 234250 259954
rect 234486 259718 234570 259954
rect 234806 259718 253930 259954
rect 254166 259718 254250 259954
rect 254486 259718 254570 259954
rect 254806 259718 273930 259954
rect 274166 259718 274250 259954
rect 274486 259718 274570 259954
rect 274806 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 493930 259954
rect 494166 259718 494250 259954
rect 494486 259718 494570 259954
rect 494806 259718 513930 259954
rect 514166 259718 514250 259954
rect 514486 259718 514570 259954
rect 514806 259718 533930 259954
rect 534166 259718 534250 259954
rect 534486 259718 534570 259954
rect 534806 259718 553930 259954
rect 554166 259718 554250 259954
rect 554486 259718 554570 259954
rect 554806 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 213930 259634
rect 214166 259398 214250 259634
rect 214486 259398 214570 259634
rect 214806 259398 233930 259634
rect 234166 259398 234250 259634
rect 234486 259398 234570 259634
rect 234806 259398 253930 259634
rect 254166 259398 254250 259634
rect 254486 259398 254570 259634
rect 254806 259398 273930 259634
rect 274166 259398 274250 259634
rect 274486 259398 274570 259634
rect 274806 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 493930 259634
rect 494166 259398 494250 259634
rect 494486 259398 494570 259634
rect 494806 259398 513930 259634
rect 514166 259398 514250 259634
rect 514486 259398 514570 259634
rect 514806 259398 533930 259634
rect 534166 259398 534250 259634
rect 534486 259398 534570 259634
rect 534806 259398 553930 259634
rect 554166 259398 554250 259634
rect 554486 259398 554570 259634
rect 554806 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 203930 255454
rect 204166 255218 204250 255454
rect 204486 255218 204570 255454
rect 204806 255218 223930 255454
rect 224166 255218 224250 255454
rect 224486 255218 224570 255454
rect 224806 255218 243930 255454
rect 244166 255218 244250 255454
rect 244486 255218 244570 255454
rect 244806 255218 263930 255454
rect 264166 255218 264250 255454
rect 264486 255218 264570 255454
rect 264806 255218 283930 255454
rect 284166 255218 284250 255454
rect 284486 255218 284570 255454
rect 284806 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 483930 255454
rect 484166 255218 484250 255454
rect 484486 255218 484570 255454
rect 484806 255218 503930 255454
rect 504166 255218 504250 255454
rect 504486 255218 504570 255454
rect 504806 255218 523930 255454
rect 524166 255218 524250 255454
rect 524486 255218 524570 255454
rect 524806 255218 543930 255454
rect 544166 255218 544250 255454
rect 544486 255218 544570 255454
rect 544806 255218 563930 255454
rect 564166 255218 564250 255454
rect 564486 255218 564570 255454
rect 564806 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 203930 255134
rect 204166 254898 204250 255134
rect 204486 254898 204570 255134
rect 204806 254898 223930 255134
rect 224166 254898 224250 255134
rect 224486 254898 224570 255134
rect 224806 254898 243930 255134
rect 244166 254898 244250 255134
rect 244486 254898 244570 255134
rect 244806 254898 263930 255134
rect 264166 254898 264250 255134
rect 264486 254898 264570 255134
rect 264806 254898 283930 255134
rect 284166 254898 284250 255134
rect 284486 254898 284570 255134
rect 284806 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 483930 255134
rect 484166 254898 484250 255134
rect 484486 254898 484570 255134
rect 484806 254898 503930 255134
rect 504166 254898 504250 255134
rect 504486 254898 504570 255134
rect 504806 254898 523930 255134
rect 524166 254898 524250 255134
rect 524486 254898 524570 255134
rect 524806 254898 543930 255134
rect 544166 254898 544250 255134
rect 544486 254898 544570 255134
rect 544806 254898 563930 255134
rect 564166 254898 564250 255134
rect 564486 254898 564570 255134
rect 564806 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 213930 223954
rect 214166 223718 214250 223954
rect 214486 223718 214570 223954
rect 214806 223718 233930 223954
rect 234166 223718 234250 223954
rect 234486 223718 234570 223954
rect 234806 223718 253930 223954
rect 254166 223718 254250 223954
rect 254486 223718 254570 223954
rect 254806 223718 273930 223954
rect 274166 223718 274250 223954
rect 274486 223718 274570 223954
rect 274806 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 493930 223954
rect 494166 223718 494250 223954
rect 494486 223718 494570 223954
rect 494806 223718 513930 223954
rect 514166 223718 514250 223954
rect 514486 223718 514570 223954
rect 514806 223718 533930 223954
rect 534166 223718 534250 223954
rect 534486 223718 534570 223954
rect 534806 223718 553930 223954
rect 554166 223718 554250 223954
rect 554486 223718 554570 223954
rect 554806 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 213930 223634
rect 214166 223398 214250 223634
rect 214486 223398 214570 223634
rect 214806 223398 233930 223634
rect 234166 223398 234250 223634
rect 234486 223398 234570 223634
rect 234806 223398 253930 223634
rect 254166 223398 254250 223634
rect 254486 223398 254570 223634
rect 254806 223398 273930 223634
rect 274166 223398 274250 223634
rect 274486 223398 274570 223634
rect 274806 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 493930 223634
rect 494166 223398 494250 223634
rect 494486 223398 494570 223634
rect 494806 223398 513930 223634
rect 514166 223398 514250 223634
rect 514486 223398 514570 223634
rect 514806 223398 533930 223634
rect 534166 223398 534250 223634
rect 534486 223398 534570 223634
rect 534806 223398 553930 223634
rect 554166 223398 554250 223634
rect 554486 223398 554570 223634
rect 554806 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 203930 219454
rect 204166 219218 204250 219454
rect 204486 219218 204570 219454
rect 204806 219218 223930 219454
rect 224166 219218 224250 219454
rect 224486 219218 224570 219454
rect 224806 219218 243930 219454
rect 244166 219218 244250 219454
rect 244486 219218 244570 219454
rect 244806 219218 263930 219454
rect 264166 219218 264250 219454
rect 264486 219218 264570 219454
rect 264806 219218 283930 219454
rect 284166 219218 284250 219454
rect 284486 219218 284570 219454
rect 284806 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 483930 219454
rect 484166 219218 484250 219454
rect 484486 219218 484570 219454
rect 484806 219218 503930 219454
rect 504166 219218 504250 219454
rect 504486 219218 504570 219454
rect 504806 219218 523930 219454
rect 524166 219218 524250 219454
rect 524486 219218 524570 219454
rect 524806 219218 543930 219454
rect 544166 219218 544250 219454
rect 544486 219218 544570 219454
rect 544806 219218 563930 219454
rect 564166 219218 564250 219454
rect 564486 219218 564570 219454
rect 564806 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 203930 219134
rect 204166 218898 204250 219134
rect 204486 218898 204570 219134
rect 204806 218898 223930 219134
rect 224166 218898 224250 219134
rect 224486 218898 224570 219134
rect 224806 218898 243930 219134
rect 244166 218898 244250 219134
rect 244486 218898 244570 219134
rect 244806 218898 263930 219134
rect 264166 218898 264250 219134
rect 264486 218898 264570 219134
rect 264806 218898 283930 219134
rect 284166 218898 284250 219134
rect 284486 218898 284570 219134
rect 284806 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 483930 219134
rect 484166 218898 484250 219134
rect 484486 218898 484570 219134
rect 484806 218898 503930 219134
rect 504166 218898 504250 219134
rect 504486 218898 504570 219134
rect 504806 218898 523930 219134
rect 524166 218898 524250 219134
rect 524486 218898 524570 219134
rect 524806 218898 543930 219134
rect 544166 218898 544250 219134
rect 544486 218898 544570 219134
rect 544806 218898 563930 219134
rect 564166 218898 564250 219134
rect 564486 218898 564570 219134
rect 564806 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 203930 183454
rect 204166 183218 204250 183454
rect 204486 183218 204570 183454
rect 204806 183218 223930 183454
rect 224166 183218 224250 183454
rect 224486 183218 224570 183454
rect 224806 183218 243930 183454
rect 244166 183218 244250 183454
rect 244486 183218 244570 183454
rect 244806 183218 263930 183454
rect 264166 183218 264250 183454
rect 264486 183218 264570 183454
rect 264806 183218 283930 183454
rect 284166 183218 284250 183454
rect 284486 183218 284570 183454
rect 284806 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 483930 183454
rect 484166 183218 484250 183454
rect 484486 183218 484570 183454
rect 484806 183218 503930 183454
rect 504166 183218 504250 183454
rect 504486 183218 504570 183454
rect 504806 183218 523930 183454
rect 524166 183218 524250 183454
rect 524486 183218 524570 183454
rect 524806 183218 543930 183454
rect 544166 183218 544250 183454
rect 544486 183218 544570 183454
rect 544806 183218 563930 183454
rect 564166 183218 564250 183454
rect 564486 183218 564570 183454
rect 564806 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 203930 183134
rect 204166 182898 204250 183134
rect 204486 182898 204570 183134
rect 204806 182898 223930 183134
rect 224166 182898 224250 183134
rect 224486 182898 224570 183134
rect 224806 182898 243930 183134
rect 244166 182898 244250 183134
rect 244486 182898 244570 183134
rect 244806 182898 263930 183134
rect 264166 182898 264250 183134
rect 264486 182898 264570 183134
rect 264806 182898 283930 183134
rect 284166 182898 284250 183134
rect 284486 182898 284570 183134
rect 284806 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 483930 183134
rect 484166 182898 484250 183134
rect 484486 182898 484570 183134
rect 484806 182898 503930 183134
rect 504166 182898 504250 183134
rect 504486 182898 504570 183134
rect 504806 182898 523930 183134
rect 524166 182898 524250 183134
rect 524486 182898 524570 183134
rect 524806 182898 543930 183134
rect 544166 182898 544250 183134
rect 544486 182898 544570 183134
rect 544806 182898 563930 183134
rect 564166 182898 564250 183134
rect 564486 182898 564570 183134
rect 564806 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 213930 151954
rect 214166 151718 214250 151954
rect 214486 151718 214570 151954
rect 214806 151718 233930 151954
rect 234166 151718 234250 151954
rect 234486 151718 234570 151954
rect 234806 151718 253930 151954
rect 254166 151718 254250 151954
rect 254486 151718 254570 151954
rect 254806 151718 273930 151954
rect 274166 151718 274250 151954
rect 274486 151718 274570 151954
rect 274806 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 493930 151954
rect 494166 151718 494250 151954
rect 494486 151718 494570 151954
rect 494806 151718 513930 151954
rect 514166 151718 514250 151954
rect 514486 151718 514570 151954
rect 514806 151718 533930 151954
rect 534166 151718 534250 151954
rect 534486 151718 534570 151954
rect 534806 151718 553930 151954
rect 554166 151718 554250 151954
rect 554486 151718 554570 151954
rect 554806 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 213930 151634
rect 214166 151398 214250 151634
rect 214486 151398 214570 151634
rect 214806 151398 233930 151634
rect 234166 151398 234250 151634
rect 234486 151398 234570 151634
rect 234806 151398 253930 151634
rect 254166 151398 254250 151634
rect 254486 151398 254570 151634
rect 254806 151398 273930 151634
rect 274166 151398 274250 151634
rect 274486 151398 274570 151634
rect 274806 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 493930 151634
rect 494166 151398 494250 151634
rect 494486 151398 494570 151634
rect 494806 151398 513930 151634
rect 514166 151398 514250 151634
rect 514486 151398 514570 151634
rect 514806 151398 533930 151634
rect 534166 151398 534250 151634
rect 534486 151398 534570 151634
rect 534806 151398 553930 151634
rect 554166 151398 554250 151634
rect 554486 151398 554570 151634
rect 554806 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 203930 147454
rect 204166 147218 204250 147454
rect 204486 147218 204570 147454
rect 204806 147218 223930 147454
rect 224166 147218 224250 147454
rect 224486 147218 224570 147454
rect 224806 147218 243930 147454
rect 244166 147218 244250 147454
rect 244486 147218 244570 147454
rect 244806 147218 263930 147454
rect 264166 147218 264250 147454
rect 264486 147218 264570 147454
rect 264806 147218 283930 147454
rect 284166 147218 284250 147454
rect 284486 147218 284570 147454
rect 284806 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 483930 147454
rect 484166 147218 484250 147454
rect 484486 147218 484570 147454
rect 484806 147218 503930 147454
rect 504166 147218 504250 147454
rect 504486 147218 504570 147454
rect 504806 147218 523930 147454
rect 524166 147218 524250 147454
rect 524486 147218 524570 147454
rect 524806 147218 543930 147454
rect 544166 147218 544250 147454
rect 544486 147218 544570 147454
rect 544806 147218 563930 147454
rect 564166 147218 564250 147454
rect 564486 147218 564570 147454
rect 564806 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 203930 147134
rect 204166 146898 204250 147134
rect 204486 146898 204570 147134
rect 204806 146898 223930 147134
rect 224166 146898 224250 147134
rect 224486 146898 224570 147134
rect 224806 146898 243930 147134
rect 244166 146898 244250 147134
rect 244486 146898 244570 147134
rect 244806 146898 263930 147134
rect 264166 146898 264250 147134
rect 264486 146898 264570 147134
rect 264806 146898 283930 147134
rect 284166 146898 284250 147134
rect 284486 146898 284570 147134
rect 284806 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 483930 147134
rect 484166 146898 484250 147134
rect 484486 146898 484570 147134
rect 484806 146898 503930 147134
rect 504166 146898 504250 147134
rect 504486 146898 504570 147134
rect 504806 146898 523930 147134
rect 524166 146898 524250 147134
rect 524486 146898 524570 147134
rect 524806 146898 543930 147134
rect 544166 146898 544250 147134
rect 544486 146898 544570 147134
rect 544806 146898 563930 147134
rect 564166 146898 564250 147134
rect 564486 146898 564570 147134
rect 564806 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 213930 115954
rect 214166 115718 214250 115954
rect 214486 115718 214570 115954
rect 214806 115718 233930 115954
rect 234166 115718 234250 115954
rect 234486 115718 234570 115954
rect 234806 115718 253930 115954
rect 254166 115718 254250 115954
rect 254486 115718 254570 115954
rect 254806 115718 273930 115954
rect 274166 115718 274250 115954
rect 274486 115718 274570 115954
rect 274806 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 493930 115954
rect 494166 115718 494250 115954
rect 494486 115718 494570 115954
rect 494806 115718 513930 115954
rect 514166 115718 514250 115954
rect 514486 115718 514570 115954
rect 514806 115718 533930 115954
rect 534166 115718 534250 115954
rect 534486 115718 534570 115954
rect 534806 115718 553930 115954
rect 554166 115718 554250 115954
rect 554486 115718 554570 115954
rect 554806 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 213930 115634
rect 214166 115398 214250 115634
rect 214486 115398 214570 115634
rect 214806 115398 233930 115634
rect 234166 115398 234250 115634
rect 234486 115398 234570 115634
rect 234806 115398 253930 115634
rect 254166 115398 254250 115634
rect 254486 115398 254570 115634
rect 254806 115398 273930 115634
rect 274166 115398 274250 115634
rect 274486 115398 274570 115634
rect 274806 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 493930 115634
rect 494166 115398 494250 115634
rect 494486 115398 494570 115634
rect 494806 115398 513930 115634
rect 514166 115398 514250 115634
rect 514486 115398 514570 115634
rect 514806 115398 533930 115634
rect 534166 115398 534250 115634
rect 534486 115398 534570 115634
rect 534806 115398 553930 115634
rect 554166 115398 554250 115634
rect 554486 115398 554570 115634
rect 554806 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 203930 111454
rect 204166 111218 204250 111454
rect 204486 111218 204570 111454
rect 204806 111218 223930 111454
rect 224166 111218 224250 111454
rect 224486 111218 224570 111454
rect 224806 111218 243930 111454
rect 244166 111218 244250 111454
rect 244486 111218 244570 111454
rect 244806 111218 263930 111454
rect 264166 111218 264250 111454
rect 264486 111218 264570 111454
rect 264806 111218 283930 111454
rect 284166 111218 284250 111454
rect 284486 111218 284570 111454
rect 284806 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 483930 111454
rect 484166 111218 484250 111454
rect 484486 111218 484570 111454
rect 484806 111218 503930 111454
rect 504166 111218 504250 111454
rect 504486 111218 504570 111454
rect 504806 111218 523930 111454
rect 524166 111218 524250 111454
rect 524486 111218 524570 111454
rect 524806 111218 543930 111454
rect 544166 111218 544250 111454
rect 544486 111218 544570 111454
rect 544806 111218 563930 111454
rect 564166 111218 564250 111454
rect 564486 111218 564570 111454
rect 564806 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 203930 111134
rect 204166 110898 204250 111134
rect 204486 110898 204570 111134
rect 204806 110898 223930 111134
rect 224166 110898 224250 111134
rect 224486 110898 224570 111134
rect 224806 110898 243930 111134
rect 244166 110898 244250 111134
rect 244486 110898 244570 111134
rect 244806 110898 263930 111134
rect 264166 110898 264250 111134
rect 264486 110898 264570 111134
rect 264806 110898 283930 111134
rect 284166 110898 284250 111134
rect 284486 110898 284570 111134
rect 284806 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 483930 111134
rect 484166 110898 484250 111134
rect 484486 110898 484570 111134
rect 484806 110898 503930 111134
rect 504166 110898 504250 111134
rect 504486 110898 504570 111134
rect 504806 110898 523930 111134
rect 524166 110898 524250 111134
rect 524486 110898 524570 111134
rect 524806 110898 543930 111134
rect 544166 110898 544250 111134
rect 544486 110898 544570 111134
rect 544806 110898 563930 111134
rect 564166 110898 564250 111134
rect 564486 110898 564570 111134
rect 564806 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 167930 43954
rect 168166 43718 168250 43954
rect 168486 43718 168570 43954
rect 168806 43718 187930 43954
rect 188166 43718 188250 43954
rect 188486 43718 188570 43954
rect 188806 43718 207930 43954
rect 208166 43718 208250 43954
rect 208486 43718 208570 43954
rect 208806 43718 227930 43954
rect 228166 43718 228250 43954
rect 228486 43718 228570 43954
rect 228806 43718 247930 43954
rect 248166 43718 248250 43954
rect 248486 43718 248570 43954
rect 248806 43718 267930 43954
rect 268166 43718 268250 43954
rect 268486 43718 268570 43954
rect 268806 43718 287930 43954
rect 288166 43718 288250 43954
rect 288486 43718 288570 43954
rect 288806 43718 307930 43954
rect 308166 43718 308250 43954
rect 308486 43718 308570 43954
rect 308806 43718 327930 43954
rect 328166 43718 328250 43954
rect 328486 43718 328570 43954
rect 328806 43718 347930 43954
rect 348166 43718 348250 43954
rect 348486 43718 348570 43954
rect 348806 43718 367930 43954
rect 368166 43718 368250 43954
rect 368486 43718 368570 43954
rect 368806 43718 387930 43954
rect 388166 43718 388250 43954
rect 388486 43718 388570 43954
rect 388806 43718 407930 43954
rect 408166 43718 408250 43954
rect 408486 43718 408570 43954
rect 408806 43718 427930 43954
rect 428166 43718 428250 43954
rect 428486 43718 428570 43954
rect 428806 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 167930 43634
rect 168166 43398 168250 43634
rect 168486 43398 168570 43634
rect 168806 43398 187930 43634
rect 188166 43398 188250 43634
rect 188486 43398 188570 43634
rect 188806 43398 207930 43634
rect 208166 43398 208250 43634
rect 208486 43398 208570 43634
rect 208806 43398 227930 43634
rect 228166 43398 228250 43634
rect 228486 43398 228570 43634
rect 228806 43398 247930 43634
rect 248166 43398 248250 43634
rect 248486 43398 248570 43634
rect 248806 43398 267930 43634
rect 268166 43398 268250 43634
rect 268486 43398 268570 43634
rect 268806 43398 287930 43634
rect 288166 43398 288250 43634
rect 288486 43398 288570 43634
rect 288806 43398 307930 43634
rect 308166 43398 308250 43634
rect 308486 43398 308570 43634
rect 308806 43398 327930 43634
rect 328166 43398 328250 43634
rect 328486 43398 328570 43634
rect 328806 43398 347930 43634
rect 348166 43398 348250 43634
rect 348486 43398 348570 43634
rect 348806 43398 367930 43634
rect 368166 43398 368250 43634
rect 368486 43398 368570 43634
rect 368806 43398 387930 43634
rect 388166 43398 388250 43634
rect 388486 43398 388570 43634
rect 388806 43398 407930 43634
rect 408166 43398 408250 43634
rect 408486 43398 408570 43634
rect 408806 43398 427930 43634
rect 428166 43398 428250 43634
rect 428486 43398 428570 43634
rect 428806 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 157930 39454
rect 158166 39218 158250 39454
rect 158486 39218 158570 39454
rect 158806 39218 177930 39454
rect 178166 39218 178250 39454
rect 178486 39218 178570 39454
rect 178806 39218 197930 39454
rect 198166 39218 198250 39454
rect 198486 39218 198570 39454
rect 198806 39218 217930 39454
rect 218166 39218 218250 39454
rect 218486 39218 218570 39454
rect 218806 39218 237930 39454
rect 238166 39218 238250 39454
rect 238486 39218 238570 39454
rect 238806 39218 257930 39454
rect 258166 39218 258250 39454
rect 258486 39218 258570 39454
rect 258806 39218 277930 39454
rect 278166 39218 278250 39454
rect 278486 39218 278570 39454
rect 278806 39218 297930 39454
rect 298166 39218 298250 39454
rect 298486 39218 298570 39454
rect 298806 39218 317930 39454
rect 318166 39218 318250 39454
rect 318486 39218 318570 39454
rect 318806 39218 337930 39454
rect 338166 39218 338250 39454
rect 338486 39218 338570 39454
rect 338806 39218 357930 39454
rect 358166 39218 358250 39454
rect 358486 39218 358570 39454
rect 358806 39218 377930 39454
rect 378166 39218 378250 39454
rect 378486 39218 378570 39454
rect 378806 39218 397930 39454
rect 398166 39218 398250 39454
rect 398486 39218 398570 39454
rect 398806 39218 417930 39454
rect 418166 39218 418250 39454
rect 418486 39218 418570 39454
rect 418806 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 157930 39134
rect 158166 38898 158250 39134
rect 158486 38898 158570 39134
rect 158806 38898 177930 39134
rect 178166 38898 178250 39134
rect 178486 38898 178570 39134
rect 178806 38898 197930 39134
rect 198166 38898 198250 39134
rect 198486 38898 198570 39134
rect 198806 38898 217930 39134
rect 218166 38898 218250 39134
rect 218486 38898 218570 39134
rect 218806 38898 237930 39134
rect 238166 38898 238250 39134
rect 238486 38898 238570 39134
rect 238806 38898 257930 39134
rect 258166 38898 258250 39134
rect 258486 38898 258570 39134
rect 258806 38898 277930 39134
rect 278166 38898 278250 39134
rect 278486 38898 278570 39134
rect 278806 38898 297930 39134
rect 298166 38898 298250 39134
rect 298486 38898 298570 39134
rect 298806 38898 317930 39134
rect 318166 38898 318250 39134
rect 318486 38898 318570 39134
rect 318806 38898 337930 39134
rect 338166 38898 338250 39134
rect 338486 38898 338570 39134
rect 338806 38898 357930 39134
rect 358166 38898 358250 39134
rect 358486 38898 358570 39134
rect 358806 38898 377930 39134
rect 378166 38898 378250 39134
rect 378486 38898 378570 39134
rect 378806 38898 397930 39134
rect 398166 38898 398250 39134
rect 398486 38898 398570 39134
rect 398806 38898 417930 39134
rect 418166 38898 418250 39134
rect 418486 38898 418570 39134
rect 418806 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use controller_unit  controller_unit_mod
timestamp 0
transform 1 0 154000 0 1 24000
box -800 -800 280800 28800
use driver_core  driver_core_0
timestamp 0
transform 1 0 20000 0 1 78000
box 1066 -800 268862 107760
use driver_core  driver_core_1
timestamp 0
transform 1 0 20000 0 1 206000
box 1066 -800 268862 107760
use driver_core  driver_core_2
timestamp 0
transform 1 0 20000 0 1 334000
box 1066 -800 268862 107760
use driver_core  driver_core_3
timestamp 0
transform 1 0 20000 0 1 462000
box 1066 -800 268862 107760
use driver_core  driver_core_4
timestamp 0
transform 1 0 20000 0 1 588000
box 1066 -800 268862 107760
use driver_core  driver_core_5
timestamp 0
transform 1 0 300000 0 1 588000
box 1066 -800 268862 107760
use driver_core  driver_core_6
timestamp 0
transform 1 0 300000 0 1 462000
box 1066 -800 268862 107760
use driver_core  driver_core_7
timestamp 0
transform 1 0 300000 0 1 334000
box 1066 -800 268862 107760
use driver_core  driver_core_8
timestamp 0
transform 1 0 300000 0 1 206000
box 1066 -800 268862 107760
use driver_core  driver_core_9
timestamp 0
transform 1 0 300000 0 1 78000
box 1066 -800 268862 107760
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 54000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 700000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 700000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 700000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 700000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 700000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 700000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 700000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 700000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 700000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 700000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 700000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 700000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 700000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 700000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 700000 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
