VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO driver_core
  CLASS BLOCK ;
  FOREIGN driver_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 550.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 -4.000 382.630 4.000 ;
    END
  END clock
  PIN clock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 -4.000 363.310 4.000 ;
    END
  END clock_a
  PIN col_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 -4.000 730.390 4.000 ;
    END
  END col_select_a[0]
  PIN col_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 -4.000 749.710 4.000 ;
    END
  END col_select_a[1]
  PIN col_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 -4.000 769.030 4.000 ;
    END
  END col_select_a[2]
  PIN col_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 -4.000 788.350 4.000 ;
    END
  END col_select_a[3]
  PIN col_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 -4.000 807.670 4.000 ;
    END
  END col_select_a[4]
  PIN col_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 -4.000 826.990 4.000 ;
    END
  END col_select_a[5]
  PIN data_in_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -4.000 54.190 4.000 ;
    END
  END data_in_a[0]
  PIN data_in_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 -4.000 247.390 4.000 ;
    END
  END data_in_a[10]
  PIN data_in_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 -4.000 266.710 4.000 ;
    END
  END data_in_a[11]
  PIN data_in_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 -4.000 286.030 4.000 ;
    END
  END data_in_a[12]
  PIN data_in_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 -4.000 305.350 4.000 ;
    END
  END data_in_a[13]
  PIN data_in_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 -4.000 324.670 4.000 ;
    END
  END data_in_a[14]
  PIN data_in_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 -4.000 343.990 4.000 ;
    END
  END data_in_a[15]
  PIN data_in_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END data_in_a[1]
  PIN data_in_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END data_in_a[2]
  PIN data_in_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 -4.000 112.150 4.000 ;
    END
  END data_in_a[3]
  PIN data_in_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 -4.000 131.470 4.000 ;
    END
  END data_in_a[4]
  PIN data_in_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 -4.000 150.790 4.000 ;
    END
  END data_in_a[5]
  PIN data_in_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 -4.000 170.110 4.000 ;
    END
  END data_in_a[6]
  PIN data_in_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 -4.000 189.430 4.000 ;
    END
  END data_in_a[7]
  PIN data_in_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 -4.000 208.750 4.000 ;
    END
  END data_in_a[8]
  PIN data_in_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 -4.000 228.070 4.000 ;
    END
  END data_in_a[9]
  PIN driver_io[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 -4.000 15.550 4.000 ;
    END
  END driver_io[0]
  PIN driver_io[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END driver_io[1]
  PIN inverter_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 -4.000 884.950 4.000 ;
    END
  END inverter_select_a
  PIN mem_address_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 -4.000 401.950 4.000 ;
    END
  END mem_address_a[0]
  PIN mem_address_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 -4.000 421.270 4.000 ;
    END
  END mem_address_a[1]
  PIN mem_address_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 -4.000 440.590 4.000 ;
    END
  END mem_address_a[2]
  PIN mem_address_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 -4.000 459.910 4.000 ;
    END
  END mem_address_a[3]
  PIN mem_address_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 -4.000 479.230 4.000 ;
    END
  END mem_address_a[4]
  PIN mem_address_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 -4.000 498.550 4.000 ;
    END
  END mem_address_a[5]
  PIN mem_address_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 -4.000 517.870 4.000 ;
    END
  END mem_address_a[6]
  PIN mem_address_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 -4.000 537.190 4.000 ;
    END
  END mem_address_a[7]
  PIN mem_address_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 -4.000 556.510 4.000 ;
    END
  END mem_address_a[8]
  PIN mem_address_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 -4.000 575.830 4.000 ;
    END
  END mem_address_a[9]
  PIN mem_write_n_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 -4.000 595.150 4.000 ;
    END
  END mem_write_n_a
  PIN output_active_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 -4.000 865.630 4.000 ;
    END
  END output_active_a
  PIN row_col_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 -4.000 846.310 4.000 ;
    END
  END row_col_select_a
  PIN row_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 -4.000 614.470 4.000 ;
    END
  END row_select_a[0]
  PIN row_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 -4.000 633.790 4.000 ;
    END
  END row_select_a[1]
  PIN row_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 -4.000 653.110 4.000 ;
    END
  END row_select_a[2]
  PIN row_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 -4.000 672.430 4.000 ;
    END
  END row_select_a[3]
  PIN row_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 -4.000 691.750 4.000 ;
    END
  END row_select_a[4]
  PIN row_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 -4.000 711.070 4.000 ;
    END
  END row_select_a[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.340 10.640 624.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.340 10.640 724.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.340 10.640 824.340 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 669.340 10.640 674.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.340 10.640 774.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 869.340 10.640 874.340 538.800 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 538.645 ;
      LAYER met1 ;
        RECT 5.520 8.200 894.240 538.800 ;
      LAYER met2 ;
        RECT 15.280 4.280 889.080 538.745 ;
        RECT 15.830 3.670 34.310 4.280 ;
        RECT 35.150 3.670 53.630 4.280 ;
        RECT 54.470 3.670 72.950 4.280 ;
        RECT 73.790 3.670 92.270 4.280 ;
        RECT 93.110 3.670 111.590 4.280 ;
        RECT 112.430 3.670 130.910 4.280 ;
        RECT 131.750 3.670 150.230 4.280 ;
        RECT 151.070 3.670 169.550 4.280 ;
        RECT 170.390 3.670 188.870 4.280 ;
        RECT 189.710 3.670 208.190 4.280 ;
        RECT 209.030 3.670 227.510 4.280 ;
        RECT 228.350 3.670 246.830 4.280 ;
        RECT 247.670 3.670 266.150 4.280 ;
        RECT 266.990 3.670 285.470 4.280 ;
        RECT 286.310 3.670 304.790 4.280 ;
        RECT 305.630 3.670 324.110 4.280 ;
        RECT 324.950 3.670 343.430 4.280 ;
        RECT 344.270 3.670 362.750 4.280 ;
        RECT 363.590 3.670 382.070 4.280 ;
        RECT 382.910 3.670 401.390 4.280 ;
        RECT 402.230 3.670 420.710 4.280 ;
        RECT 421.550 3.670 440.030 4.280 ;
        RECT 440.870 3.670 459.350 4.280 ;
        RECT 460.190 3.670 478.670 4.280 ;
        RECT 479.510 3.670 497.990 4.280 ;
        RECT 498.830 3.670 517.310 4.280 ;
        RECT 518.150 3.670 536.630 4.280 ;
        RECT 537.470 3.670 555.950 4.280 ;
        RECT 556.790 3.670 575.270 4.280 ;
        RECT 576.110 3.670 594.590 4.280 ;
        RECT 595.430 3.670 613.910 4.280 ;
        RECT 614.750 3.670 633.230 4.280 ;
        RECT 634.070 3.670 652.550 4.280 ;
        RECT 653.390 3.670 671.870 4.280 ;
        RECT 672.710 3.670 691.190 4.280 ;
        RECT 692.030 3.670 710.510 4.280 ;
        RECT 711.350 3.670 729.830 4.280 ;
        RECT 730.670 3.670 749.150 4.280 ;
        RECT 749.990 3.670 768.470 4.280 ;
        RECT 769.310 3.670 787.790 4.280 ;
        RECT 788.630 3.670 807.110 4.280 ;
        RECT 807.950 3.670 826.430 4.280 ;
        RECT 827.270 3.670 845.750 4.280 ;
        RECT 846.590 3.670 865.070 4.280 ;
        RECT 865.910 3.670 884.390 4.280 ;
        RECT 885.230 3.670 889.080 4.280 ;
      LAYER met3 ;
        RECT 19.450 10.715 886.355 538.725 ;
      LAYER met4 ;
        RECT 142.895 26.695 168.940 352.745 ;
        RECT 174.740 26.695 218.940 352.745 ;
        RECT 224.740 26.695 268.940 352.745 ;
        RECT 274.740 26.695 318.940 352.745 ;
        RECT 324.740 26.695 368.940 352.745 ;
        RECT 374.740 26.695 418.940 352.745 ;
        RECT 424.740 26.695 468.940 352.745 ;
        RECT 474.740 26.695 518.940 352.745 ;
        RECT 524.740 26.695 568.940 352.745 ;
        RECT 574.740 26.695 618.940 352.745 ;
        RECT 624.740 26.695 668.940 352.745 ;
        RECT 674.740 26.695 718.940 352.745 ;
        RECT 724.740 26.695 768.940 352.745 ;
        RECT 774.740 26.695 807.465 352.745 ;
  END
END driver_core
END LIBRARY

