VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO driver_core
  CLASS BLOCK ;
  FOREIGN driver_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 400.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 -4.000 254.750 4.000 ;
    END
  END clock
  PIN clock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 -4.000 241.870 4.000 ;
    END
  END clock_a
  PIN col_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 -4.000 486.590 4.000 ;
    END
  END col_select_a[0]
  PIN col_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 -4.000 499.470 4.000 ;
    END
  END col_select_a[1]
  PIN col_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 -4.000 512.350 4.000 ;
    END
  END col_select_a[2]
  PIN col_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 -4.000 525.230 4.000 ;
    END
  END col_select_a[3]
  PIN col_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 -4.000 538.110 4.000 ;
    END
  END col_select_a[4]
  PIN col_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 -4.000 550.990 4.000 ;
    END
  END col_select_a[5]
  PIN data_in_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END data_in_a[0]
  PIN data_in_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 -4.000 164.590 4.000 ;
    END
  END data_in_a[10]
  PIN data_in_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 -4.000 177.470 4.000 ;
    END
  END data_in_a[11]
  PIN data_in_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 -4.000 190.350 4.000 ;
    END
  END data_in_a[12]
  PIN data_in_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 -4.000 203.230 4.000 ;
    END
  END data_in_a[13]
  PIN data_in_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 -4.000 216.110 4.000 ;
    END
  END data_in_a[14]
  PIN data_in_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 -4.000 228.990 4.000 ;
    END
  END data_in_a[15]
  PIN data_in_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END data_in_a[1]
  PIN data_in_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 -4.000 61.550 4.000 ;
    END
  END data_in_a[2]
  PIN data_in_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 -4.000 74.430 4.000 ;
    END
  END data_in_a[3]
  PIN data_in_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 -4.000 87.310 4.000 ;
    END
  END data_in_a[4]
  PIN data_in_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 -4.000 100.190 4.000 ;
    END
  END data_in_a[5]
  PIN data_in_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 -4.000 113.070 4.000 ;
    END
  END data_in_a[6]
  PIN data_in_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 -4.000 125.950 4.000 ;
    END
  END data_in_a[7]
  PIN data_in_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 -4.000 138.830 4.000 ;
    END
  END data_in_a[8]
  PIN data_in_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 -4.000 151.710 4.000 ;
    END
  END data_in_a[9]
  PIN driver_io[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 -4.000 10.030 4.000 ;
    END
  END driver_io[0]
  PIN driver_io[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END driver_io[1]
  PIN inverter_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 -4.000 589.630 4.000 ;
    END
  END inverter_select_a
  PIN mem_address_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 -4.000 267.630 4.000 ;
    END
  END mem_address_a[0]
  PIN mem_address_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 -4.000 280.510 4.000 ;
    END
  END mem_address_a[1]
  PIN mem_address_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 -4.000 293.390 4.000 ;
    END
  END mem_address_a[2]
  PIN mem_address_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 -4.000 306.270 4.000 ;
    END
  END mem_address_a[3]
  PIN mem_address_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 -4.000 319.150 4.000 ;
    END
  END mem_address_a[4]
  PIN mem_address_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 -4.000 332.030 4.000 ;
    END
  END mem_address_a[5]
  PIN mem_address_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 -4.000 344.910 4.000 ;
    END
  END mem_address_a[6]
  PIN mem_address_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 -4.000 357.790 4.000 ;
    END
  END mem_address_a[7]
  PIN mem_address_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 -4.000 370.670 4.000 ;
    END
  END mem_address_a[8]
  PIN mem_address_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 -4.000 383.550 4.000 ;
    END
  END mem_address_a[9]
  PIN mem_write_n_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 -4.000 396.430 4.000 ;
    END
  END mem_write_n_a
  PIN output_active_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 -4.000 576.750 4.000 ;
    END
  END output_active_a
  PIN row_col_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 -4.000 563.870 4.000 ;
    END
  END row_col_select_a
  PIN row_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 -4.000 409.310 4.000 ;
    END
  END row_select_a[0]
  PIN row_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 -4.000 422.190 4.000 ;
    END
  END row_select_a[1]
  PIN row_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 -4.000 435.070 4.000 ;
    END
  END row_select_a[2]
  PIN row_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 -4.000 447.950 4.000 ;
    END
  END row_select_a[3]
  PIN row_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 -4.000 460.830 4.000 ;
    END
  END row_select_a[4]
  PIN row_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 -4.000 473.710 4.000 ;
    END
  END row_select_a[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 389.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 387.545 594.510 389.150 ;
        RECT 5.330 382.105 594.510 384.935 ;
        RECT 5.330 376.665 594.510 379.495 ;
        RECT 5.330 371.225 594.510 374.055 ;
        RECT 5.330 365.785 594.510 368.615 ;
        RECT 5.330 360.345 594.510 363.175 ;
        RECT 5.330 354.905 594.510 357.735 ;
        RECT 5.330 349.465 594.510 352.295 ;
        RECT 5.330 344.025 594.510 346.855 ;
        RECT 5.330 338.585 594.510 341.415 ;
        RECT 5.330 333.145 594.510 335.975 ;
        RECT 5.330 327.705 594.510 330.535 ;
        RECT 5.330 322.265 594.510 325.095 ;
        RECT 5.330 316.825 594.510 319.655 ;
        RECT 5.330 311.385 594.510 314.215 ;
        RECT 5.330 305.945 594.510 308.775 ;
        RECT 5.330 300.505 594.510 303.335 ;
        RECT 5.330 295.065 594.510 297.895 ;
        RECT 5.330 289.625 594.510 292.455 ;
        RECT 5.330 284.185 594.510 287.015 ;
        RECT 5.330 278.745 594.510 281.575 ;
        RECT 5.330 273.305 594.510 276.135 ;
        RECT 5.330 267.865 594.510 270.695 ;
        RECT 5.330 262.425 594.510 265.255 ;
        RECT 5.330 256.985 594.510 259.815 ;
        RECT 5.330 251.545 594.510 254.375 ;
        RECT 5.330 246.105 594.510 248.935 ;
        RECT 5.330 240.665 594.510 243.495 ;
        RECT 5.330 235.225 594.510 238.055 ;
        RECT 5.330 229.785 594.510 232.615 ;
        RECT 5.330 224.345 594.510 227.175 ;
        RECT 5.330 218.905 594.510 221.735 ;
        RECT 5.330 213.465 594.510 216.295 ;
        RECT 5.330 208.025 594.510 210.855 ;
        RECT 5.330 202.585 594.510 205.415 ;
        RECT 5.330 197.145 594.510 199.975 ;
        RECT 5.330 191.705 594.510 194.535 ;
        RECT 5.330 186.265 594.510 189.095 ;
        RECT 5.330 180.825 594.510 183.655 ;
        RECT 5.330 175.385 594.510 178.215 ;
        RECT 5.330 169.945 594.510 172.775 ;
        RECT 5.330 164.505 594.510 167.335 ;
        RECT 5.330 159.065 594.510 161.895 ;
        RECT 5.330 153.625 594.510 156.455 ;
        RECT 5.330 148.185 594.510 151.015 ;
        RECT 5.330 142.745 594.510 145.575 ;
        RECT 5.330 137.305 594.510 140.135 ;
        RECT 5.330 131.865 594.510 134.695 ;
        RECT 5.330 126.425 594.510 129.255 ;
        RECT 5.330 120.985 594.510 123.815 ;
        RECT 5.330 115.545 594.510 118.375 ;
        RECT 5.330 110.105 594.510 112.935 ;
        RECT 5.330 104.665 594.510 107.495 ;
        RECT 5.330 99.225 594.510 102.055 ;
        RECT 5.330 93.785 594.510 96.615 ;
        RECT 5.330 88.345 594.510 91.175 ;
        RECT 5.330 82.905 594.510 85.735 ;
        RECT 5.330 77.465 594.510 80.295 ;
        RECT 5.330 72.025 594.510 74.855 ;
        RECT 5.330 66.585 594.510 69.415 ;
        RECT 5.330 61.145 594.510 63.975 ;
        RECT 5.330 55.705 594.510 58.535 ;
        RECT 5.330 50.265 594.510 53.095 ;
        RECT 5.330 44.825 594.510 47.655 ;
        RECT 5.330 39.385 594.510 42.215 ;
        RECT 5.330 33.945 594.510 36.775 ;
        RECT 5.330 28.505 594.510 31.335 ;
        RECT 5.330 23.065 594.510 25.895 ;
        RECT 5.330 17.625 594.510 20.455 ;
        RECT 5.330 12.185 594.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 594.320 389.045 ;
      LAYER met1 ;
        RECT 5.520 6.160 594.320 389.200 ;
      LAYER met2 ;
        RECT 7.920 4.280 591.000 389.145 ;
        RECT 7.920 3.670 9.470 4.280 ;
        RECT 10.310 3.670 22.350 4.280 ;
        RECT 23.190 3.670 35.230 4.280 ;
        RECT 36.070 3.670 48.110 4.280 ;
        RECT 48.950 3.670 60.990 4.280 ;
        RECT 61.830 3.670 73.870 4.280 ;
        RECT 74.710 3.670 86.750 4.280 ;
        RECT 87.590 3.670 99.630 4.280 ;
        RECT 100.470 3.670 112.510 4.280 ;
        RECT 113.350 3.670 125.390 4.280 ;
        RECT 126.230 3.670 138.270 4.280 ;
        RECT 139.110 3.670 151.150 4.280 ;
        RECT 151.990 3.670 164.030 4.280 ;
        RECT 164.870 3.670 176.910 4.280 ;
        RECT 177.750 3.670 189.790 4.280 ;
        RECT 190.630 3.670 202.670 4.280 ;
        RECT 203.510 3.670 215.550 4.280 ;
        RECT 216.390 3.670 228.430 4.280 ;
        RECT 229.270 3.670 241.310 4.280 ;
        RECT 242.150 3.670 254.190 4.280 ;
        RECT 255.030 3.670 267.070 4.280 ;
        RECT 267.910 3.670 279.950 4.280 ;
        RECT 280.790 3.670 292.830 4.280 ;
        RECT 293.670 3.670 305.710 4.280 ;
        RECT 306.550 3.670 318.590 4.280 ;
        RECT 319.430 3.670 331.470 4.280 ;
        RECT 332.310 3.670 344.350 4.280 ;
        RECT 345.190 3.670 357.230 4.280 ;
        RECT 358.070 3.670 370.110 4.280 ;
        RECT 370.950 3.670 382.990 4.280 ;
        RECT 383.830 3.670 395.870 4.280 ;
        RECT 396.710 3.670 408.750 4.280 ;
        RECT 409.590 3.670 421.630 4.280 ;
        RECT 422.470 3.670 434.510 4.280 ;
        RECT 435.350 3.670 447.390 4.280 ;
        RECT 448.230 3.670 460.270 4.280 ;
        RECT 461.110 3.670 473.150 4.280 ;
        RECT 473.990 3.670 486.030 4.280 ;
        RECT 486.870 3.670 498.910 4.280 ;
        RECT 499.750 3.670 511.790 4.280 ;
        RECT 512.630 3.670 524.670 4.280 ;
        RECT 525.510 3.670 537.550 4.280 ;
        RECT 538.390 3.670 550.430 4.280 ;
        RECT 551.270 3.670 563.310 4.280 ;
        RECT 564.150 3.670 576.190 4.280 ;
        RECT 577.030 3.670 589.070 4.280 ;
        RECT 589.910 3.670 591.000 4.280 ;
      LAYER met3 ;
        RECT 19.450 7.655 590.575 389.125 ;
      LAYER met4 ;
        RECT 74.815 15.815 118.940 364.985 ;
        RECT 124.740 15.815 168.940 364.985 ;
        RECT 174.740 15.815 218.940 364.985 ;
        RECT 224.740 15.815 268.940 364.985 ;
        RECT 274.740 15.815 318.940 364.985 ;
        RECT 324.740 15.815 368.940 364.985 ;
        RECT 374.740 15.815 418.940 364.985 ;
        RECT 424.740 15.815 468.940 364.985 ;
        RECT 474.740 15.815 513.065 364.985 ;
  END
END driver_core
END LIBRARY

