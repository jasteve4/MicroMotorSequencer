magic
tech sky130B
magscale 1 2
timestamp 1661812818
<< metal1 >>
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 202782 700992 202788 701004
rect 137888 700964 202788 700992
rect 137888 700952 137894 700964
rect 202782 700952 202788 700964
rect 202840 700952 202846 701004
rect 397454 700952 397460 701004
rect 397512 700992 397518 701004
rect 462314 700992 462320 701004
rect 397512 700964 462320 700992
rect 397512 700952 397518 700964
rect 462314 700952 462320 700964
rect 462372 700952 462378 701004
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 16482 700516 16488 700528
rect 8168 700488 16488 700516
rect 8168 700476 8174 700488
rect 16482 700476 16488 700488
rect 16540 700516 16546 700528
rect 72970 700516 72976 700528
rect 16540 700488 72976 700516
rect 16540 700476 16546 700488
rect 72970 700476 72976 700488
rect 73028 700476 73034 700528
rect 295242 700476 295248 700528
rect 295300 700516 295306 700528
rect 397454 700516 397460 700528
rect 295300 700488 397460 700516
rect 295300 700476 295306 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 20622 700408 20628 700460
rect 20680 700448 20686 700460
rect 89162 700448 89168 700460
rect 20680 700420 89168 700448
rect 20680 700408 20686 700420
rect 89162 700408 89168 700420
rect 89220 700408 89226 700460
rect 300578 700408 300584 700460
rect 300636 700448 300642 700460
rect 413646 700448 413652 700460
rect 300636 700420 413652 700448
rect 300636 700408 300642 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 20438 700340 20444 700392
rect 20496 700380 20502 700392
rect 154114 700380 154120 700392
rect 20496 700352 154120 700380
rect 20496 700340 20502 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 300670 700340 300676 700392
rect 300728 700380 300734 700392
rect 478506 700380 478512 700392
rect 300728 700352 478512 700380
rect 300728 700340 300734 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 20346 700272 20352 700324
rect 20404 700312 20410 700324
rect 218974 700312 218980 700324
rect 20404 700284 218980 700312
rect 20404 700272 20410 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 300762 700272 300768 700324
rect 300820 700312 300826 700324
rect 543458 700312 543464 700324
rect 300820 700284 543464 700312
rect 300820 700272 300826 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 20530 699660 20536 699712
rect 20588 699700 20594 699712
rect 24302 699700 24308 699712
rect 20588 699672 24308 699700
rect 20588 699660 20594 699672
rect 24302 699660 24308 699672
rect 24360 699660 24366 699712
rect 527174 697552 527180 697604
rect 527232 697592 527238 697604
rect 574094 697592 574100 697604
rect 527232 697564 574100 697592
rect 527232 697552 527238 697564
rect 574094 697552 574100 697564
rect 574152 697552 574158 697604
rect 574094 696940 574100 696992
rect 574152 696980 574158 696992
rect 580166 696980 580172 696992
rect 574152 696952 580172 696980
rect 574152 696940 574158 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 671032 3424 671084
rect 3476 671072 3482 671084
rect 7650 671072 7656 671084
rect 3476 671044 7656 671072
rect 3476 671032 3482 671044
rect 7650 671032 7656 671044
rect 7708 671032 7714 671084
rect 2866 618876 2872 618928
rect 2924 618916 2930 618928
rect 4982 618916 4988 618928
rect 2924 618888 4988 618916
rect 2924 618876 2930 618888
rect 4982 618876 4988 618888
rect 5040 618876 5046 618928
rect 300578 588616 300584 588668
rect 300636 588656 300642 588668
rect 304166 588656 304172 588668
rect 300636 588628 304172 588656
rect 300636 588616 300642 588628
rect 304166 588616 304172 588628
rect 304224 588616 304230 588668
rect 300670 586508 300676 586560
rect 300728 586548 300734 586560
rect 310330 586548 310336 586560
rect 300728 586520 310336 586548
rect 300728 586508 300734 586520
rect 310330 586508 310336 586520
rect 310388 586508 310394 586560
rect 20438 586440 20444 586492
rect 20496 586480 20502 586492
rect 24210 586480 24216 586492
rect 20496 586452 24216 586480
rect 20496 586440 20502 586452
rect 24210 586440 24216 586452
rect 24268 586440 24274 586492
rect 129182 586440 129188 586492
rect 129240 586480 129246 586492
rect 134334 586480 134340 586492
rect 129240 586452 134340 586480
rect 129240 586440 129246 586452
rect 134334 586440 134340 586452
rect 134392 586440 134398 586492
rect 198642 586440 198648 586492
rect 198700 586480 198706 586492
rect 292574 586480 292580 586492
rect 198700 586452 292580 586480
rect 198700 586440 198706 586452
rect 292574 586440 292580 586452
rect 292632 586440 292638 586492
rect 408862 586440 408868 586492
rect 408920 586480 408926 586492
rect 414658 586480 414664 586492
rect 408920 586452 414664 586480
rect 408920 586440 408926 586452
rect 414658 586440 414664 586452
rect 414716 586440 414722 586492
rect 20346 586372 20352 586424
rect 20404 586412 20410 586424
rect 30006 586412 30012 586424
rect 20404 586384 30012 586412
rect 20404 586372 20410 586384
rect 30006 586372 30012 586384
rect 30064 586372 30070 586424
rect 559558 586168 559564 586220
rect 559616 586208 559622 586220
rect 569954 586208 569960 586220
rect 559616 586180 569960 586208
rect 559616 586168 559622 586180
rect 569954 586168 569960 586180
rect 570012 586168 570018 586220
rect 22002 586100 22008 586152
rect 22060 586140 22066 586152
rect 47394 586140 47400 586152
rect 22060 586112 47400 586140
rect 22060 586100 22066 586112
rect 47394 586100 47400 586112
rect 47452 586100 47458 586152
rect 300486 586100 300492 586152
rect 300544 586140 300550 586152
rect 316126 586140 316132 586152
rect 300544 586112 316132 586140
rect 300544 586100 300550 586112
rect 316126 586100 316132 586112
rect 316184 586100 316190 586152
rect 553762 586100 553768 586152
rect 553820 586140 553826 586152
rect 572714 586140 572720 586152
rect 553820 586112 572720 586140
rect 553820 586100 553826 586112
rect 572714 586100 572720 586112
rect 572772 586100 572778 586152
rect 20438 586032 20444 586084
rect 20496 586072 20502 586084
rect 53190 586072 53196 586084
rect 20496 586044 53196 586072
rect 20496 586032 20502 586044
rect 53190 586032 53196 586044
rect 53248 586032 53254 586084
rect 279878 586032 279884 586084
rect 279936 586072 279942 586084
rect 289998 586072 290004 586084
rect 279936 586044 290004 586072
rect 279936 586032 279942 586044
rect 289998 586032 290004 586044
rect 290056 586032 290062 586084
rect 300670 586032 300676 586084
rect 300728 586072 300734 586084
rect 321922 586072 321928 586084
rect 300728 586044 321928 586072
rect 300728 586032 300734 586044
rect 321922 586032 321928 586044
rect 321980 586032 321986 586084
rect 547966 586032 547972 586084
rect 548024 586072 548030 586084
rect 570138 586072 570144 586084
rect 548024 586044 570144 586072
rect 548024 586032 548030 586044
rect 570138 586032 570144 586044
rect 570196 586032 570202 586084
rect 17862 585964 17868 586016
rect 17920 586004 17926 586016
rect 58986 586004 58992 586016
rect 17920 585976 58992 586004
rect 17920 585964 17926 585976
rect 58986 585964 58992 585976
rect 59044 585964 59050 586016
rect 268286 585964 268292 586016
rect 268344 586004 268350 586016
rect 289906 586004 289912 586016
rect 268344 585976 289912 586004
rect 268344 585964 268350 585976
rect 289906 585964 289912 585976
rect 289964 585964 289970 586016
rect 302142 585964 302148 586016
rect 302200 586004 302206 586016
rect 327718 586004 327724 586016
rect 302200 585976 327724 586004
rect 302200 585964 302206 585976
rect 327718 585964 327724 585976
rect 327776 585964 327782 586016
rect 542170 585964 542176 586016
rect 542228 586004 542234 586016
rect 570046 586004 570052 586016
rect 542228 585976 570052 586004
rect 542228 585964 542234 585976
rect 570046 585964 570052 585976
rect 570104 585964 570110 586016
rect 20346 585896 20352 585948
rect 20404 585936 20410 585948
rect 35894 585936 35900 585948
rect 20404 585908 35900 585936
rect 20404 585896 20410 585908
rect 35894 585896 35900 585908
rect 35952 585896 35958 585948
rect 37918 585896 37924 585948
rect 37976 585936 37982 585948
rect 105354 585936 105360 585948
rect 37976 585908 105360 585936
rect 37976 585896 37982 585908
rect 105354 585896 105360 585908
rect 105412 585896 105418 585948
rect 262122 585896 262128 585948
rect 262180 585936 262186 585948
rect 289814 585936 289820 585948
rect 262180 585908 289820 585936
rect 262180 585896 262186 585908
rect 289814 585896 289820 585908
rect 289872 585896 289878 585948
rect 300578 585896 300584 585948
rect 300636 585936 300642 585948
rect 333514 585936 333520 585948
rect 300636 585908 333520 585936
rect 300636 585896 300642 585908
rect 333514 585896 333520 585908
rect 333572 585896 333578 585948
rect 536374 585896 536380 585948
rect 536432 585936 536438 585948
rect 568574 585936 568580 585948
rect 536432 585908 568580 585936
rect 536432 585896 536438 585908
rect 568574 585896 568580 585908
rect 568632 585896 568638 585948
rect 31018 585828 31024 585880
rect 31076 585868 31082 585880
rect 99558 585868 99564 585880
rect 31076 585840 99564 585868
rect 31076 585828 31082 585840
rect 99558 585828 99564 585840
rect 99616 585828 99622 585880
rect 256602 585828 256608 585880
rect 256660 585868 256666 585880
rect 288434 585868 288440 585880
rect 256660 585840 288440 585868
rect 256660 585828 256666 585840
rect 288434 585828 288440 585840
rect 288492 585828 288498 585880
rect 297818 585828 297824 585880
rect 297876 585868 297882 585880
rect 339310 585868 339316 585880
rect 297876 585840 339316 585868
rect 297876 585828 297882 585840
rect 339310 585828 339316 585840
rect 339368 585828 339374 585880
rect 524782 585828 524788 585880
rect 524840 585868 524846 585880
rect 569310 585868 569316 585880
rect 524840 585840 569316 585868
rect 524840 585828 524846 585840
rect 569310 585828 569316 585840
rect 569368 585828 569374 585880
rect 20254 585760 20260 585812
rect 20312 585800 20318 585812
rect 41598 585800 41604 585812
rect 20312 585772 41604 585800
rect 20312 585760 20318 585772
rect 41598 585760 41604 585772
rect 41656 585760 41662 585812
rect 43438 585760 43444 585812
rect 43496 585800 43502 585812
rect 116946 585800 116952 585812
rect 43496 585772 116952 585800
rect 43496 585760 43502 585772
rect 116946 585760 116952 585772
rect 117004 585760 117010 585812
rect 250898 585760 250904 585812
rect 250956 585800 250962 585812
rect 288618 585800 288624 585812
rect 250956 585772 288624 585800
rect 250956 585760 250962 585772
rect 288618 585760 288624 585772
rect 288676 585760 288682 585812
rect 299382 585760 299388 585812
rect 299440 585800 299446 585812
rect 345106 585800 345112 585812
rect 299440 585772 345112 585800
rect 299440 585760 299446 585772
rect 345106 585760 345112 585772
rect 345164 585760 345170 585812
rect 507394 585760 507400 585812
rect 507452 585800 507458 585812
rect 568666 585800 568672 585812
rect 507452 585772 568672 585800
rect 507452 585760 507458 585772
rect 568666 585760 568672 585772
rect 568724 585760 568730 585812
rect 17678 583380 17684 583432
rect 17736 583420 17742 583432
rect 76374 583420 76380 583432
rect 17736 583392 76380 583420
rect 17736 583380 17742 583392
rect 76374 583380 76380 583392
rect 76432 583380 76438 583432
rect 233142 583380 233148 583432
rect 233200 583420 233206 583432
rect 291286 583420 291292 583432
rect 233200 583392 291292 583420
rect 233200 583380 233206 583392
rect 291286 583380 291292 583392
rect 291344 583380 291350 583432
rect 17770 583312 17776 583364
rect 17828 583352 17834 583364
rect 87966 583352 87972 583364
rect 17828 583324 87972 583352
rect 17828 583312 17834 583324
rect 87966 583312 87972 583324
rect 88024 583312 88030 583364
rect 221918 583312 221924 583364
rect 221976 583352 221982 583364
rect 292758 583352 292764 583364
rect 221976 583324 292764 583352
rect 221976 583312 221982 583324
rect 292758 583312 292764 583324
rect 292816 583312 292822 583364
rect 513190 583312 513196 583364
rect 513248 583352 513254 583364
rect 571518 583352 571524 583364
rect 513248 583324 571524 583352
rect 513248 583312 513254 583324
rect 571518 583312 571524 583324
rect 571576 583312 571582 583364
rect 19150 583244 19156 583296
rect 19208 583284 19214 583296
rect 93854 583284 93860 583296
rect 19208 583256 93860 583284
rect 19208 583244 19214 583256
rect 93854 583244 93860 583256
rect 93912 583244 93918 583296
rect 216122 583244 216128 583296
rect 216180 583284 216186 583296
rect 291194 583284 291200 583296
rect 216180 583256 291200 583284
rect 216180 583244 216186 583256
rect 291194 583244 291200 583256
rect 291252 583244 291258 583296
rect 297726 583244 297732 583296
rect 297784 583284 297790 583296
rect 356698 583284 356704 583296
rect 297784 583256 356704 583284
rect 297784 583244 297790 583256
rect 356698 583244 356704 583256
rect 356756 583244 356762 583296
rect 501598 583244 501604 583296
rect 501656 583284 501662 583296
rect 571426 583284 571432 583296
rect 501656 583256 571432 583284
rect 501656 583244 501662 583256
rect 571426 583244 571432 583256
rect 571484 583244 571490 583296
rect 15010 583176 15016 583228
rect 15068 583216 15074 583228
rect 111150 583216 111156 583228
rect 15068 583188 111156 583216
rect 15068 583176 15074 583188
rect 111150 583176 111156 583188
rect 111208 583176 111214 583228
rect 210326 583176 210332 583228
rect 210384 583216 210390 583228
rect 292574 583216 292580 583228
rect 210384 583188 292580 583216
rect 210384 583176 210390 583188
rect 292574 583176 292580 583188
rect 292632 583176 292638 583228
rect 298830 583176 298836 583228
rect 298888 583216 298894 583228
rect 368290 583216 368296 583228
rect 298888 583188 368296 583216
rect 298888 583176 298894 583188
rect 368290 583176 368296 583188
rect 368348 583176 368354 583228
rect 490006 583176 490012 583228
rect 490064 583216 490070 583228
rect 574186 583216 574192 583228
rect 490064 583188 574192 583216
rect 490064 583176 490070 583188
rect 574186 583176 574192 583188
rect 574244 583176 574250 583228
rect 19058 583108 19064 583160
rect 19116 583148 19122 583160
rect 122834 583148 122840 583160
rect 19116 583120 122840 583148
rect 19116 583108 19122 583120
rect 122834 583108 122840 583120
rect 122892 583108 122898 583160
rect 204162 583108 204168 583160
rect 204220 583148 204226 583160
rect 291378 583148 291384 583160
rect 204220 583120 291384 583148
rect 204220 583108 204226 583120
rect 291378 583108 291384 583120
rect 291436 583108 291442 583160
rect 299198 583108 299204 583160
rect 299256 583148 299262 583160
rect 374086 583148 374092 583160
rect 299256 583120 374092 583148
rect 299256 583108 299262 583120
rect 374086 583108 374092 583120
rect 374144 583108 374150 583160
rect 484210 583108 484216 583160
rect 484268 583148 484274 583160
rect 571610 583148 571616 583160
rect 484268 583120 571616 583148
rect 484268 583108 484274 583120
rect 571610 583108 571616 583120
rect 571668 583108 571674 583160
rect 15102 583040 15108 583092
rect 15160 583080 15166 583092
rect 140130 583080 140136 583092
rect 15160 583052 140136 583080
rect 15160 583040 15166 583052
rect 140130 583040 140136 583052
rect 140188 583040 140194 583092
rect 192938 583040 192944 583092
rect 192996 583080 193002 583092
rect 293954 583080 293960 583092
rect 192996 583052 293960 583080
rect 192996 583040 193002 583052
rect 293954 583040 293960 583052
rect 294012 583040 294018 583092
rect 297910 583040 297916 583092
rect 297968 583080 297974 583092
rect 379882 583080 379888 583092
rect 297968 583052 379888 583080
rect 297968 583040 297974 583052
rect 379882 583040 379888 583052
rect 379940 583040 379946 583092
rect 472618 583040 472624 583092
rect 472676 583080 472682 583092
rect 572806 583080 572812 583092
rect 472676 583052 572812 583080
rect 472676 583040 472682 583052
rect 572806 583040 572812 583052
rect 572864 583040 572870 583092
rect 16390 582972 16396 583024
rect 16448 583012 16454 583024
rect 151814 583012 151820 583024
rect 16448 582984 151820 583012
rect 16448 582972 16454 582984
rect 151814 582972 151820 582984
rect 151872 582972 151878 583024
rect 175182 582972 175188 583024
rect 175240 583012 175246 583024
rect 291838 583012 291844 583024
rect 175240 582984 291844 583012
rect 175240 582972 175246 582984
rect 291838 582972 291844 582984
rect 291896 582972 291902 583024
rect 296622 582972 296628 583024
rect 296680 583012 296686 583024
rect 391474 583012 391480 583024
rect 296680 582984 391480 583012
rect 296680 582972 296686 582984
rect 391474 582972 391480 582984
rect 391532 582972 391538 583024
rect 455230 582972 455236 583024
rect 455288 583012 455294 583024
rect 571334 583012 571340 583024
rect 455288 582984 571340 583012
rect 455288 582972 455294 582984
rect 571334 582972 571340 582984
rect 571392 582972 571398 583024
rect 296530 580524 296536 580576
rect 296588 580564 296594 580576
rect 397270 580564 397276 580576
rect 296588 580536 397276 580564
rect 296588 580524 296594 580536
rect 397270 580524 397276 580536
rect 397328 580524 397334 580576
rect 300394 580456 300400 580508
rect 300452 580496 300458 580508
rect 403066 580496 403072 580508
rect 300452 580468 403072 580496
rect 300452 580456 300458 580468
rect 403066 580456 403072 580468
rect 403124 580456 403130 580508
rect 181346 580388 181352 580440
rect 181404 580428 181410 580440
rect 293218 580428 293224 580440
rect 181404 580400 293224 580428
rect 181404 580388 181410 580400
rect 293218 580388 293224 580400
rect 293276 580388 293282 580440
rect 296438 580388 296444 580440
rect 296496 580428 296502 580440
rect 420454 580428 420460 580440
rect 296496 580400 420460 580428
rect 296496 580388 296502 580400
rect 420454 580388 420460 580400
rect 420512 580388 420518 580440
rect 158162 580320 158168 580372
rect 158220 580360 158226 580372
rect 288526 580360 288532 580372
rect 158220 580332 288532 580360
rect 158220 580320 158226 580332
rect 288526 580320 288532 580332
rect 288584 580320 288590 580372
rect 298002 580320 298008 580372
rect 298060 580360 298066 580372
rect 426250 580360 426256 580372
rect 298060 580332 426256 580360
rect 298060 580320 298066 580332
rect 426250 580320 426256 580332
rect 426308 580320 426314 580372
rect 14918 580252 14924 580304
rect 14976 580292 14982 580304
rect 145926 580292 145932 580304
rect 14976 580264 145932 580292
rect 14976 580252 14982 580264
rect 145926 580252 145932 580264
rect 145984 580252 145990 580304
rect 163958 580252 163964 580304
rect 164016 580292 164022 580304
rect 294046 580292 294052 580304
rect 164016 580264 294052 580292
rect 164016 580252 164022 580264
rect 294046 580252 294052 580264
rect 294104 580252 294110 580304
rect 299106 580252 299112 580304
rect 299164 580292 299170 580304
rect 432046 580292 432052 580304
rect 299164 580264 432052 580292
rect 299164 580252 299170 580264
rect 432046 580252 432052 580264
rect 432104 580252 432110 580304
rect 449434 580252 449440 580304
rect 449492 580292 449498 580304
rect 572898 580292 572904 580304
rect 449492 580264 572904 580292
rect 449492 580252 449498 580264
rect 572898 580252 572904 580264
rect 572956 580252 572962 580304
rect 273254 572160 273260 572212
rect 273312 572200 273318 572212
rect 294598 572200 294604 572212
rect 273312 572172 294604 572200
rect 273312 572160 273318 572172
rect 294598 572160 294604 572172
rect 294656 572160 294662 572212
rect 529934 572160 529940 572212
rect 529992 572200 529998 572212
rect 570230 572200 570236 572212
rect 529992 572172 570236 572200
rect 529992 572160 529998 572172
rect 570230 572160 570236 572172
rect 570288 572160 570294 572212
rect 18598 572092 18604 572144
rect 18656 572132 18662 572144
rect 31018 572132 31024 572144
rect 18656 572104 31024 572132
rect 18656 572092 18662 572104
rect 31018 572092 31024 572104
rect 31076 572092 31082 572144
rect 244274 572092 244280 572144
rect 244332 572132 244338 572144
rect 290090 572132 290096 572144
rect 244332 572104 290096 572132
rect 244332 572092 244338 572104
rect 290090 572092 290096 572104
rect 290148 572092 290154 572144
rect 495434 572092 495440 572144
rect 495492 572132 495498 572144
rect 571702 572132 571708 572144
rect 495492 572104 571708 572132
rect 495492 572092 495498 572104
rect 571702 572092 571708 572104
rect 571760 572092 571766 572144
rect 17586 572024 17592 572076
rect 17644 572064 17650 572076
rect 37918 572064 37924 572076
rect 17644 572036 37924 572064
rect 17644 572024 17650 572036
rect 37918 572024 37924 572036
rect 37976 572024 37982 572076
rect 186314 572024 186320 572076
rect 186372 572064 186378 572076
rect 290182 572064 290188 572076
rect 186372 572036 290188 572064
rect 186372 572024 186378 572036
rect 290182 572024 290188 572036
rect 290240 572024 290246 572076
rect 460934 572024 460940 572076
rect 460992 572064 460998 572076
rect 572990 572064 572996 572076
rect 460992 572036 572996 572064
rect 460992 572024 460998 572036
rect 572990 572024 572996 572036
rect 573048 572024 573054 572076
rect 18690 571956 18696 572008
rect 18748 571996 18754 572008
rect 43438 571996 43444 572008
rect 18748 571968 43444 571996
rect 18748 571956 18754 571968
rect 43438 571956 43444 571968
rect 43496 571956 43502 572008
rect 168374 571956 168380 572008
rect 168432 571996 168438 572008
rect 293310 571996 293316 572008
rect 168432 571968 293316 571996
rect 168432 571956 168438 571968
rect 293310 571956 293316 571968
rect 293368 571956 293374 572008
rect 442994 571956 443000 572008
rect 443052 571996 443058 572008
rect 575566 571996 575572 572008
rect 443052 571968 575572 571996
rect 443052 571956 443058 571968
rect 575566 571956 575572 571968
rect 575624 571956 575630 572008
rect 569218 485052 569224 485104
rect 569276 485092 569282 485104
rect 580534 485092 580540 485104
rect 569276 485064 580540 485092
rect 569276 485052 569282 485064
rect 580534 485052 580540 485064
rect 580592 485092 580598 485104
rect 580902 485092 580908 485104
rect 580592 485064 580908 485092
rect 580592 485052 580598 485064
rect 580902 485052 580908 485064
rect 580960 485052 580966 485104
rect 19058 463360 19064 463412
rect 19116 463400 19122 463412
rect 23382 463400 23388 463412
rect 19116 463372 23388 463400
rect 19116 463360 19122 463372
rect 23382 463360 23388 463372
rect 23440 463360 23446 463412
rect 291838 462544 291844 462596
rect 291896 462584 291902 462596
rect 292942 462584 292948 462596
rect 291896 462556 292948 462584
rect 291896 462544 291902 462556
rect 292942 462544 292948 462556
rect 293000 462544 293006 462596
rect 2774 462408 2780 462460
rect 2832 462448 2838 462460
rect 4798 462448 4804 462460
rect 2832 462420 4804 462448
rect 2832 462408 2838 462420
rect 4798 462408 4804 462420
rect 4856 462408 4862 462460
rect 24854 462408 24860 462460
rect 24912 462448 24918 462460
rect 140130 462448 140136 462460
rect 24912 462420 140136 462448
rect 24912 462408 24918 462420
rect 140130 462408 140136 462420
rect 140188 462408 140194 462460
rect 296622 462408 296628 462460
rect 296680 462448 296686 462460
rect 391198 462448 391204 462460
rect 296680 462420 391204 462448
rect 296680 462408 296686 462420
rect 391198 462408 391204 462420
rect 391256 462408 391262 462460
rect 438210 462408 438216 462460
rect 438268 462448 438274 462460
rect 568758 462448 568764 462460
rect 438268 462420 568764 462448
rect 438268 462408 438274 462420
rect 568758 462408 568764 462420
rect 568816 462448 568822 462460
rect 575474 462448 575480 462460
rect 568816 462420 575480 462448
rect 568816 462408 568822 462420
rect 575474 462408 575480 462420
rect 575532 462408 575538 462460
rect 151906 462380 151912 462392
rect 26206 462352 151912 462380
rect 14826 462272 14832 462324
rect 14884 462312 14890 462324
rect 15010 462312 15016 462324
rect 14884 462284 15016 462312
rect 14884 462272 14890 462284
rect 15010 462272 15016 462284
rect 15068 462272 15074 462324
rect 16390 462272 16396 462324
rect 16448 462312 16454 462324
rect 26206 462312 26234 462352
rect 151906 462340 151912 462352
rect 151964 462340 151970 462392
rect 292574 462340 292580 462392
rect 292632 462380 292638 462392
rect 293218 462380 293224 462392
rect 292632 462352 293224 462380
rect 292632 462340 292638 462352
rect 293218 462340 293224 462352
rect 293276 462380 293282 462392
rect 296714 462380 296720 462392
rect 293276 462352 296720 462380
rect 293276 462340 293282 462352
rect 296714 462340 296720 462352
rect 296772 462340 296778 462392
rect 300118 462340 300124 462392
rect 300176 462380 300182 462392
rect 402882 462380 402888 462392
rect 300176 462352 402888 462380
rect 300176 462340 300182 462352
rect 402882 462340 402888 462352
rect 402940 462340 402946 462392
rect 443730 462340 443736 462392
rect 443788 462380 443794 462392
rect 575566 462380 575572 462392
rect 443788 462352 575572 462380
rect 443788 462340 443794 462352
rect 575566 462340 575572 462352
rect 575624 462340 575630 462392
rect 16448 462284 26234 462312
rect 16448 462272 16454 462284
rect 288250 462272 288256 462324
rect 288308 462312 288314 462324
rect 288526 462312 288532 462324
rect 288308 462284 288532 462312
rect 288308 462272 288314 462284
rect 288526 462272 288532 462284
rect 288584 462272 288590 462324
rect 291470 462272 291476 462324
rect 291528 462312 291534 462324
rect 294046 462312 294052 462324
rect 291528 462284 294052 462312
rect 291528 462272 291534 462284
rect 294046 462272 294052 462284
rect 294104 462272 294110 462324
rect 297818 462272 297824 462324
rect 297876 462312 297882 462324
rect 300210 462312 300216 462324
rect 297876 462284 300216 462312
rect 297876 462272 297882 462284
rect 300210 462272 300216 462284
rect 300268 462272 300274 462324
rect 300762 462272 300768 462324
rect 300820 462312 300826 462324
rect 304166 462312 304172 462324
rect 300820 462284 304172 462312
rect 300820 462272 300826 462284
rect 304166 462272 304172 462284
rect 304224 462272 304230 462324
rect 570322 462272 570328 462324
rect 570380 462312 570386 462324
rect 571610 462312 571616 462324
rect 570380 462284 571616 462312
rect 570380 462272 570386 462284
rect 571610 462272 571616 462284
rect 571668 462272 571674 462324
rect 20530 462204 20536 462256
rect 20588 462244 20594 462256
rect 24210 462244 24216 462256
rect 20588 462216 24216 462244
rect 20588 462204 20594 462216
rect 24210 462204 24216 462216
rect 24268 462204 24274 462256
rect 297726 462204 297732 462256
rect 297784 462244 297790 462256
rect 298738 462244 298744 462256
rect 297784 462216 298744 462244
rect 297784 462204 297790 462216
rect 298738 462204 298744 462216
rect 298796 462204 298802 462256
rect 300670 462204 300676 462256
rect 300728 462244 300734 462256
rect 302142 462244 302148 462256
rect 300728 462216 302148 462244
rect 300728 462204 300734 462216
rect 302142 462204 302148 462216
rect 302200 462204 302206 462256
rect 300302 461864 300308 461916
rect 300360 461904 300366 461916
rect 300578 461904 300584 461916
rect 300360 461876 300584 461904
rect 300360 461864 300366 461876
rect 300578 461864 300584 461876
rect 300636 461864 300642 461916
rect 15102 461592 15108 461644
rect 15160 461632 15166 461644
rect 17402 461632 17408 461644
rect 15160 461604 17408 461632
rect 15160 461592 15166 461604
rect 17402 461592 17408 461604
rect 17460 461632 17466 461644
rect 24854 461632 24860 461644
rect 17460 461604 24860 461632
rect 17460 461592 17466 461604
rect 24854 461592 24860 461604
rect 24912 461592 24918 461644
rect 291286 461320 291292 461372
rect 291344 461360 291350 461372
rect 291562 461360 291568 461372
rect 291344 461332 291568 461360
rect 291344 461320 291350 461332
rect 291562 461320 291568 461332
rect 291620 461320 291626 461372
rect 455322 461320 455328 461372
rect 455380 461360 455386 461372
rect 567102 461360 567108 461372
rect 455380 461332 567108 461360
rect 455380 461320 455386 461332
rect 567102 461320 567108 461332
rect 567160 461360 567166 461372
rect 571334 461360 571340 461372
rect 567160 461332 571340 461360
rect 567160 461320 567166 461332
rect 571334 461320 571340 461332
rect 571392 461320 571398 461372
rect 158162 461252 158168 461304
rect 158220 461292 158226 461304
rect 288250 461292 288256 461304
rect 158220 461264 288256 461292
rect 158220 461252 158226 461264
rect 288250 461252 288256 461264
rect 288308 461252 288314 461304
rect 233326 461184 233332 461236
rect 233384 461224 233390 461236
rect 291304 461224 291332 461320
rect 513282 461252 513288 461304
rect 513340 461292 513346 461304
rect 571518 461292 571524 461304
rect 513340 461264 571524 461292
rect 513340 461252 513346 461264
rect 571518 461252 571524 461264
rect 571576 461252 571582 461304
rect 233384 461196 291332 461224
rect 233384 461184 233390 461196
rect 300210 461184 300216 461236
rect 300268 461224 300274 461236
rect 336734 461224 336740 461236
rect 300268 461196 336740 461224
rect 300268 461184 300274 461196
rect 336734 461184 336740 461196
rect 336792 461184 336798 461236
rect 507762 461184 507768 461236
rect 507820 461224 507826 461236
rect 567746 461224 567752 461236
rect 507820 461196 567752 461224
rect 507820 461184 507826 461196
rect 567746 461184 567752 461196
rect 567804 461224 567810 461236
rect 568666 461224 568672 461236
rect 567804 461196 568672 461224
rect 567804 461184 567810 461196
rect 568666 461184 568672 461196
rect 568724 461184 568730 461236
rect 181346 461116 181352 461168
rect 181404 461156 181410 461168
rect 292574 461156 292580 461168
rect 181404 461128 292580 461156
rect 181404 461116 181410 461128
rect 292574 461116 292580 461128
rect 292632 461116 292638 461168
rect 299290 461116 299296 461168
rect 299348 461156 299354 461168
rect 302050 461156 302056 461168
rect 299348 461128 302056 461156
rect 299348 461116 299354 461128
rect 302050 461116 302056 461128
rect 302108 461156 302114 461168
rect 327350 461156 327356 461168
rect 302108 461128 327356 461156
rect 302108 461116 302114 461128
rect 327350 461116 327356 461128
rect 327408 461116 327414 461168
rect 501874 461116 501880 461168
rect 501932 461156 501938 461168
rect 571426 461156 571432 461168
rect 501932 461128 571432 461156
rect 501932 461116 501938 461128
rect 571426 461116 571432 461128
rect 571484 461156 571490 461168
rect 574646 461156 574652 461168
rect 571484 461128 574652 461156
rect 571484 461116 571490 461128
rect 574646 461116 574652 461128
rect 574704 461116 574710 461168
rect 175228 461048 175234 461100
rect 175286 461088 175292 461100
rect 291838 461088 291844 461100
rect 175286 461060 291844 461088
rect 175286 461048 175292 461060
rect 291838 461048 291844 461060
rect 291896 461048 291902 461100
rect 300302 461048 300308 461100
rect 300360 461088 300366 461100
rect 333514 461088 333520 461100
rect 300360 461060 333520 461088
rect 300360 461048 300366 461060
rect 333514 461048 333520 461060
rect 333572 461048 333578 461100
rect 484210 461048 484216 461100
rect 484268 461088 484274 461100
rect 570322 461088 570328 461100
rect 484268 461060 570328 461088
rect 484268 461048 484274 461060
rect 570322 461048 570328 461060
rect 570380 461048 570386 461100
rect 14826 460980 14832 461032
rect 14884 461020 14890 461032
rect 26234 461020 26240 461032
rect 14884 460992 26240 461020
rect 14884 460980 14890 460992
rect 26234 460980 26240 460992
rect 26292 460980 26298 461032
rect 163636 460980 163642 461032
rect 163694 461020 163700 461032
rect 291470 461020 291476 461032
rect 163694 460992 291476 461020
rect 163694 460980 163700 460992
rect 291470 460980 291476 460992
rect 291528 460980 291534 461032
rect 303522 460980 303528 461032
rect 303580 461020 303586 461032
rect 350902 461020 350908 461032
rect 303580 460992 350908 461020
rect 303580 460980 303586 460992
rect 350902 460980 350908 460992
rect 350960 460980 350966 461032
rect 561582 460980 561588 461032
rect 561640 461020 561646 461032
rect 574186 461020 574192 461032
rect 561640 460992 574192 461020
rect 561640 460980 561646 460992
rect 574186 460980 574192 460992
rect 574244 460980 574250 461032
rect 145926 460952 145932 460964
rect 24872 460924 145932 460952
rect 14918 460844 14924 460896
rect 14976 460884 14982 460896
rect 24872 460884 24900 460924
rect 145926 460912 145932 460924
rect 145984 460912 145990 460964
rect 280706 460912 280712 460964
rect 280764 460952 280770 460964
rect 292482 460952 292488 460964
rect 280764 460924 292488 460952
rect 280764 460912 280770 460924
rect 292482 460912 292488 460924
rect 292540 460912 292546 460964
rect 298738 460912 298744 460964
rect 298796 460952 298802 460964
rect 356698 460952 356704 460964
rect 298796 460924 356704 460952
rect 298796 460912 298802 460924
rect 356698 460912 356704 460924
rect 356756 460912 356762 460964
rect 449434 460912 449440 460964
rect 449492 460952 449498 460964
rect 572898 460952 572904 460964
rect 449492 460924 572904 460952
rect 449492 460912 449498 460924
rect 572898 460912 572904 460924
rect 572956 460912 572962 460964
rect 14976 460856 24900 460884
rect 14976 460844 14982 460856
rect 192938 460844 192944 460896
rect 192996 460884 193002 460896
rect 293954 460884 293960 460896
rect 192996 460856 293960 460884
rect 192996 460844 193002 460856
rect 293954 460844 293960 460856
rect 294012 460844 294018 460896
rect 296530 460844 296536 460896
rect 296588 460884 296594 460896
rect 397270 460884 397276 460896
rect 296588 460856 397276 460884
rect 296588 460844 296594 460856
rect 397270 460844 397276 460856
rect 397328 460844 397334 460896
rect 461026 460844 461032 460896
rect 461084 460884 461090 460896
rect 572990 460884 572996 460896
rect 461084 460856 572996 460884
rect 461084 460844 461090 460856
rect 572990 460844 572996 460856
rect 573048 460844 573054 460896
rect 15010 459620 15016 459672
rect 15068 459660 15074 459672
rect 18690 459660 18696 459672
rect 15068 459632 18696 459660
rect 15068 459620 15074 459632
rect 18690 459620 18696 459632
rect 18748 459620 18754 459672
rect 16298 459552 16304 459604
rect 16356 459592 16362 459604
rect 18598 459592 18604 459604
rect 16356 459564 18604 459592
rect 16356 459552 16362 459564
rect 18598 459552 18604 459564
rect 18656 459552 18662 459604
rect 20254 459552 20260 459604
rect 20312 459592 20318 459604
rect 20312 459564 40080 459592
rect 20312 459552 20318 459564
rect 20622 459484 20628 459536
rect 20680 459524 20686 459536
rect 30006 459524 30012 459536
rect 20680 459496 30012 459524
rect 20680 459484 20686 459496
rect 30006 459484 30012 459496
rect 30064 459484 30070 459536
rect 40052 459524 40080 459564
rect 293954 459552 293960 459604
rect 294012 459592 294018 459604
rect 295426 459592 295432 459604
rect 294012 459564 295432 459592
rect 294012 459552 294018 459564
rect 295426 459552 295432 459564
rect 295484 459552 295490 459604
rect 569310 459552 569316 459604
rect 569368 459592 569374 459604
rect 571610 459592 571616 459604
rect 569368 459564 571616 459592
rect 569368 459552 569374 459564
rect 571610 459552 571616 459564
rect 571668 459552 571674 459604
rect 572990 459552 572996 459604
rect 573048 459592 573054 459604
rect 574278 459592 574284 459604
rect 573048 459564 574284 459592
rect 573048 459552 573054 459564
rect 574278 459552 574284 459564
rect 574336 459552 574342 459604
rect 41598 459524 41604 459536
rect 40052 459496 41604 459524
rect 41598 459484 41604 459496
rect 41656 459484 41662 459536
rect 129182 459484 129188 459536
rect 129240 459524 129246 459536
rect 134334 459524 134340 459536
rect 129240 459496 134340 459524
rect 129240 459484 129246 459496
rect 134334 459484 134340 459496
rect 134392 459484 134398 459536
rect 187142 459484 187148 459536
rect 187200 459524 187206 459536
rect 290274 459524 290280 459536
rect 187200 459496 290280 459524
rect 187200 459484 187206 459496
rect 290274 459484 290280 459496
rect 290332 459484 290338 459536
rect 318794 459484 318800 459536
rect 318852 459524 318858 459536
rect 321922 459524 321928 459536
rect 318852 459496 321928 459524
rect 318852 459484 318858 459496
rect 321922 459484 321928 459496
rect 321980 459484 321986 459536
rect 336734 459484 336740 459536
rect 336792 459524 336798 459536
rect 339310 459524 339316 459536
rect 336792 459496 339316 459524
rect 336792 459484 336798 459496
rect 339310 459484 339316 459496
rect 339368 459484 339374 459536
rect 408862 459484 408868 459536
rect 408920 459524 408926 459536
rect 414658 459524 414664 459536
rect 408920 459496 414664 459524
rect 408920 459484 408926 459496
rect 414658 459484 414664 459496
rect 414716 459484 414722 459536
rect 466822 459484 466828 459536
rect 466880 459524 466886 459536
rect 567930 459524 567936 459536
rect 466880 459496 567936 459524
rect 466880 459484 466886 459496
rect 567930 459484 567936 459496
rect 567988 459524 567994 459536
rect 568482 459524 568488 459536
rect 567988 459496 568488 459524
rect 567988 459484 567994 459496
rect 568482 459484 568488 459496
rect 568540 459484 568546 459536
rect 204162 459416 204168 459468
rect 204220 459456 204226 459468
rect 291378 459456 291384 459468
rect 204220 459428 291384 459456
rect 204220 459416 204226 459428
rect 291378 459416 291384 459428
rect 291436 459416 291442 459468
rect 297818 459416 297824 459468
rect 297876 459456 297882 459468
rect 379882 459456 379888 459468
rect 297876 459428 379888 459456
rect 297876 459416 297882 459428
rect 379882 459416 379888 459428
rect 379940 459416 379946 459468
rect 559558 459416 559564 459468
rect 559616 459456 559622 459468
rect 569954 459456 569960 459468
rect 559616 459428 569960 459456
rect 559616 459416 559622 459428
rect 569954 459416 569960 459428
rect 570012 459416 570018 459468
rect 18598 459348 18604 459400
rect 18656 459388 18662 459400
rect 99558 459388 99564 459400
rect 18656 459360 99564 459388
rect 18656 459348 18662 459360
rect 99558 459348 99564 459360
rect 99616 459348 99622 459400
rect 216122 459348 216128 459400
rect 216180 459388 216186 459400
rect 291194 459388 291200 459400
rect 216180 459360 291200 459388
rect 216180 459348 216186 459360
rect 291194 459348 291200 459360
rect 291252 459348 291258 459400
rect 299014 459348 299020 459400
rect 299072 459388 299078 459400
rect 374086 459388 374092 459400
rect 299072 459360 374092 459388
rect 299072 459348 299078 459360
rect 374086 459348 374092 459360
rect 374144 459348 374150 459400
rect 524782 459348 524788 459400
rect 524840 459388 524846 459400
rect 569310 459388 569316 459400
rect 524840 459360 569316 459388
rect 524840 459348 524846 459360
rect 569310 459348 569316 459360
rect 569368 459348 569374 459400
rect 17770 459280 17776 459332
rect 17828 459320 17834 459332
rect 87966 459320 87972 459332
rect 17828 459292 87972 459320
rect 17828 459280 17834 459292
rect 87966 459280 87972 459292
rect 88024 459280 88030 459332
rect 221918 459280 221924 459332
rect 221976 459320 221982 459332
rect 292758 459320 292764 459332
rect 221976 459292 292764 459320
rect 221976 459280 221982 459292
rect 292758 459280 292764 459292
rect 292816 459280 292822 459332
rect 299382 459280 299388 459332
rect 299440 459320 299446 459332
rect 345106 459320 345112 459332
rect 299440 459292 345112 459320
rect 299440 459280 299446 459292
rect 345106 459280 345112 459292
rect 345164 459280 345170 459332
rect 530578 459280 530584 459332
rect 530636 459320 530642 459332
rect 570230 459320 570236 459332
rect 530636 459292 570236 459320
rect 530636 459280 530642 459292
rect 570230 459280 570236 459292
rect 570288 459280 570294 459332
rect 18690 459212 18696 459264
rect 18748 459252 18754 459264
rect 116946 459252 116952 459264
rect 18748 459224 116952 459252
rect 18748 459212 18754 459224
rect 116946 459212 116952 459224
rect 117004 459212 117010 459264
rect 210326 459212 210332 459264
rect 210384 459252 210390 459264
rect 280706 459252 280712 459264
rect 210384 459224 280712 459252
rect 210384 459212 210390 459224
rect 280706 459212 280712 459224
rect 280764 459212 280770 459264
rect 304994 459212 305000 459264
rect 305052 459252 305058 459264
rect 316126 459252 316132 459264
rect 305052 459224 316132 459252
rect 305052 459212 305058 459224
rect 316126 459212 316132 459224
rect 316184 459212 316190 459264
rect 547966 459212 547972 459264
rect 548024 459252 548030 459264
rect 570138 459252 570144 459264
rect 548024 459224 570144 459252
rect 548024 459212 548030 459224
rect 570138 459212 570144 459224
rect 570196 459212 570202 459264
rect 17586 459144 17592 459196
rect 17644 459184 17650 459196
rect 105354 459184 105360 459196
rect 17644 459156 105360 459184
rect 17644 459144 17650 459156
rect 105354 459144 105360 459156
rect 105412 459144 105418 459196
rect 279878 459144 279884 459196
rect 279936 459184 279942 459196
rect 289998 459184 290004 459196
rect 279936 459156 290004 459184
rect 279936 459144 279942 459156
rect 289998 459144 290004 459156
rect 290056 459144 290062 459196
rect 299198 459144 299204 459196
rect 299256 459184 299262 459196
rect 385678 459184 385684 459196
rect 299256 459156 385684 459184
rect 299256 459144 299262 459156
rect 385678 459144 385684 459156
rect 385736 459144 385742 459196
rect 490006 459144 490012 459196
rect 490064 459184 490070 459196
rect 561582 459184 561588 459196
rect 490064 459156 561588 459184
rect 490064 459144 490070 459156
rect 561582 459144 561588 459156
rect 561640 459144 561646 459196
rect 30926 459008 30932 459060
rect 30984 459048 30990 459060
rect 35894 459048 35900 459060
rect 30984 459020 35900 459048
rect 30984 459008 30990 459020
rect 35894 459008 35900 459020
rect 35952 459008 35958 459060
rect 274082 458872 274088 458924
rect 274140 458912 274146 458924
rect 294690 458912 294696 458924
rect 274140 458884 294696 458912
rect 274140 458872 274146 458884
rect 294690 458872 294696 458884
rect 294748 458872 294754 458924
rect 300394 458872 300400 458924
rect 300452 458912 300458 458924
rect 368290 458912 368296 458924
rect 300452 458884 368296 458912
rect 300452 458872 300458 458884
rect 368290 458872 368296 458884
rect 368348 458872 368354 458924
rect 64874 458844 64880 458856
rect 26206 458816 64880 458844
rect 19242 458668 19248 458720
rect 19300 458708 19306 458720
rect 20530 458708 20536 458720
rect 19300 458680 20536 458708
rect 19300 458668 19306 458680
rect 20530 458668 20536 458680
rect 20588 458708 20594 458720
rect 26206 458708 26234 458816
rect 64874 458804 64880 458816
rect 64932 458804 64938 458856
rect 268286 458804 268292 458856
rect 268344 458844 268350 458856
rect 280062 458844 280068 458856
rect 268344 458816 280068 458844
rect 268344 458804 268350 458816
rect 280062 458804 280068 458816
rect 280120 458804 280126 458856
rect 289078 458804 289084 458856
rect 289136 458844 289142 458856
rect 408862 458844 408868 458856
rect 289136 458816 408868 458844
rect 289136 458804 289142 458816
rect 408862 458804 408868 458816
rect 408920 458804 408926 458856
rect 495802 458804 495808 458856
rect 495860 458844 495866 458856
rect 569310 458844 569316 458856
rect 495860 458816 569316 458844
rect 495860 458804 495866 458816
rect 569310 458804 569316 458816
rect 569368 458844 569374 458856
rect 571702 458844 571708 458856
rect 569368 458816 571708 458844
rect 569368 458804 569374 458816
rect 571702 458804 571708 458816
rect 571760 458804 571766 458856
rect 20588 458680 26234 458708
rect 20588 458668 20594 458680
rect 298830 458668 298836 458720
rect 298888 458708 298894 458720
rect 300394 458708 300400 458720
rect 298888 458680 300400 458708
rect 298888 458668 298894 458680
rect 300394 458668 300400 458680
rect 300452 458668 300458 458720
rect 569954 458532 569960 458584
rect 570012 458572 570018 458584
rect 570414 458572 570420 458584
rect 570012 458544 570420 458572
rect 570012 458532 570018 458544
rect 570414 458532 570420 458544
rect 570472 458532 570478 458584
rect 569954 458396 569960 458448
rect 570012 458436 570018 458448
rect 570138 458436 570144 458448
rect 570012 458408 570144 458436
rect 570012 458396 570018 458408
rect 570138 458396 570144 458408
rect 570196 458396 570202 458448
rect 291194 458260 291200 458312
rect 291252 458300 291258 458312
rect 292850 458300 292856 458312
rect 291252 458272 292856 458300
rect 291252 458260 291258 458272
rect 292850 458260 292856 458272
rect 292908 458260 292914 458312
rect 17494 458192 17500 458244
rect 17552 458232 17558 458244
rect 17770 458232 17776 458244
rect 17552 458204 17776 458232
rect 17552 458192 17558 458204
rect 17770 458192 17776 458204
rect 17828 458192 17834 458244
rect 291378 458192 291384 458244
rect 291436 458232 291442 458244
rect 292666 458232 292672 458244
rect 291436 458204 292672 458232
rect 291436 458192 291442 458204
rect 292666 458192 292672 458204
rect 292724 458192 292730 458244
rect 293310 458192 293316 458244
rect 293368 458232 293374 458244
rect 293954 458232 293960 458244
rect 293368 458204 293960 458232
rect 293368 458192 293374 458204
rect 293954 458192 293960 458204
rect 294012 458192 294018 458244
rect 299106 458192 299112 458244
rect 299164 458232 299170 458244
rect 299382 458232 299388 458244
rect 299164 458204 299388 458232
rect 299164 458192 299170 458204
rect 299382 458192 299388 458204
rect 299440 458192 299446 458244
rect 565354 458192 565360 458244
rect 565412 458232 565418 458244
rect 568942 458232 568948 458244
rect 565412 458204 568948 458232
rect 565412 458192 565418 458204
rect 568942 458192 568948 458204
rect 569000 458192 569006 458244
rect 570230 458192 570236 458244
rect 570288 458232 570294 458244
rect 571518 458232 571524 458244
rect 570288 458204 571524 458232
rect 570288 458192 570294 458204
rect 571518 458192 571524 458204
rect 571576 458192 571582 458244
rect 26234 458124 26240 458176
rect 26292 458164 26298 458176
rect 111150 458164 111156 458176
rect 26292 458136 111156 458164
rect 26292 458124 26298 458136
rect 111150 458124 111156 458136
rect 111208 458124 111214 458176
rect 169662 458124 169668 458176
rect 169720 458164 169726 458176
rect 293328 458164 293356 458192
rect 169720 458136 293356 458164
rect 169720 458124 169726 458136
rect 518986 458124 518992 458176
rect 519044 458164 519050 458176
rect 565814 458164 565820 458176
rect 519044 458136 565820 458164
rect 519044 458124 519050 458136
rect 565814 458124 565820 458136
rect 565872 458124 565878 458176
rect 570414 458124 570420 458176
rect 570472 458164 570478 458176
rect 571702 458164 571708 458176
rect 570472 458136 571708 458164
rect 570472 458124 570478 458136
rect 571702 458124 571708 458136
rect 571760 458124 571766 458176
rect 19150 458056 19156 458108
rect 19208 458096 19214 458108
rect 93854 458096 93860 458108
rect 19208 458068 93860 458096
rect 19208 458056 19214 458068
rect 93854 458056 93860 458068
rect 93912 458056 93918 458108
rect 245102 458056 245108 458108
rect 245160 458096 245166 458108
rect 290090 458096 290096 458108
rect 245160 458068 290096 458096
rect 245160 458056 245166 458068
rect 290090 458056 290096 458068
rect 290148 458056 290154 458108
rect 536374 458056 536380 458108
rect 536432 458096 536438 458108
rect 568666 458096 568672 458108
rect 536432 458068 568672 458096
rect 536432 458056 536438 458068
rect 568666 458056 568672 458068
rect 568724 458056 568730 458108
rect 17678 457988 17684 458040
rect 17736 458028 17742 458040
rect 76374 458028 76380 458040
rect 17736 458000 76380 458028
rect 17736 457988 17742 458000
rect 76374 457988 76380 458000
rect 76432 457988 76438 458040
rect 250898 457988 250904 458040
rect 250956 458028 250962 458040
rect 288618 458028 288624 458040
rect 250956 458000 288624 458028
rect 250956 457988 250962 458000
rect 288618 457988 288624 458000
rect 288676 458028 288682 458040
rect 291378 458028 291384 458040
rect 288676 458000 291384 458028
rect 288676 457988 288682 458000
rect 291378 457988 291384 458000
rect 291436 457988 291442 458040
rect 542170 457988 542176 458040
rect 542228 458028 542234 458040
rect 570046 458028 570052 458040
rect 542228 458000 570052 458028
rect 542228 457988 542234 458000
rect 570046 457988 570052 458000
rect 570104 457988 570110 458040
rect 20438 457920 20444 457972
rect 20496 457960 20502 457972
rect 53190 457960 53196 457972
rect 20496 457932 53196 457960
rect 20496 457920 20502 457932
rect 53190 457920 53196 457932
rect 53248 457920 53254 457972
rect 256602 457920 256608 457972
rect 256660 457960 256666 457972
rect 287606 457960 287612 457972
rect 256660 457932 287612 457960
rect 256660 457920 256666 457932
rect 287606 457920 287612 457932
rect 287664 457960 287670 457972
rect 288434 457960 288440 457972
rect 287664 457932 288440 457960
rect 287664 457920 287670 457932
rect 288434 457920 288440 457932
rect 288492 457920 288498 457972
rect 21910 457852 21916 457904
rect 21968 457892 21974 457904
rect 47394 457892 47400 457904
rect 21968 457864 47400 457892
rect 21968 457852 21974 457864
rect 47394 457852 47400 457864
rect 47452 457852 47458 457904
rect 262122 457852 262128 457904
rect 262180 457892 262186 457904
rect 289814 457892 289820 457904
rect 262180 457864 289820 457892
rect 262180 457852 262186 457864
rect 289814 457852 289820 457864
rect 289872 457852 289878 457904
rect 280062 457444 280068 457496
rect 280120 457484 280126 457496
rect 289170 457484 289176 457496
rect 280120 457456 289176 457484
rect 280120 457444 280126 457456
rect 289170 457444 289176 457456
rect 289228 457484 289234 457496
rect 289906 457484 289912 457496
rect 289228 457456 289912 457484
rect 289228 457444 289234 457456
rect 289906 457444 289912 457456
rect 289964 457444 289970 457496
rect 304994 457444 305000 457496
rect 305052 457484 305058 457496
rect 426434 457484 426440 457496
rect 305052 457456 426440 457484
rect 305052 457444 305058 457456
rect 426434 457444 426440 457456
rect 426492 457444 426498 457496
rect 55950 456832 55956 456884
rect 56008 456872 56014 456884
rect 58986 456872 58992 456884
rect 56008 456844 58992 456872
rect 56008 456832 56014 456844
rect 58986 456832 58992 456844
rect 59044 456832 59050 456884
rect 306374 456696 306380 456748
rect 306432 456736 306438 456748
rect 420454 456736 420460 456748
rect 306432 456708 420460 456736
rect 306432 456696 306438 456708
rect 420454 456696 420460 456708
rect 420512 456696 420518 456748
rect 298002 456492 298008 456544
rect 298060 456532 298066 456544
rect 299198 456532 299204 456544
rect 298060 456504 299204 456532
rect 298060 456492 298066 456504
rect 299198 456492 299204 456504
rect 299256 456532 299262 456544
rect 304994 456532 305000 456544
rect 299256 456504 305000 456532
rect 299256 456492 299262 456504
rect 304994 456492 305000 456504
rect 305052 456492 305058 456544
rect 288250 456288 288256 456340
rect 288308 456328 288314 456340
rect 290182 456328 290188 456340
rect 288308 456300 290188 456328
rect 288308 456288 288314 456300
rect 290182 456288 290188 456300
rect 290240 456288 290246 456340
rect 17862 456016 17868 456068
rect 17920 456056 17926 456068
rect 19150 456056 19156 456068
rect 17920 456028 19156 456056
rect 17920 456016 17926 456028
rect 19150 456016 19156 456028
rect 19208 456056 19214 456068
rect 55950 456056 55956 456068
rect 19208 456028 55956 456056
rect 19208 456016 19214 456028
rect 55950 456016 55956 456028
rect 56008 456016 56014 456068
rect 307662 456016 307668 456068
rect 307720 456056 307726 456068
rect 432046 456056 432052 456068
rect 307720 456028 432052 456056
rect 307720 456016 307726 456028
rect 432046 456016 432052 456028
rect 432104 456016 432110 456068
rect 297910 455336 297916 455388
rect 297968 455376 297974 455388
rect 302234 455376 302240 455388
rect 297968 455348 302240 455376
rect 297968 455336 297974 455348
rect 302234 455336 302240 455348
rect 302292 455376 302298 455388
rect 307662 455376 307668 455388
rect 302292 455348 307668 455376
rect 302292 455336 302298 455348
rect 307662 455336 307668 455348
rect 307720 455336 307726 455388
rect 471974 444320 471980 444372
rect 472032 444360 472038 444372
rect 572806 444360 572812 444372
rect 472032 444332 572812 444360
rect 472032 444320 472038 444332
rect 572806 444320 572812 444332
rect 572864 444320 572870 444372
rect 284294 443640 284300 443692
rect 284352 443680 284358 443692
rect 297358 443680 297364 443692
rect 284352 443652 297364 443680
rect 284352 443640 284358 443652
rect 297358 443640 297364 443652
rect 297416 443640 297422 443692
rect 567102 443640 567108 443692
rect 567160 443680 567166 443692
rect 570230 443680 570236 443692
rect 567160 443652 570236 443680
rect 567160 443640 567166 443652
rect 570230 443640 570236 443652
rect 570288 443640 570294 443692
rect 19058 443368 19064 443420
rect 19116 443408 19122 443420
rect 23474 443408 23480 443420
rect 19116 443380 23480 443408
rect 19116 443368 19122 443380
rect 23474 443368 23480 443380
rect 23532 443368 23538 443420
rect 2866 409912 2872 409964
rect 2924 409952 2930 409964
rect 4890 409952 4896 409964
rect 2924 409924 4896 409952
rect 2924 409912 2930 409924
rect 4890 409912 4896 409924
rect 4948 409912 4954 409964
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 7558 398732 7564 398744
rect 2832 398704 7564 398732
rect 2832 398692 2838 398704
rect 7558 398692 7564 398704
rect 7616 398692 7622 398744
rect 570598 378768 570604 378820
rect 570656 378808 570662 378820
rect 580442 378808 580448 378820
rect 570656 378780 580448 378808
rect 570656 378768 570662 378780
rect 580442 378768 580448 378780
rect 580500 378808 580506 378820
rect 580902 378808 580908 378820
rect 580500 378780 580908 378808
rect 580500 378768 580506 378780
rect 580902 378768 580908 378780
rect 580960 378768 580966 378820
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 18598 357456 18604 357468
rect 3384 357428 18604 357456
rect 3384 357416 3390 357428
rect 18598 357416 18604 357428
rect 18656 357416 18662 357468
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 18690 345080 18696 345092
rect 3384 345052 18696 345080
rect 3384 345040 3390 345052
rect 18690 345040 18696 345052
rect 18748 345040 18754 345092
rect 14918 333956 14924 334008
rect 14976 333996 14982 334008
rect 27522 333996 27528 334008
rect 14976 333968 27528 333996
rect 14976 333956 14982 333968
rect 27522 333956 27528 333968
rect 27580 333956 27586 334008
rect 292482 333956 292488 334008
rect 292540 333996 292546 334008
rect 295610 333996 295616 334008
rect 292540 333968 295616 333996
rect 292540 333956 292546 333968
rect 295610 333956 295616 333968
rect 295668 333956 295674 334008
rect 19150 333276 19156 333328
rect 19208 333316 19214 333328
rect 21818 333316 21824 333328
rect 19208 333288 21824 333316
rect 19208 333276 19214 333288
rect 21818 333276 21824 333288
rect 21876 333316 21882 333328
rect 21876 333288 35894 333316
rect 21876 333276 21882 333288
rect 17402 333208 17408 333260
rect 17460 333248 17466 333260
rect 26234 333248 26240 333260
rect 17460 333220 26240 333248
rect 17460 333208 17466 333220
rect 26234 333208 26240 333220
rect 26292 333208 26298 333260
rect 35866 332976 35894 333288
rect 286962 333276 286968 333328
rect 287020 333316 287026 333328
rect 291470 333316 291476 333328
rect 287020 333288 291476 333316
rect 287020 333276 287026 333288
rect 291470 333276 291476 333288
rect 291528 333276 291534 333328
rect 291746 333276 291752 333328
rect 291804 333316 291810 333328
rect 292850 333316 292856 333328
rect 291804 333288 292856 333316
rect 291804 333276 291810 333288
rect 292850 333276 292856 333288
rect 292908 333276 292914 333328
rect 281442 333208 281448 333260
rect 281500 333248 281506 333260
rect 290274 333248 290280 333260
rect 281500 333220 290280 333248
rect 281500 333208 281506 333220
rect 290274 333208 290280 333220
rect 290332 333208 290338 333260
rect 296622 333208 296628 333260
rect 296680 333248 296686 333260
rect 306374 333248 306380 333260
rect 296680 333220 306380 333248
rect 296680 333208 296686 333220
rect 306374 333208 306380 333220
rect 306432 333208 306438 333260
rect 567102 333208 567108 333260
rect 567160 333248 567166 333260
rect 570322 333248 570328 333260
rect 567160 333220 570328 333248
rect 567160 333208 567166 333220
rect 570322 333208 570328 333220
rect 570380 333208 570386 333260
rect 300210 333140 300216 333192
rect 300268 333180 300274 333192
rect 300762 333180 300768 333192
rect 300268 333152 300768 333180
rect 300268 333140 300274 333152
rect 300762 333140 300768 333152
rect 300820 333140 300826 333192
rect 56502 332976 56508 332988
rect 35866 332948 56508 332976
rect 56502 332936 56508 332948
rect 56560 332936 56566 332988
rect 250898 332936 250904 332988
rect 250956 332976 250962 332988
rect 291286 332976 291292 332988
rect 250956 332948 291292 332976
rect 250956 332936 250962 332948
rect 291286 332936 291292 332948
rect 291344 332936 291350 332988
rect 300762 332936 300768 332988
rect 300820 332976 300826 332988
rect 338942 332976 338948 332988
rect 300820 332948 338948 332976
rect 300820 332936 300826 332948
rect 338942 332936 338948 332948
rect 339000 332936 339006 332988
rect 19058 332868 19064 332920
rect 19116 332908 19122 332920
rect 122742 332908 122748 332920
rect 19116 332880 122748 332908
rect 19116 332868 19122 332880
rect 122742 332868 122748 332880
rect 122800 332868 122806 332920
rect 239306 332868 239312 332920
rect 239364 332908 239370 332920
rect 282178 332908 282184 332920
rect 239364 332880 282184 332908
rect 239364 332868 239370 332880
rect 282178 332868 282184 332880
rect 282236 332868 282242 332920
rect 299106 332868 299112 332920
rect 299164 332908 299170 332920
rect 342254 332908 342260 332920
rect 299164 332880 342260 332908
rect 299164 332868 299170 332880
rect 342254 332868 342260 332880
rect 342312 332868 342318 332920
rect 571334 332908 571340 332920
rect 567166 332880 571340 332908
rect 22002 332800 22008 332852
rect 22060 332840 22066 332852
rect 82170 332840 82176 332852
rect 22060 332812 82176 332840
rect 22060 332800 22066 332812
rect 82170 332800 82176 332812
rect 82228 332800 82234 332852
rect 169754 332800 169760 332852
rect 169812 332840 169818 332852
rect 294046 332840 294052 332852
rect 169812 332812 294052 332840
rect 169812 332800 169818 332812
rect 294046 332800 294052 332812
rect 294104 332800 294110 332852
rect 299014 332800 299020 332852
rect 299072 332840 299078 332852
rect 373902 332840 373908 332852
rect 299072 332812 373908 332840
rect 299072 332800 299078 332812
rect 373902 332800 373908 332812
rect 373960 332800 373966 332852
rect 16298 332732 16304 332784
rect 16356 332772 16362 332784
rect 99558 332772 99564 332784
rect 16356 332744 99564 332772
rect 16356 332732 16362 332744
rect 99558 332732 99564 332744
rect 99616 332732 99622 332784
rect 216122 332732 216128 332784
rect 216180 332772 216186 332784
rect 291746 332772 291752 332784
rect 216180 332744 291752 332772
rect 216180 332732 216186 332744
rect 291746 332732 291752 332744
rect 291804 332732 291810 332784
rect 302050 332732 302056 332784
rect 302108 332772 302114 332784
rect 368290 332772 368296 332784
rect 302108 332744 368296 332772
rect 302108 332732 302114 332744
rect 368290 332732 368296 332744
rect 368348 332732 368354 332784
rect 513190 332732 513196 332784
rect 513248 332772 513254 332784
rect 567166 332772 567194 332880
rect 571334 332868 571340 332880
rect 571392 332868 571398 332920
rect 572806 332772 572812 332784
rect 513248 332744 567194 332772
rect 567304 332744 572812 332772
rect 513248 332732 513254 332744
rect 4982 332664 4988 332716
rect 5040 332704 5046 332716
rect 24210 332704 24216 332716
rect 5040 332676 24216 332704
rect 5040 332664 5046 332676
rect 24210 332664 24216 332676
rect 24268 332664 24274 332716
rect 27522 332664 27528 332716
rect 27580 332704 27586 332716
rect 111150 332704 111156 332716
rect 27580 332676 111156 332704
rect 27580 332664 27586 332676
rect 111150 332664 111156 332676
rect 111208 332664 111214 332716
rect 210326 332664 210332 332716
rect 210384 332704 210390 332716
rect 292482 332704 292488 332716
rect 210384 332676 292488 332704
rect 210384 332664 210390 332676
rect 292482 332664 292488 332676
rect 292540 332664 292546 332716
rect 296254 332664 296260 332716
rect 296312 332704 296318 332716
rect 297818 332704 297824 332716
rect 296312 332676 297824 332704
rect 296312 332664 296318 332676
rect 297818 332664 297824 332676
rect 297876 332704 297882 332716
rect 379882 332704 379888 332716
rect 297876 332676 379888 332704
rect 297876 332664 297882 332676
rect 379882 332664 379888 332676
rect 379940 332664 379946 332716
rect 472618 332664 472624 332716
rect 472676 332704 472682 332716
rect 567304 332704 567332 332744
rect 572806 332732 572812 332744
rect 572864 332772 572870 332784
rect 574554 332772 574560 332784
rect 572864 332744 574560 332772
rect 572864 332732 572870 332744
rect 574554 332732 574560 332744
rect 574612 332732 574618 332784
rect 472676 332676 567332 332704
rect 472676 332664 472682 332676
rect 571334 332664 571340 332716
rect 571392 332704 571398 332716
rect 572990 332704 572996 332716
rect 571392 332676 572996 332704
rect 571392 332664 571398 332676
rect 572990 332664 572996 332676
rect 573048 332664 573054 332716
rect 17586 332596 17592 332648
rect 17644 332636 17650 332648
rect 105354 332636 105360 332648
rect 17644 332608 105360 332636
rect 17644 332596 17650 332608
rect 105354 332596 105360 332608
rect 105412 332596 105418 332648
rect 181346 332596 181352 332648
rect 181404 332636 181410 332648
rect 292574 332636 292580 332648
rect 181404 332608 292580 332636
rect 181404 332596 181410 332608
rect 292574 332596 292580 332608
rect 292632 332636 292638 332648
rect 296714 332636 296720 332648
rect 292632 332608 296720 332636
rect 292632 332596 292638 332608
rect 296714 332596 296720 332608
rect 296772 332596 296778 332648
rect 298830 332596 298836 332648
rect 298888 332636 298894 332648
rect 299014 332636 299020 332648
rect 298888 332608 299020 332636
rect 298888 332596 298894 332608
rect 299014 332596 299020 332608
rect 299072 332596 299078 332648
rect 304534 332596 304540 332648
rect 304592 332636 304598 332648
rect 580350 332636 580356 332648
rect 304592 332608 580356 332636
rect 304592 332596 304598 332608
rect 580350 332596 580356 332608
rect 580408 332596 580414 332648
rect 7650 332528 7656 332580
rect 7708 332568 7714 332580
rect 30006 332568 30012 332580
rect 7708 332540 30012 332568
rect 7708 332528 7714 332540
rect 30006 332528 30012 332540
rect 30064 332528 30070 332580
rect 31018 332568 31024 332580
rect 30576 332540 31024 332568
rect 21910 332460 21916 332512
rect 21968 332500 21974 332512
rect 30576 332500 30604 332540
rect 31018 332528 31024 332540
rect 31076 332528 31082 332580
rect 56502 332528 56508 332580
rect 56560 332568 56566 332580
rect 58986 332568 58992 332580
rect 56560 332540 58992 332568
rect 56560 332528 56566 332540
rect 58986 332528 58992 332540
rect 59044 332528 59050 332580
rect 129182 332528 129188 332580
rect 129240 332568 129246 332580
rect 134978 332568 134984 332580
rect 129240 332540 134984 332568
rect 129240 332528 129246 332540
rect 134978 332528 134984 332540
rect 135036 332528 135042 332580
rect 256602 332528 256608 332580
rect 256660 332568 256666 332580
rect 287790 332568 287796 332580
rect 256660 332540 287796 332568
rect 256660 332528 256666 332540
rect 287790 332528 287796 332540
rect 287848 332528 287854 332580
rect 342254 332528 342260 332580
rect 342312 332568 342318 332580
rect 345106 332568 345112 332580
rect 342312 332540 345112 332568
rect 342312 332528 342318 332540
rect 345106 332528 345112 332540
rect 345164 332528 345170 332580
rect 408862 332528 408868 332580
rect 408920 332568 408926 332580
rect 414658 332568 414664 332580
rect 408920 332540 414664 332568
rect 408920 332528 408926 332540
rect 414658 332528 414664 332540
rect 414716 332528 414722 332580
rect 524782 332528 524788 332580
rect 524840 332568 524846 332580
rect 571610 332568 571616 332580
rect 524840 332540 571616 332568
rect 524840 332528 524846 332540
rect 571610 332528 571616 332540
rect 571668 332528 571674 332580
rect 64966 332500 64972 332512
rect 21968 332472 30604 332500
rect 30668 332472 64972 332500
rect 21968 332460 21974 332472
rect 20530 332392 20536 332444
rect 20588 332432 20594 332444
rect 30668 332432 30696 332472
rect 64966 332460 64972 332472
rect 65024 332460 65030 332512
rect 262122 332460 262128 332512
rect 262180 332500 262186 332512
rect 289814 332500 289820 332512
rect 262180 332472 289820 332500
rect 262180 332460 262186 332472
rect 289814 332460 289820 332472
rect 289872 332460 289878 332512
rect 300302 332460 300308 332512
rect 300360 332500 300366 332512
rect 333514 332500 333520 332512
rect 300360 332472 333520 332500
rect 300360 332460 300366 332472
rect 333514 332460 333520 332472
rect 333572 332460 333578 332512
rect 518986 332460 518992 332512
rect 519044 332500 519050 332512
rect 565814 332500 565820 332512
rect 519044 332472 565820 332500
rect 519044 332460 519050 332472
rect 565814 332460 565820 332472
rect 565872 332460 565878 332512
rect 53190 332432 53196 332444
rect 20588 332404 30696 332432
rect 30760 332404 53196 332432
rect 20588 332392 20594 332404
rect 20438 332324 20444 332376
rect 20496 332364 20502 332376
rect 30760 332364 30788 332404
rect 53190 332392 53196 332404
rect 53248 332392 53254 332444
rect 268286 332392 268292 332444
rect 268344 332432 268350 332444
rect 289170 332432 289176 332444
rect 268344 332404 289176 332432
rect 268344 332392 268350 332404
rect 289170 332392 289176 332404
rect 289228 332432 289234 332444
rect 293034 332432 293040 332444
rect 289228 332404 293040 332432
rect 289228 332392 289234 332404
rect 293034 332392 293040 332404
rect 293092 332392 293098 332444
rect 299290 332392 299296 332444
rect 299348 332432 299354 332444
rect 327718 332432 327724 332444
rect 299348 332404 327724 332432
rect 299348 332392 299354 332404
rect 327718 332392 327724 332404
rect 327776 332392 327782 332444
rect 536374 332392 536380 332444
rect 536432 332432 536438 332444
rect 568666 332432 568672 332444
rect 536432 332404 568672 332432
rect 536432 332392 536438 332404
rect 568666 332392 568672 332404
rect 568724 332392 568730 332444
rect 20496 332336 30788 332364
rect 20496 332324 20502 332336
rect 31018 332324 31024 332376
rect 31076 332364 31082 332376
rect 47394 332364 47400 332376
rect 31076 332336 47400 332364
rect 31076 332324 31082 332336
rect 47394 332324 47400 332336
rect 47452 332324 47458 332376
rect 279878 332324 279884 332376
rect 279936 332364 279942 332376
rect 289998 332364 290004 332376
rect 279936 332336 290004 332364
rect 279936 332324 279942 332336
rect 289998 332324 290004 332336
rect 290056 332324 290062 332376
rect 302142 332324 302148 332376
rect 302200 332364 302206 332376
rect 321922 332364 321928 332376
rect 302200 332336 321928 332364
rect 302200 332324 302206 332336
rect 321922 332324 321928 332336
rect 321980 332324 321986 332376
rect 542170 332324 542176 332376
rect 542228 332364 542234 332376
rect 570046 332364 570052 332376
rect 542228 332336 570052 332364
rect 542228 332324 542234 332336
rect 570046 332324 570052 332336
rect 570104 332324 570110 332376
rect 20254 332256 20260 332308
rect 20312 332296 20318 332308
rect 41598 332296 41604 332308
rect 20312 332268 41604 332296
rect 20312 332256 20318 332268
rect 41598 332256 41604 332268
rect 41656 332256 41662 332308
rect 300578 332256 300584 332308
rect 300636 332296 300642 332308
rect 316126 332296 316132 332308
rect 300636 332268 316132 332296
rect 300636 332256 300642 332268
rect 316126 332256 316132 332268
rect 316184 332256 316190 332308
rect 547966 332256 547972 332308
rect 548024 332296 548030 332308
rect 569954 332296 569960 332308
rect 548024 332268 569960 332296
rect 548024 332256 548030 332268
rect 569954 332256 569960 332268
rect 570012 332256 570018 332308
rect 20346 332188 20352 332240
rect 20404 332228 20410 332240
rect 35986 332228 35992 332240
rect 20404 332200 35992 332228
rect 20404 332188 20410 332200
rect 35986 332188 35992 332200
rect 36044 332188 36050 332240
rect 303522 332188 303528 332240
rect 303580 332228 303586 332240
rect 350902 332228 350908 332240
rect 303580 332200 350908 332228
rect 303580 332188 303586 332200
rect 350902 332188 350908 332200
rect 350960 332188 350966 332240
rect 559558 332188 559564 332240
rect 559616 332228 559622 332240
rect 571886 332228 571892 332240
rect 559616 332200 571892 332228
rect 559616 332188 559622 332200
rect 571886 332188 571892 332200
rect 571944 332188 571950 332240
rect 23382 332120 23388 332172
rect 23440 332160 23446 332172
rect 70578 332160 70584 332172
rect 23440 332132 70584 332160
rect 23440 332120 23446 332132
rect 70578 332120 70584 332132
rect 70636 332120 70642 332172
rect 289814 332052 289820 332104
rect 289872 332092 289878 332104
rect 293954 332092 293960 332104
rect 289872 332064 293960 332092
rect 289872 332052 289878 332064
rect 293954 332052 293960 332064
rect 294012 332052 294018 332104
rect 285582 331984 285588 332036
rect 285640 332024 285646 332036
rect 290550 332024 290556 332036
rect 285640 331996 290556 332024
rect 285640 331984 285646 331996
rect 290550 331984 290556 331996
rect 290608 331984 290614 332036
rect 198642 331916 198648 331968
rect 198700 331956 198706 331968
rect 289814 331956 289820 331968
rect 198700 331928 289820 331956
rect 198700 331916 198706 331928
rect 289814 331916 289820 331928
rect 289872 331916 289878 331968
rect 290458 331916 290464 331968
rect 290516 331956 290522 331968
rect 408862 331956 408868 331968
rect 290516 331928 408868 331956
rect 290516 331916 290522 331928
rect 408862 331916 408868 331928
rect 408920 331916 408926 331968
rect 443638 331916 443644 331968
rect 443696 331956 443702 331968
rect 561582 331956 561588 331968
rect 443696 331928 561588 331956
rect 443696 331916 443702 331928
rect 561582 331916 561588 331928
rect 561640 331916 561646 331968
rect 134978 331848 134984 331900
rect 135036 331888 135042 331900
rect 288434 331888 288440 331900
rect 135036 331860 288440 331888
rect 135036 331848 135042 331860
rect 288434 331848 288440 331860
rect 288492 331848 288498 331900
rect 297450 331848 297456 331900
rect 297508 331888 297514 331900
rect 478414 331888 478420 331900
rect 297508 331860 478420 331888
rect 297508 331848 297514 331860
rect 478414 331848 478420 331860
rect 478472 331848 478478 331900
rect 565354 331848 565360 331900
rect 565412 331888 565418 331900
rect 571334 331888 571340 331900
rect 565412 331860 571340 331888
rect 565412 331848 565418 331860
rect 571334 331848 571340 331860
rect 571392 331848 571398 331900
rect 282178 331712 282184 331764
rect 282236 331752 282242 331764
rect 285582 331752 285588 331764
rect 282236 331724 285588 331752
rect 282236 331712 282242 331724
rect 285582 331712 285588 331724
rect 285640 331712 285646 331764
rect 20070 331372 20076 331424
rect 20128 331412 20134 331424
rect 20438 331412 20444 331424
rect 20128 331384 20444 331412
rect 20128 331372 20134 331384
rect 20438 331372 20444 331384
rect 20496 331372 20502 331424
rect 20162 331304 20168 331356
rect 20220 331344 20226 331356
rect 20530 331344 20536 331356
rect 20220 331316 20536 331344
rect 20220 331304 20226 331316
rect 20530 331304 20536 331316
rect 20588 331304 20594 331356
rect 20438 331236 20444 331288
rect 20496 331276 20502 331288
rect 21910 331276 21916 331288
rect 20496 331248 21916 331276
rect 20496 331236 20502 331248
rect 21910 331236 21916 331248
rect 21968 331236 21974 331288
rect 245102 331236 245108 331288
rect 245160 331276 245166 331288
rect 246298 331276 246304 331288
rect 245160 331248 246304 331276
rect 245160 331236 245166 331248
rect 246298 331236 246304 331248
rect 246356 331236 246362 331288
rect 299014 331236 299020 331288
rect 299072 331276 299078 331288
rect 299290 331276 299296 331288
rect 299072 331248 299296 331276
rect 299072 331236 299078 331248
rect 299290 331236 299296 331248
rect 299348 331236 299354 331288
rect 453942 331236 453948 331288
rect 454000 331276 454006 331288
rect 455230 331276 455236 331288
rect 454000 331248 455236 331276
rect 454000 331236 454006 331248
rect 455230 331236 455236 331248
rect 455288 331236 455294 331288
rect 482922 331236 482928 331288
rect 482980 331276 482986 331288
rect 484210 331276 484216 331288
rect 482980 331248 484216 331276
rect 482980 331236 482986 331248
rect 484210 331236 484216 331248
rect 484268 331236 484274 331288
rect 571610 331236 571616 331288
rect 571668 331276 571674 331288
rect 573082 331276 573088 331288
rect 571668 331248 573088 331276
rect 571668 331236 571674 331248
rect 573082 331236 573088 331248
rect 573140 331236 573146 331288
rect 192938 331168 192944 331220
rect 192996 331208 193002 331220
rect 295426 331208 295432 331220
rect 192996 331180 295432 331208
rect 192996 331168 193002 331180
rect 295426 331168 295432 331180
rect 295484 331168 295490 331220
rect 561582 331168 561588 331220
rect 561640 331208 561646 331220
rect 575566 331208 575572 331220
rect 561640 331180 575572 331208
rect 561640 331168 561646 331180
rect 575566 331168 575572 331180
rect 575624 331208 575630 331220
rect 576210 331208 576216 331220
rect 575624 331180 576216 331208
rect 575624 331168 575630 331180
rect 576210 331168 576216 331180
rect 576268 331168 576274 331220
rect 221918 331100 221924 331152
rect 221976 331140 221982 331152
rect 292758 331140 292764 331152
rect 221976 331112 292764 331140
rect 221976 331100 221982 331112
rect 292758 331100 292764 331112
rect 292816 331100 292822 331152
rect 24854 330488 24860 330540
rect 24912 330528 24918 330540
rect 145926 330528 145932 330540
rect 24912 330500 145932 330528
rect 24912 330488 24918 330500
rect 145926 330488 145932 330500
rect 145984 330488 145990 330540
rect 204162 330488 204168 330540
rect 204220 330528 204226 330540
rect 289722 330528 289728 330540
rect 204220 330500 289728 330528
rect 204220 330488 204226 330500
rect 289722 330488 289728 330500
rect 289780 330528 289786 330540
rect 292666 330528 292672 330540
rect 289780 330500 292672 330528
rect 289780 330488 289786 330500
rect 292666 330488 292672 330500
rect 292724 330488 292730 330540
rect 299198 330488 299204 330540
rect 299256 330528 299262 330540
rect 307662 330528 307668 330540
rect 299256 330500 307668 330528
rect 299256 330488 299262 330500
rect 307662 330488 307668 330500
rect 307720 330488 307726 330540
rect 576210 330352 576216 330404
rect 576268 330392 576274 330404
rect 576854 330392 576860 330404
rect 576268 330364 576860 330392
rect 576268 330352 576274 330364
rect 576854 330352 576860 330364
rect 576912 330352 576918 330404
rect 15010 329740 15016 329792
rect 15068 329780 15074 329792
rect 116946 329780 116952 329792
rect 15068 329752 116952 329780
rect 15068 329740 15074 329752
rect 116946 329740 116952 329752
rect 117004 329740 117010 329792
rect 307662 329740 307668 329792
rect 307720 329780 307726 329792
rect 425698 329780 425704 329792
rect 307720 329752 425704 329780
rect 307720 329740 307726 329752
rect 425698 329740 425704 329752
rect 425756 329780 425762 329792
rect 426250 329780 426256 329792
rect 425756 329752 426256 329780
rect 425756 329740 425762 329752
rect 426250 329740 426256 329752
rect 426308 329740 426314 329792
rect 461026 329740 461032 329792
rect 461084 329780 461090 329792
rect 574278 329780 574284 329792
rect 461084 329752 574284 329780
rect 461084 329740 461090 329752
rect 574278 329740 574284 329752
rect 574336 329740 574342 329792
rect 574462 329740 574468 329792
rect 574520 329780 574526 329792
rect 575658 329780 575664 329792
rect 574520 329752 575664 329780
rect 574520 329740 574526 329752
rect 575658 329740 575664 329752
rect 575716 329740 575722 329792
rect 17494 329672 17500 329724
rect 17552 329712 17558 329724
rect 87966 329712 87972 329724
rect 17552 329684 87972 329712
rect 17552 329672 17558 329684
rect 87966 329672 87972 329684
rect 88024 329672 88030 329724
rect 490006 329672 490012 329724
rect 490064 329712 490070 329724
rect 574480 329712 574508 329740
rect 490064 329684 574508 329712
rect 490064 329672 490070 329684
rect 15102 329604 15108 329656
rect 15160 329644 15166 329656
rect 24854 329644 24860 329656
rect 15160 329616 24860 329644
rect 15160 329604 15166 329616
rect 24854 329604 24860 329616
rect 24912 329604 24918 329656
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 17218 318832 17224 318844
rect 3384 318804 17224 318832
rect 3384 318792 3390 318804
rect 17218 318792 17224 318804
rect 17276 318792 17282 318844
rect 437474 318112 437480 318164
rect 437532 318152 437538 318164
rect 562318 318152 562324 318164
rect 437532 318124 562324 318152
rect 437532 318112 437538 318124
rect 562318 318112 562324 318124
rect 562376 318112 562382 318164
rect 307662 318044 307668 318096
rect 307720 318084 307726 318096
rect 431954 318084 431960 318096
rect 307720 318056 431960 318084
rect 307720 318044 307726 318056
rect 431954 318044 431960 318056
rect 432012 318084 432018 318096
rect 578234 318084 578240 318096
rect 432012 318056 578240 318084
rect 432012 318044 432018 318056
rect 578234 318044 578240 318056
rect 578292 318044 578298 318096
rect 298738 317432 298744 317484
rect 298796 317472 298802 317484
rect 304994 317472 305000 317484
rect 298796 317444 305000 317472
rect 298796 317432 298802 317444
rect 304994 317432 305000 317444
rect 305052 317432 305058 317484
rect 297910 317364 297916 317416
rect 297968 317404 297974 317416
rect 307662 317404 307668 317416
rect 297968 317376 307668 317404
rect 297968 317364 297974 317376
rect 307662 317364 307668 317376
rect 307720 317364 307726 317416
rect 562318 317364 562324 317416
rect 562376 317404 562382 317416
rect 575474 317404 575480 317416
rect 562376 317376 575480 317404
rect 562376 317364 562382 317376
rect 575474 317364 575480 317376
rect 575532 317364 575538 317416
rect 425698 316684 425704 316736
rect 425756 316724 425762 316736
rect 565814 316724 565820 316736
rect 425756 316696 565820 316724
rect 425756 316684 425762 316696
rect 565814 316684 565820 316696
rect 565872 316684 565878 316736
rect 281442 316004 281448 316056
rect 281500 316044 281506 316056
rect 295518 316044 295524 316056
rect 281500 316016 295524 316044
rect 281500 316004 281506 316016
rect 295518 316004 295524 316016
rect 295576 316004 295582 316056
rect 26326 315936 26332 315988
rect 26384 315976 26390 315988
rect 139394 315976 139400 315988
rect 26384 315948 139400 315976
rect 26384 315936 26390 315948
rect 139394 315936 139400 315948
rect 139452 315936 139458 315988
rect 157334 315936 157340 315988
rect 157392 315976 157398 315988
rect 280798 315976 280804 315988
rect 157392 315948 280804 315976
rect 157392 315936 157398 315948
rect 280798 315936 280804 315948
rect 280856 315936 280862 315988
rect 19242 315868 19248 315920
rect 19300 315908 19306 315920
rect 93854 315908 93860 315920
rect 19300 315880 93860 315908
rect 19300 315868 19306 315880
rect 93854 315868 93860 315880
rect 93912 315868 93918 315920
rect 186222 315868 186228 315920
rect 186280 315908 186286 315920
rect 281460 315908 281488 316004
rect 304994 315936 305000 315988
rect 305052 315976 305058 315988
rect 419534 315976 419540 315988
rect 305052 315948 419540 315976
rect 305052 315936 305058 315948
rect 419534 315936 419540 315948
rect 419592 315936 419598 315988
rect 448514 315936 448520 315988
rect 448572 315976 448578 315988
rect 572898 315976 572904 315988
rect 448572 315948 572904 315976
rect 448572 315936 448578 315948
rect 572898 315936 572904 315948
rect 572956 315936 572962 315988
rect 186280 315880 281488 315908
rect 186280 315868 186286 315880
rect 300118 315868 300124 315920
rect 300176 315908 300182 315920
rect 402974 315908 402980 315920
rect 300176 315880 402980 315908
rect 300176 315868 300182 315880
rect 402974 315868 402980 315880
rect 403032 315868 403038 315920
rect 482922 315868 482928 315920
rect 482980 315908 482986 315920
rect 567102 315908 567108 315920
rect 482980 315880 567108 315908
rect 482980 315868 482986 315880
rect 567102 315868 567108 315880
rect 567160 315868 567166 315920
rect 226334 315800 226340 315852
rect 226392 315840 226398 315852
rect 288526 315840 288532 315852
rect 226392 315812 288532 315840
rect 226392 315800 226398 315812
rect 288526 315800 288532 315812
rect 288584 315800 288590 315852
rect 296346 315800 296352 315852
rect 296404 315840 296410 315852
rect 396074 315840 396080 315852
rect 296404 315812 396080 315840
rect 296404 315800 296410 315812
rect 396074 315800 396080 315812
rect 396132 315800 396138 315852
rect 495434 315800 495440 315852
rect 495492 315840 495498 315852
rect 569310 315840 569316 315852
rect 495492 315812 569316 315840
rect 495492 315800 495498 315812
rect 569310 315800 569316 315812
rect 569368 315800 569374 315852
rect 231854 315732 231860 315784
rect 231912 315772 231918 315784
rect 291562 315772 291568 315784
rect 231912 315744 291568 315772
rect 231912 315732 231918 315744
rect 291562 315732 291568 315744
rect 291620 315732 291626 315784
rect 307662 315732 307668 315784
rect 307720 315772 307726 315784
rect 390554 315772 390560 315784
rect 307720 315744 390560 315772
rect 307720 315732 307726 315744
rect 390554 315732 390560 315744
rect 390612 315732 390618 315784
rect 500862 315732 500868 315784
rect 500920 315772 500926 315784
rect 574646 315772 574652 315784
rect 500920 315744 574652 315772
rect 500920 315732 500926 315744
rect 574646 315732 574652 315744
rect 574704 315732 574710 315784
rect 246298 315664 246304 315716
rect 246356 315704 246362 315716
rect 290090 315704 290096 315716
rect 246356 315676 290096 315704
rect 246356 315664 246362 315676
rect 290090 315664 290096 315676
rect 290148 315664 290154 315716
rect 302050 315664 302056 315716
rect 302108 315704 302114 315716
rect 361574 315704 361580 315716
rect 302108 315676 361580 315704
rect 302108 315664 302114 315676
rect 361574 315664 361580 315676
rect 361632 315664 361638 315716
rect 506474 315664 506480 315716
rect 506532 315704 506538 315716
rect 567470 315704 567476 315716
rect 506532 315676 567476 315704
rect 506532 315664 506538 315676
rect 567470 315664 567476 315676
rect 567528 315664 567534 315716
rect 298922 315596 298928 315648
rect 298980 315636 298986 315648
rect 356054 315636 356060 315648
rect 298980 315608 356060 315636
rect 298980 315596 298986 315608
rect 356054 315596 356060 315608
rect 356112 315596 356118 315648
rect 529934 315596 529940 315648
rect 529992 315636 529998 315648
rect 571794 315636 571800 315648
rect 529992 315608 571800 315636
rect 529992 315596 529998 315608
rect 571794 315596 571800 315608
rect 571852 315596 571858 315648
rect 14826 315392 14832 315444
rect 14884 315432 14890 315444
rect 26326 315432 26332 315444
rect 14884 315404 26332 315432
rect 14884 315392 14890 315404
rect 26326 315392 26332 315404
rect 26384 315392 26390 315444
rect 27522 315324 27528 315376
rect 27580 315364 27586 315376
rect 151814 315364 151820 315376
rect 27580 315336 151820 315364
rect 27580 315324 27586 315336
rect 151814 315324 151820 315336
rect 151872 315324 151878 315376
rect 285582 315324 285588 315376
rect 285640 315364 285646 315376
rect 292942 315364 292948 315376
rect 285640 315336 292948 315364
rect 285640 315324 285646 315336
rect 292942 315324 292948 315336
rect 293000 315324 293006 315376
rect 298002 315324 298008 315376
rect 298060 315364 298066 315376
rect 306374 315364 306380 315376
rect 298060 315336 306380 315364
rect 298060 315324 298066 315336
rect 306374 315324 306380 315336
rect 306432 315364 306438 315376
rect 307662 315364 307668 315376
rect 306432 315336 307668 315364
rect 306432 315324 306438 315336
rect 307662 315324 307668 315336
rect 307720 315324 307726 315376
rect 17586 315256 17592 315308
rect 17644 315296 17650 315308
rect 157334 315296 157340 315308
rect 17644 315268 157340 315296
rect 17644 315256 17650 315268
rect 157334 315256 157340 315268
rect 157392 315256 157398 315308
rect 273254 315256 273260 315308
rect 273312 315296 273318 315308
rect 297542 315296 297548 315308
rect 273312 315268 297548 315296
rect 273312 315256 273318 315268
rect 297542 315256 297548 315268
rect 297600 315256 297606 315308
rect 298094 315256 298100 315308
rect 298152 315296 298158 315308
rect 385034 315296 385040 315308
rect 298152 315268 385040 315296
rect 298152 315256 298158 315268
rect 385034 315256 385040 315268
rect 385092 315256 385098 315308
rect 466454 315256 466460 315308
rect 466512 315296 466518 315308
rect 571426 315296 571432 315308
rect 466512 315268 571432 315296
rect 466512 315256 466518 315268
rect 571426 315256 571432 315268
rect 571484 315256 571490 315308
rect 300118 315052 300124 315104
rect 300176 315092 300182 315104
rect 300394 315092 300400 315104
rect 300176 315064 300400 315092
rect 300176 315052 300182 315064
rect 300394 315052 300400 315064
rect 300452 315052 300458 315104
rect 572898 314712 572904 314764
rect 572956 314752 572962 314764
rect 576946 314752 576952 314764
rect 572956 314724 576952 314752
rect 572956 314712 572962 314724
rect 576946 314712 576952 314724
rect 577004 314712 577010 314764
rect 290090 314644 290096 314696
rect 290148 314684 290154 314696
rect 291194 314684 291200 314696
rect 290148 314656 291200 314684
rect 290148 314644 290154 314656
rect 291194 314644 291200 314656
rect 291252 314644 291258 314696
rect 291562 314644 291568 314696
rect 291620 314684 291626 314696
rect 292850 314684 292856 314696
rect 291620 314656 292856 314684
rect 291620 314644 291626 314656
rect 292850 314644 292856 314656
rect 292908 314644 292914 314696
rect 298922 314644 298928 314696
rect 298980 314684 298986 314696
rect 299290 314684 299296 314696
rect 298980 314656 299296 314684
rect 298980 314644 298986 314656
rect 299290 314644 299296 314656
rect 299348 314644 299354 314696
rect 567102 314644 567108 314696
rect 567160 314684 567166 314696
rect 568850 314684 568856 314696
rect 567160 314656 568856 314684
rect 567160 314644 567166 314656
rect 568850 314644 568856 314656
rect 568908 314644 568914 314696
rect 569310 314644 569316 314696
rect 569368 314684 569374 314696
rect 571518 314684 571524 314696
rect 569368 314656 571524 314684
rect 569368 314644 569374 314656
rect 571518 314644 571524 314656
rect 571576 314644 571582 314696
rect 574186 314644 574192 314696
rect 574244 314684 574250 314696
rect 574646 314684 574652 314696
rect 574244 314656 574652 314684
rect 574244 314644 574250 314656
rect 574646 314644 574652 314656
rect 574704 314644 574710 314696
rect 16390 314576 16396 314628
rect 16448 314616 16454 314628
rect 27522 314616 27528 314628
rect 16448 314588 27528 314616
rect 16448 314576 16454 314588
rect 27522 314576 27528 314588
rect 27580 314576 27586 314628
rect 162854 314576 162860 314628
rect 162912 314616 162918 314628
rect 285766 314616 285772 314628
rect 162912 314588 285772 314616
rect 162912 314576 162918 314588
rect 285766 314576 285772 314588
rect 285824 314576 285830 314628
rect 453942 314576 453948 314628
rect 454000 314616 454006 314628
rect 568482 314616 568488 314628
rect 454000 314588 568488 314616
rect 454000 314576 454006 314588
rect 568482 314576 568488 314588
rect 568540 314616 568546 314628
rect 571702 314616 571708 314628
rect 568540 314588 571708 314616
rect 568540 314576 568546 314588
rect 571702 314576 571708 314588
rect 571760 314576 571766 314628
rect 285766 313896 285772 313948
rect 285824 313936 285830 313948
rect 286962 313936 286968 313948
rect 285824 313908 286968 313936
rect 285824 313896 285830 313908
rect 286962 313896 286968 313908
rect 287020 313936 287026 313948
rect 296714 313936 296720 313948
rect 287020 313908 296720 313936
rect 287020 313896 287026 313908
rect 296714 313896 296720 313908
rect 296772 313896 296778 313948
rect 565814 313896 565820 313948
rect 565872 313936 565878 313948
rect 575474 313936 575480 313948
rect 565872 313908 575480 313936
rect 565872 313896 565878 313908
rect 575474 313896 575480 313908
rect 575532 313896 575538 313948
rect 289722 313284 289728 313336
rect 289780 313324 289786 313336
rect 289906 313324 289912 313336
rect 289780 313296 289912 313324
rect 289780 313284 289786 313296
rect 289906 313284 289912 313296
rect 289964 313284 289970 313336
rect 571242 313284 571248 313336
rect 571300 313324 571306 313336
rect 571426 313324 571432 313336
rect 571300 313296 571432 313324
rect 571300 313284 571306 313296
rect 571426 313284 571432 313296
rect 571484 313284 571490 313336
rect 2774 292612 2780 292664
rect 2832 292652 2838 292664
rect 4982 292652 4988 292664
rect 2832 292624 4988 292652
rect 2832 292612 2838 292624
rect 4982 292612 4988 292624
rect 5040 292612 5046 292664
rect 3142 266432 3148 266484
rect 3200 266472 3206 266484
rect 6178 266472 6184 266484
rect 3200 266444 6184 266472
rect 3200 266432 3206 266444
rect 6178 266432 6184 266444
rect 6236 266432 6242 266484
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 5074 240224 5080 240236
rect 2832 240196 5080 240224
rect 2832 240184 2838 240196
rect 5074 240184 5080 240196
rect 5132 240184 5138 240236
rect 2958 213936 2964 213988
rect 3016 213976 3022 213988
rect 6270 213976 6276 213988
rect 3016 213948 6276 213976
rect 3016 213936 3022 213948
rect 6270 213936 6276 213948
rect 6328 213936 6334 213988
rect 300394 206592 300400 206644
rect 300452 206632 300458 206644
rect 307018 206632 307024 206644
rect 300452 206604 307024 206632
rect 300452 206592 300458 206604
rect 307018 206592 307024 206604
rect 307076 206592 307082 206644
rect 560202 206320 560208 206372
rect 560260 206360 560266 206372
rect 571702 206360 571708 206372
rect 560260 206332 571708 206360
rect 560260 206320 560266 206332
rect 571702 206320 571708 206332
rect 571760 206320 571766 206372
rect 14918 206252 14924 206304
rect 14976 206292 14982 206304
rect 24946 206292 24952 206304
rect 14976 206264 24952 206292
rect 14976 206252 14982 206264
rect 24946 206252 24952 206264
rect 25004 206252 25010 206304
rect 495434 206252 495440 206304
rect 495492 206292 495498 206304
rect 575474 206292 575480 206304
rect 495492 206264 575480 206292
rect 495492 206252 495498 206264
rect 575474 206252 575480 206264
rect 575532 206252 575538 206304
rect 298002 205708 298008 205760
rect 298060 205748 298066 205760
rect 304994 205748 305000 205760
rect 298060 205720 305000 205748
rect 298060 205708 298066 205720
rect 304994 205708 305000 205720
rect 305052 205708 305058 205760
rect 302878 205640 302884 205692
rect 302936 205680 302942 205692
rect 310422 205680 310428 205692
rect 302936 205652 310428 205680
rect 302936 205640 302942 205652
rect 310422 205640 310428 205652
rect 310480 205640 310486 205692
rect 283282 204960 283288 205012
rect 283340 205000 283346 205012
rect 289998 205000 290004 205012
rect 283340 204972 290004 205000
rect 283340 204960 283346 204972
rect 289998 204960 290004 204972
rect 290056 205000 290062 205012
rect 293126 205000 293132 205012
rect 290056 204972 293132 205000
rect 290056 204960 290062 204972
rect 293126 204960 293132 204972
rect 293184 204960 293190 205012
rect 540882 204960 540888 205012
rect 540940 205000 540946 205012
rect 578234 205000 578240 205012
rect 540940 204972 578240 205000
rect 540940 204960 540946 204972
rect 578234 204960 578240 204972
rect 578292 204960 578298 205012
rect 14826 204892 14832 204944
rect 14884 204932 14890 204944
rect 24854 204932 24860 204944
rect 14884 204904 24860 204932
rect 14884 204892 14890 204904
rect 24854 204892 24860 204904
rect 24912 204892 24918 204944
rect 289170 204892 289176 204944
rect 289228 204932 289234 204944
rect 295518 204932 295524 204944
rect 289228 204904 295524 204932
rect 289228 204892 289234 204904
rect 295518 204892 295524 204904
rect 295576 204892 295582 204944
rect 296530 204892 296536 204944
rect 296588 204932 296594 204944
rect 298830 204932 298836 204944
rect 296588 204904 298836 204932
rect 296588 204892 296594 204904
rect 298830 204892 298836 204904
rect 298888 204932 298894 204944
rect 373994 204932 374000 204944
rect 298888 204904 374000 204932
rect 298888 204892 298894 204904
rect 373994 204892 374000 204904
rect 374052 204892 374058 204944
rect 467098 204892 467104 204944
rect 467156 204932 467162 204944
rect 571242 204932 571248 204944
rect 467156 204904 571248 204932
rect 467156 204892 467162 204904
rect 571242 204892 571248 204904
rect 571300 204932 571306 204944
rect 575474 204932 575480 204944
rect 571300 204904 575480 204932
rect 571300 204892 571306 204904
rect 575474 204892 575480 204904
rect 575532 204892 575538 204944
rect 292758 204756 292764 204808
rect 292816 204796 292822 204808
rect 295334 204796 295340 204808
rect 292816 204768 295340 204796
rect 292816 204756 292822 204768
rect 295334 204756 295340 204768
rect 295392 204756 295398 204808
rect 571426 204756 571432 204808
rect 571484 204796 571490 204808
rect 571794 204796 571800 204808
rect 571484 204768 571800 204796
rect 571484 204756 571490 204768
rect 571794 204756 571800 204768
rect 571852 204756 571858 204808
rect 17494 204688 17500 204740
rect 17552 204728 17558 204740
rect 17678 204728 17684 204740
rect 17552 204700 17684 204728
rect 17552 204688 17558 204700
rect 17678 204688 17684 204700
rect 17736 204688 17742 204740
rect 245102 204552 245108 204604
rect 245160 204592 245166 204604
rect 291194 204592 291200 204604
rect 245160 204564 291200 204592
rect 245160 204552 245166 204564
rect 291194 204552 291200 204564
rect 291252 204592 291258 204604
rect 291654 204592 291660 204604
rect 291252 204564 291660 204592
rect 291252 204552 291258 204564
rect 291654 204552 291660 204564
rect 291712 204552 291718 204604
rect 221918 204484 221924 204536
rect 221976 204524 221982 204536
rect 292758 204524 292764 204536
rect 221976 204496 292764 204524
rect 221976 204484 221982 204496
rect 292758 204484 292764 204496
rect 292816 204484 292822 204536
rect 530946 204484 530952 204536
rect 531004 204524 531010 204536
rect 571426 204524 571432 204536
rect 531004 204496 571432 204524
rect 531004 204484 531010 204496
rect 571426 204484 571432 204496
rect 571484 204484 571490 204536
rect 204162 204416 204168 204468
rect 204220 204456 204226 204468
rect 288250 204456 288256 204468
rect 204220 204428 288256 204456
rect 204220 204416 204226 204428
rect 288250 204416 288256 204428
rect 288308 204456 288314 204468
rect 289906 204456 289912 204468
rect 288308 204428 289912 204456
rect 288308 204416 288314 204428
rect 289906 204416 289912 204428
rect 289964 204416 289970 204468
rect 299382 204416 299388 204468
rect 299440 204456 299446 204468
rect 340874 204456 340880 204468
rect 299440 204428 340880 204456
rect 299440 204416 299446 204428
rect 340874 204416 340880 204428
rect 340932 204416 340938 204468
rect 571518 204456 571524 204468
rect 497660 204428 571524 204456
rect 192938 204348 192944 204400
rect 192996 204388 193002 204400
rect 288342 204388 288348 204400
rect 192996 204360 288348 204388
rect 192996 204348 193002 204360
rect 288342 204348 288348 204360
rect 288400 204388 288406 204400
rect 295426 204388 295432 204400
rect 288400 204360 295432 204388
rect 288400 204348 288406 204360
rect 295426 204348 295432 204360
rect 295484 204348 295490 204400
rect 302050 204348 302056 204400
rect 302108 204388 302114 204400
rect 366266 204388 366272 204400
rect 302108 204360 366272 204388
rect 302108 204348 302114 204360
rect 366266 204348 366272 204360
rect 366324 204348 366330 204400
rect 17494 204280 17500 204332
rect 17552 204320 17558 204332
rect 87966 204320 87972 204332
rect 17552 204292 87972 204320
rect 17552 204280 17558 204292
rect 87966 204280 87972 204292
rect 88024 204280 88030 204332
rect 175182 204280 175188 204332
rect 175240 204320 175246 204332
rect 287330 204320 287336 204332
rect 175240 204292 287336 204320
rect 175240 204280 175246 204292
rect 287330 204280 287336 204292
rect 287388 204320 287394 204332
rect 291470 204320 291476 204332
rect 287388 204292 291476 204320
rect 287388 204280 287394 204292
rect 291470 204280 291476 204292
rect 291528 204280 291534 204332
rect 304258 204280 304264 204332
rect 304316 204320 304322 204332
rect 304994 204320 305000 204332
rect 304316 204292 305000 204320
rect 304316 204280 304322 204292
rect 304994 204280 305000 204292
rect 305052 204320 305058 204332
rect 391474 204320 391480 204332
rect 305052 204292 391480 204320
rect 305052 204280 305058 204292
rect 391474 204280 391480 204292
rect 391532 204280 391538 204332
rect 3510 204212 3516 204264
rect 3568 204252 3574 204264
rect 30006 204252 30012 204264
rect 3568 204224 30012 204252
rect 3568 204212 3574 204224
rect 30006 204212 30012 204224
rect 30064 204212 30070 204264
rect 33134 204212 33140 204264
rect 33192 204252 33198 204264
rect 35986 204252 35992 204264
rect 33192 204224 35992 204252
rect 33192 204212 33198 204224
rect 35986 204212 35992 204224
rect 36044 204212 36050 204264
rect 129182 204212 129188 204264
rect 129240 204252 129246 204264
rect 134978 204252 134984 204264
rect 129240 204224 134984 204252
rect 129240 204212 129246 204224
rect 134978 204212 134984 204224
rect 135036 204212 135042 204264
rect 279878 204212 279884 204264
rect 279936 204252 279942 204264
rect 283282 204252 283288 204264
rect 279936 204224 283288 204252
rect 279936 204212 279942 204224
rect 283282 204212 283288 204224
rect 283340 204212 283346 204264
rect 291194 204212 291200 204264
rect 291252 204252 291258 204264
rect 292850 204252 292856 204264
rect 291252 204224 292856 204252
rect 291252 204212 291258 204224
rect 292850 204212 292856 204224
rect 292908 204212 292914 204264
rect 299198 204212 299204 204264
rect 299256 204252 299262 204264
rect 300762 204252 300768 204264
rect 299256 204224 300768 204252
rect 299256 204212 299262 204224
rect 300762 204212 300768 204224
rect 300820 204252 300826 204264
rect 339310 204252 339316 204264
rect 300820 204224 339316 204252
rect 300820 204212 300826 204224
rect 339310 204212 339316 204224
rect 339368 204212 339374 204264
rect 340874 204212 340880 204264
rect 340932 204252 340938 204264
rect 345106 204252 345112 204264
rect 340932 204224 345112 204252
rect 340932 204212 340938 204224
rect 345106 204212 345112 204224
rect 345164 204212 345170 204264
rect 366266 204212 366272 204264
rect 366324 204252 366330 204264
rect 368290 204252 368296 204264
rect 366324 204224 368296 204252
rect 366324 204212 366330 204224
rect 368290 204212 368296 204224
rect 368348 204212 368354 204264
rect 408862 204212 408868 204264
rect 408920 204252 408926 204264
rect 414658 204252 414664 204264
rect 408920 204224 414664 204252
rect 408920 204212 408926 204224
rect 414658 204212 414664 204224
rect 414716 204212 414722 204264
rect 495802 204212 495808 204264
rect 495860 204252 495866 204264
rect 497660 204252 497688 204428
rect 571518 204416 571524 204428
rect 571576 204416 571582 204468
rect 513190 204348 513196 204400
rect 513248 204388 513254 204400
rect 568758 204388 568764 204400
rect 513248 204360 568764 204388
rect 513248 204348 513254 204360
rect 568758 204348 568764 204360
rect 568816 204388 568822 204400
rect 572990 204388 572996 204400
rect 568816 204360 572996 204388
rect 568816 204348 568822 204360
rect 572990 204348 572996 204360
rect 573048 204348 573054 204400
rect 507394 204280 507400 204332
rect 507452 204320 507458 204332
rect 567286 204320 567292 204332
rect 507452 204292 567292 204320
rect 507452 204280 507458 204292
rect 567286 204280 567292 204292
rect 567344 204280 567350 204332
rect 495860 204224 497688 204252
rect 495860 204212 495866 204224
rect 542170 204212 542176 204264
rect 542228 204252 542234 204264
rect 570046 204252 570052 204264
rect 542228 204224 570052 204252
rect 542228 204212 542234 204224
rect 570046 204212 570052 204224
rect 570104 204212 570110 204264
rect 24118 204144 24124 204196
rect 24176 204184 24182 204196
rect 24176 204156 24992 204184
rect 24176 204144 24182 204156
rect 24964 204128 24992 204156
rect 25038 204144 25044 204196
rect 25096 204184 25102 204196
rect 105354 204184 105360 204196
rect 25096 204156 105360 204184
rect 25096 204144 25102 204156
rect 105354 204144 105360 204156
rect 105412 204144 105418 204196
rect 227622 204144 227628 204196
rect 227680 204184 227686 204196
rect 288526 204184 288532 204196
rect 227680 204156 288532 204184
rect 227680 204144 227686 204156
rect 288526 204144 288532 204156
rect 288584 204144 288590 204196
rect 300302 204144 300308 204196
rect 300360 204184 300366 204196
rect 333514 204184 333520 204196
rect 300360 204156 333520 204184
rect 300360 204144 300366 204156
rect 333514 204144 333520 204156
rect 333572 204144 333578 204196
rect 426250 204144 426256 204196
rect 426308 204184 426314 204196
rect 495434 204184 495440 204196
rect 426308 204156 495440 204184
rect 426308 204144 426314 204156
rect 495434 204144 495440 204156
rect 495492 204144 495498 204196
rect 524782 204144 524788 204196
rect 524840 204184 524846 204196
rect 572898 204184 572904 204196
rect 524840 204156 572904 204184
rect 524840 204144 524846 204156
rect 572898 204144 572904 204156
rect 572956 204144 572962 204196
rect 3602 204076 3608 204128
rect 3660 204116 3666 204128
rect 24210 204116 24216 204128
rect 3660 204088 24216 204116
rect 3660 204076 3666 204088
rect 24210 204076 24216 204088
rect 24268 204076 24274 204128
rect 24946 204076 24952 204128
rect 25004 204116 25010 204128
rect 111150 204116 111156 204128
rect 25004 204088 111156 204116
rect 25004 204076 25010 204088
rect 111150 204076 111156 204088
rect 111208 204076 111214 204128
rect 239306 204076 239312 204128
rect 239364 204116 239370 204128
rect 239364 204088 287054 204116
rect 239364 204076 239370 204088
rect 16298 204008 16304 204060
rect 16356 204048 16362 204060
rect 99558 204048 99564 204060
rect 16356 204020 99564 204048
rect 16356 204008 16362 204020
rect 99558 204008 99564 204020
rect 99616 204008 99622 204060
rect 268286 204008 268292 204060
rect 268344 204048 268350 204060
rect 280062 204048 280068 204060
rect 268344 204020 280068 204048
rect 268344 204008 268350 204020
rect 280062 204008 280068 204020
rect 280120 204008 280126 204060
rect 287026 204048 287054 204088
rect 291378 204076 291384 204128
rect 291436 204116 291442 204128
rect 291746 204116 291752 204128
rect 291436 204088 291752 204116
rect 291436 204076 291442 204088
rect 291746 204076 291752 204088
rect 291804 204076 291810 204128
rect 299014 204076 299020 204128
rect 299072 204116 299078 204128
rect 327718 204116 327724 204128
rect 299072 204088 327724 204116
rect 299072 204076 299078 204088
rect 327718 204076 327724 204088
rect 327776 204076 327782 204128
rect 536374 204076 536380 204128
rect 536432 204116 536438 204128
rect 568666 204116 568672 204128
rect 536432 204088 568672 204116
rect 536432 204076 536438 204088
rect 568666 204076 568672 204088
rect 568724 204076 568730 204128
rect 292758 204048 292764 204060
rect 287026 204020 292764 204048
rect 292758 204008 292764 204020
rect 292816 204008 292822 204060
rect 302142 204008 302148 204060
rect 302200 204048 302206 204060
rect 321922 204048 321928 204060
rect 302200 204020 321928 204048
rect 302200 204008 302206 204020
rect 321922 204008 321928 204020
rect 321980 204008 321986 204060
rect 432046 204008 432052 204060
rect 432104 204048 432110 204060
rect 540882 204048 540888 204060
rect 432104 204020 540888 204048
rect 432104 204008 432110 204020
rect 540882 204008 540888 204020
rect 540940 204008 540946 204060
rect 547966 204008 547972 204060
rect 548024 204048 548030 204060
rect 569954 204048 569960 204060
rect 548024 204020 569960 204048
rect 548024 204008 548030 204020
rect 569954 204008 569960 204020
rect 570012 204008 570018 204060
rect 19242 203940 19248 203992
rect 19300 203980 19306 203992
rect 93946 203980 93952 203992
rect 19300 203952 93952 203980
rect 19300 203940 19306 203952
rect 93946 203940 93952 203952
rect 94004 203940 94010 203992
rect 216122 203940 216128 203992
rect 216180 203980 216186 203992
rect 291378 203980 291384 203992
rect 216180 203952 291384 203980
rect 216180 203940 216186 203952
rect 291378 203940 291384 203952
rect 291436 203940 291442 203992
rect 300578 203940 300584 203992
rect 300636 203980 300642 203992
rect 316126 203980 316132 203992
rect 300636 203952 316132 203980
rect 300636 203940 300642 203952
rect 316126 203940 316132 203952
rect 316184 203940 316190 203992
rect 559558 203940 559564 203992
rect 559616 203980 559622 203992
rect 571610 203980 571616 203992
rect 559616 203952 571616 203980
rect 559616 203940 559622 203952
rect 571610 203940 571616 203952
rect 571668 203940 571674 203992
rect 21818 203872 21824 203924
rect 21876 203912 21882 203924
rect 58986 203912 58992 203924
rect 21876 203884 58992 203912
rect 21876 203872 21882 203884
rect 58986 203872 58992 203884
rect 59044 203872 59050 203924
rect 24854 203804 24860 203856
rect 24912 203844 24918 203856
rect 25498 203844 25504 203856
rect 24912 203816 25504 203844
rect 24912 203804 24918 203816
rect 25498 203804 25504 203816
rect 25556 203844 25562 203856
rect 140130 203844 140136 203856
rect 25556 203816 140136 203844
rect 25556 203804 25562 203816
rect 140130 203804 140136 203816
rect 140188 203804 140194 203856
rect 17770 203736 17776 203788
rect 17828 203776 17834 203788
rect 25038 203776 25044 203788
rect 17828 203748 25044 203776
rect 17828 203736 17834 203748
rect 25038 203736 25044 203748
rect 25096 203736 25102 203788
rect 285582 203736 285588 203788
rect 285640 203776 285646 203788
rect 295978 203776 295984 203788
rect 285640 203748 295984 203776
rect 285640 203736 285646 203748
rect 295978 203736 295984 203748
rect 296036 203736 296042 203788
rect 274082 203668 274088 203720
rect 274140 203708 274146 203720
rect 300210 203708 300216 203720
rect 274140 203680 300216 203708
rect 274140 203668 274146 203680
rect 300210 203668 300216 203680
rect 300268 203668 300274 203720
rect 233142 203600 233148 203652
rect 233200 203640 233206 203652
rect 291194 203640 291200 203652
rect 233200 203612 291200 203640
rect 233200 203600 233206 203612
rect 291194 203600 291200 203612
rect 291252 203600 291258 203652
rect 300118 203600 300124 203652
rect 300176 203640 300182 203652
rect 408862 203640 408868 203652
rect 300176 203612 408868 203640
rect 300176 203600 300182 203612
rect 408862 203600 408868 203612
rect 408920 203600 408926 203652
rect 565354 203600 565360 203652
rect 565412 203640 565418 203652
rect 572990 203640 572996 203652
rect 565412 203612 572996 203640
rect 565412 203600 565418 203612
rect 572990 203600 572996 203612
rect 573048 203600 573054 203652
rect 134978 203532 134984 203584
rect 135036 203572 135042 203584
rect 289906 203572 289912 203584
rect 135036 203544 289912 203572
rect 135036 203532 135042 203544
rect 289906 203532 289912 203544
rect 289964 203532 289970 203584
rect 297634 203532 297640 203584
rect 297692 203572 297698 203584
rect 478414 203572 478420 203584
rect 297692 203544 478420 203572
rect 297692 203532 297698 203544
rect 478414 203532 478420 203544
rect 478472 203532 478478 203584
rect 553762 203532 553768 203584
rect 553820 203572 553826 203584
rect 571702 203572 571708 203584
rect 553820 203544 571708 203572
rect 553820 203532 553826 203544
rect 571702 203532 571708 203544
rect 571760 203532 571766 203584
rect 471882 202852 471888 202904
rect 471940 202892 471946 202904
rect 472618 202892 472624 202904
rect 471940 202864 472624 202892
rect 471940 202852 471946 202864
rect 472618 202852 472624 202864
rect 472676 202852 472682 202904
rect 17862 202784 17868 202836
rect 17920 202824 17926 202836
rect 19058 202824 19064 202836
rect 17920 202796 19064 202824
rect 17920 202784 17926 202796
rect 19058 202784 19064 202796
rect 19116 202784 19122 202836
rect 20070 202784 20076 202836
rect 20128 202824 20134 202836
rect 22002 202824 22008 202836
rect 20128 202796 22008 202824
rect 20128 202784 20134 202796
rect 22002 202784 22008 202796
rect 22060 202784 22066 202836
rect 23382 202784 23388 202836
rect 23440 202824 23446 202836
rect 70578 202824 70584 202836
rect 23440 202796 70584 202824
rect 23440 202784 23446 202796
rect 70578 202784 70584 202796
rect 70636 202784 70642 202836
rect 250898 202784 250904 202836
rect 250956 202824 250962 202836
rect 291470 202824 291476 202836
rect 250956 202796 291476 202824
rect 250956 202784 250962 202796
rect 291470 202784 291476 202796
rect 291528 202784 291534 202836
rect 292942 202784 292948 202836
rect 293000 202824 293006 202836
rect 293954 202824 293960 202836
rect 293000 202796 293960 202824
rect 293000 202784 293006 202796
rect 293954 202784 293960 202796
rect 294012 202784 294018 202836
rect 310422 202784 310428 202836
rect 310480 202824 310486 202836
rect 426250 202824 426256 202836
rect 310480 202796 426256 202824
rect 310480 202784 310486 202796
rect 426250 202784 426256 202796
rect 426308 202784 426314 202836
rect 20346 202716 20352 202768
rect 20404 202756 20410 202768
rect 64966 202756 64972 202768
rect 20404 202728 64972 202756
rect 20404 202716 20410 202728
rect 64966 202716 64972 202728
rect 65024 202716 65030 202768
rect 256602 202716 256608 202768
rect 256660 202756 256666 202768
rect 287882 202756 287888 202768
rect 256660 202728 287888 202756
rect 256660 202716 256666 202728
rect 287882 202716 287888 202728
rect 287940 202716 287946 202768
rect 20438 202648 20444 202700
rect 20496 202688 20502 202700
rect 47394 202688 47400 202700
rect 20496 202660 47400 202688
rect 20496 202648 20502 202660
rect 47394 202648 47400 202660
rect 47452 202648 47458 202700
rect 22002 202172 22008 202224
rect 22060 202212 22066 202224
rect 53190 202212 53196 202224
rect 22060 202184 53196 202212
rect 22060 202172 22066 202184
rect 53190 202172 53196 202184
rect 53248 202172 53254 202224
rect 19058 202104 19064 202156
rect 19116 202144 19122 202156
rect 76374 202144 76380 202156
rect 19116 202116 76380 202144
rect 19116 202104 19122 202116
rect 76374 202104 76380 202116
rect 76432 202104 76438 202156
rect 262122 202104 262128 202156
rect 262180 202144 262186 202156
rect 292942 202144 292948 202156
rect 262180 202116 292948 202144
rect 262180 202104 262186 202116
rect 292942 202104 292948 202116
rect 293000 202104 293006 202156
rect 303706 202104 303712 202156
rect 303764 202144 303770 202156
rect 432046 202144 432052 202156
rect 303764 202116 432052 202144
rect 303764 202104 303770 202116
rect 432046 202104 432052 202116
rect 432104 202104 432110 202156
rect 181438 201424 181444 201476
rect 181496 201464 181502 201476
rect 292574 201464 292580 201476
rect 181496 201436 292580 201464
rect 181496 201424 181502 201436
rect 292574 201424 292580 201436
rect 292632 201424 292638 201476
rect 303522 201424 303528 201476
rect 303580 201464 303586 201476
rect 350902 201464 350908 201476
rect 303580 201436 350908 201464
rect 303580 201424 303586 201436
rect 350902 201424 350908 201436
rect 350960 201424 350966 201476
rect 501598 201424 501604 201476
rect 501656 201464 501662 201476
rect 574186 201464 574192 201476
rect 501656 201436 574192 201464
rect 501656 201424 501662 201436
rect 574186 201424 574192 201436
rect 574244 201464 574250 201476
rect 574462 201464 574468 201476
rect 574244 201436 574468 201464
rect 574244 201424 574250 201436
rect 574462 201424 574468 201436
rect 574520 201424 574526 201476
rect 574278 201356 574284 201408
rect 574336 201396 574342 201408
rect 575658 201396 575664 201408
rect 574336 201368 575664 201396
rect 574336 201356 574342 201368
rect 575658 201356 575664 201368
rect 575716 201356 575722 201408
rect 490006 200744 490012 200796
rect 490064 200784 490070 200796
rect 574278 200784 574284 200796
rect 490064 200756 574284 200784
rect 490064 200744 490070 200756
rect 574278 200744 574284 200756
rect 574336 200744 574342 200796
rect 19150 199384 19156 199436
rect 19208 199424 19214 199436
rect 22094 199424 22100 199436
rect 19208 199396 22100 199424
rect 19208 199384 19214 199396
rect 22094 199384 22100 199396
rect 22152 199424 22158 199436
rect 122742 199424 122748 199436
rect 22152 199396 122748 199424
rect 22152 199384 22158 199396
rect 122742 199384 122748 199396
rect 122800 199384 122806 199436
rect 162854 188980 162860 189032
rect 162912 189020 162918 189032
rect 296714 189020 296720 189032
rect 162912 188992 296720 189020
rect 162912 188980 162918 188992
rect 296714 188980 296720 188992
rect 296772 188980 296778 189032
rect 298554 188980 298560 189032
rect 298612 189020 298618 189032
rect 396074 189020 396080 189032
rect 298612 188992 396080 189020
rect 298612 188980 298618 188992
rect 396074 188980 396080 188992
rect 396132 188980 396138 189032
rect 437474 188980 437480 189032
rect 437532 189020 437538 189032
rect 575566 189020 575572 189032
rect 437532 188992 575572 189020
rect 437532 188980 437538 188992
rect 575566 188980 575572 188992
rect 575624 188980 575630 189032
rect 168374 188912 168380 188964
rect 168432 188952 168438 188964
rect 276658 188952 276664 188964
rect 168432 188924 276664 188952
rect 168432 188912 168438 188924
rect 276658 188912 276664 188924
rect 276716 188912 276722 188964
rect 296438 188912 296444 188964
rect 296496 188952 296502 188964
rect 298094 188952 298100 188964
rect 296496 188924 298100 188952
rect 296496 188912 296502 188924
rect 298094 188912 298100 188924
rect 298152 188952 298158 188964
rect 385034 188952 385040 188964
rect 298152 188924 385040 188952
rect 298152 188912 298158 188924
rect 385034 188912 385040 188924
rect 385092 188912 385098 188964
rect 442902 188912 442908 188964
rect 442960 188952 442966 188964
rect 576854 188952 576860 188964
rect 442960 188924 576860 188952
rect 442960 188912 442966 188924
rect 576854 188912 576860 188924
rect 576912 188952 576918 188964
rect 577130 188952 577136 188964
rect 576912 188924 577136 188952
rect 576912 188912 576918 188924
rect 577130 188912 577136 188924
rect 577188 188912 577194 188964
rect 186314 188844 186320 188896
rect 186372 188884 186378 188896
rect 289170 188884 289176 188896
rect 186372 188856 289176 188884
rect 186372 188844 186378 188856
rect 289170 188844 289176 188856
rect 289228 188844 289234 188896
rect 460934 188844 460940 188896
rect 460992 188884 460998 188896
rect 574370 188884 574376 188896
rect 460992 188856 574376 188884
rect 460992 188844 460998 188856
rect 574370 188844 574376 188856
rect 574428 188844 574434 188896
rect 454034 188776 454040 188828
rect 454092 188816 454098 188828
rect 560202 188816 560208 188828
rect 454092 188788 560208 188816
rect 454092 188776 454098 188788
rect 560202 188776 560208 188788
rect 560260 188776 560266 188828
rect 471882 188708 471888 188760
rect 471940 188748 471946 188760
rect 574554 188748 574560 188760
rect 471940 188720 574560 188748
rect 471940 188708 471946 188720
rect 574554 188708 574560 188720
rect 574612 188708 574618 188760
rect 483014 188640 483020 188692
rect 483072 188680 483078 188692
rect 568850 188680 568856 188692
rect 483072 188652 568856 188680
rect 483072 188640 483078 188652
rect 568850 188640 568856 188652
rect 568908 188640 568914 188692
rect 575566 188572 575572 188624
rect 575624 188612 575630 188624
rect 576854 188612 576860 188624
rect 575624 188584 576860 188612
rect 575624 188572 575630 188584
rect 576854 188572 576860 188584
rect 576912 188572 576918 188624
rect 103974 188368 103980 188420
rect 104032 188408 104038 188420
rect 162854 188408 162860 188420
rect 104032 188380 162860 188408
rect 104032 188368 104038 188380
rect 162854 188368 162860 188380
rect 162912 188368 162918 188420
rect 296254 188368 296260 188420
rect 296312 188408 296318 188420
rect 298738 188408 298744 188420
rect 296312 188380 298744 188408
rect 296312 188368 296318 188380
rect 298738 188368 298744 188380
rect 298796 188408 298802 188420
rect 379514 188408 379520 188420
rect 298796 188380 379520 188408
rect 298796 188368 298802 188380
rect 379514 188368 379520 188380
rect 379572 188368 379578 188420
rect 560202 188368 560208 188420
rect 560260 188408 560266 188420
rect 577038 188408 577044 188420
rect 560260 188380 577044 188408
rect 560260 188368 560266 188380
rect 577038 188368 577044 188380
rect 577096 188368 577102 188420
rect 14918 188300 14924 188352
rect 14976 188340 14982 188352
rect 181438 188340 181444 188352
rect 14976 188312 181444 188340
rect 14976 188300 14982 188312
rect 181438 188300 181444 188312
rect 181496 188300 181502 188352
rect 307018 188300 307024 188352
rect 307076 188340 307082 188352
rect 308030 188340 308036 188352
rect 307076 188312 308036 188340
rect 307076 188300 307082 188312
rect 308030 188300 308036 188312
rect 308088 188340 308094 188352
rect 402974 188340 402980 188352
rect 308088 188312 402980 188340
rect 308088 188300 308094 188312
rect 402974 188300 402980 188312
rect 403032 188300 403038 188352
rect 448514 188300 448520 188352
rect 448572 188340 448578 188352
rect 575658 188340 575664 188352
rect 448572 188312 575664 188340
rect 448572 188300 448578 188312
rect 575658 188300 575664 188312
rect 575716 188340 575722 188352
rect 576946 188340 576952 188352
rect 575716 188312 576952 188340
rect 575716 188300 575722 188312
rect 576946 188300 576952 188312
rect 577004 188300 577010 188352
rect 574278 187892 574284 187944
rect 574336 187932 574342 187944
rect 574554 187932 574560 187944
rect 574336 187904 574560 187932
rect 574336 187892 574342 187904
rect 574554 187892 574560 187904
rect 574612 187892 574618 187944
rect 568850 187688 568856 187740
rect 568908 187728 568914 187740
rect 570138 187728 570144 187740
rect 568908 187700 570144 187728
rect 568908 187688 568914 187700
rect 570138 187688 570144 187700
rect 570196 187688 570202 187740
rect 574370 187688 574376 187740
rect 574428 187728 574434 187740
rect 575750 187728 575756 187740
rect 574428 187700 575756 187728
rect 574428 187688 574434 187700
rect 575750 187688 575756 187700
rect 575808 187688 575814 187740
rect 300762 187620 300768 187672
rect 300820 187660 300826 187672
rect 361574 187660 361580 187672
rect 300820 187632 361580 187660
rect 300820 187620 300826 187632
rect 361574 187620 361580 187632
rect 361632 187620 361638 187672
rect 299290 187552 299296 187604
rect 299348 187592 299354 187604
rect 356054 187592 356060 187604
rect 299348 187564 356060 187592
rect 299348 187552 299354 187564
rect 356054 187552 356060 187564
rect 356112 187552 356118 187604
rect 13630 187076 13636 187128
rect 13688 187116 13694 187128
rect 25498 187116 25504 187128
rect 13688 187088 25504 187116
rect 13688 187076 13694 187088
rect 25498 187076 25504 187088
rect 25556 187076 25562 187128
rect 15010 187008 15016 187060
rect 15068 187048 15074 187060
rect 103974 187048 103980 187060
rect 15068 187020 103980 187048
rect 15068 187008 15074 187020
rect 103974 187008 103980 187020
rect 104032 187008 104038 187060
rect 296622 187008 296628 187060
rect 296680 187048 296686 187060
rect 304258 187048 304264 187060
rect 296680 187020 304264 187048
rect 296680 187008 296686 187020
rect 304258 187008 304264 187020
rect 304316 187008 304322 187060
rect 13538 186940 13544 186992
rect 13596 186980 13602 186992
rect 186314 186980 186320 186992
rect 13596 186952 186320 186980
rect 13596 186940 13602 186952
rect 186314 186940 186320 186952
rect 186372 186940 186378 186992
rect 298002 186940 298008 186992
rect 298060 186980 298066 186992
rect 308030 186980 308036 186992
rect 298060 186952 308036 186980
rect 298060 186940 298066 186952
rect 308030 186940 308036 186952
rect 308088 186940 308094 186992
rect 419534 186940 419540 186992
rect 419592 186980 419598 186992
rect 578234 186980 578240 186992
rect 419592 186952 578240 186980
rect 419592 186940 419598 186952
rect 578234 186940 578240 186952
rect 578292 186940 578298 186992
rect 288250 186872 288256 186924
rect 288308 186912 288314 186924
rect 292850 186912 292856 186924
rect 288308 186884 292856 186912
rect 288308 186872 288314 186884
rect 292850 186872 292856 186884
rect 292908 186872 292914 186924
rect 17678 186396 17684 186448
rect 17736 186436 17742 186448
rect 24118 186436 24124 186448
rect 17736 186408 24124 186436
rect 17736 186396 17742 186408
rect 24118 186396 24124 186408
rect 24176 186396 24182 186448
rect 19150 186328 19156 186380
rect 19208 186368 19214 186380
rect 22094 186368 22100 186380
rect 19208 186340 22100 186368
rect 19208 186328 19214 186340
rect 22094 186328 22100 186340
rect 22152 186328 22158 186380
rect 288342 186328 288348 186380
rect 288400 186368 288406 186380
rect 294046 186368 294052 186380
rect 288400 186340 294052 186368
rect 288400 186328 288406 186340
rect 294046 186328 294052 186340
rect 294104 186328 294110 186380
rect 276658 185852 276664 185904
rect 276716 185892 276722 185904
rect 291562 185892 291568 185904
rect 276716 185864 291568 185892
rect 276716 185852 276722 185864
rect 291562 185852 291568 185864
rect 291620 185852 291626 185904
rect 2774 149472 2780 149524
rect 2832 149512 2838 149524
rect 5166 149512 5172 149524
rect 2832 149484 5172 149512
rect 2832 149472 2838 149484
rect 5166 149472 5172 149484
rect 5224 149472 5230 149524
rect 3326 136688 3332 136740
rect 3384 136728 3390 136740
rect 8938 136728 8944 136740
rect 3384 136700 8944 136728
rect 3384 136688 3390 136700
rect 8938 136688 8944 136700
rect 8996 136688 9002 136740
rect 302142 78344 302148 78396
rect 302200 78384 302206 78396
rect 313274 78384 313280 78396
rect 302200 78356 313280 78384
rect 302200 78344 302206 78356
rect 313274 78344 313280 78356
rect 313332 78344 313338 78396
rect 300578 78276 300584 78328
rect 300636 78316 300642 78328
rect 315942 78316 315948 78328
rect 300636 78288 315948 78316
rect 300636 78276 300642 78288
rect 315942 78276 315948 78288
rect 316000 78276 316006 78328
rect 299106 78208 299112 78260
rect 299164 78248 299170 78260
rect 324314 78248 324320 78260
rect 299164 78220 324320 78248
rect 299164 78208 299170 78220
rect 324314 78208 324320 78220
rect 324372 78208 324378 78260
rect 471974 78208 471980 78260
rect 472032 78248 472038 78260
rect 472986 78248 472992 78260
rect 472032 78220 472992 78248
rect 472032 78208 472038 78220
rect 472986 78208 472992 78220
rect 473044 78248 473050 78260
rect 574278 78248 574284 78260
rect 473044 78220 574284 78248
rect 473044 78208 473050 78220
rect 574278 78208 574284 78220
rect 574336 78208 574342 78260
rect 14918 78140 14924 78192
rect 14976 78180 14982 78192
rect 82814 78180 82820 78192
rect 14976 78152 82820 78180
rect 14976 78140 14982 78152
rect 82814 78140 82820 78152
rect 82872 78140 82878 78192
rect 300486 78140 300492 78192
rect 300544 78180 300550 78192
rect 328454 78180 328460 78192
rect 300544 78152 328460 78180
rect 300544 78140 300550 78152
rect 328454 78140 328460 78152
rect 328512 78180 328518 78192
rect 333238 78180 333244 78192
rect 328512 78152 333244 78180
rect 328512 78140 328518 78152
rect 333238 78140 333244 78152
rect 333296 78140 333302 78192
rect 454034 78140 454040 78192
rect 454092 78180 454098 78192
rect 455322 78180 455328 78192
rect 454092 78152 455328 78180
rect 454092 78140 454098 78152
rect 455322 78140 455328 78152
rect 455380 78180 455386 78192
rect 577038 78180 577044 78192
rect 455380 78152 577044 78180
rect 455380 78140 455386 78152
rect 577038 78140 577044 78152
rect 577096 78140 577102 78192
rect 17678 78072 17684 78124
rect 17736 78112 17742 78124
rect 111150 78112 111156 78124
rect 17736 78084 111156 78112
rect 17736 78072 17742 78084
rect 111150 78072 111156 78084
rect 111208 78072 111214 78124
rect 278774 78072 278780 78124
rect 278832 78112 278838 78124
rect 279878 78112 279884 78124
rect 278832 78084 279884 78112
rect 278832 78072 278838 78084
rect 279878 78072 279884 78084
rect 279936 78112 279942 78124
rect 293126 78112 293132 78124
rect 279936 78084 293132 78112
rect 279936 78072 279942 78084
rect 293126 78072 293132 78084
rect 293184 78072 293190 78124
rect 300210 78072 300216 78124
rect 300268 78112 300274 78124
rect 365714 78112 365720 78124
rect 300268 78084 365720 78112
rect 300268 78072 300274 78084
rect 365714 78072 365720 78084
rect 365772 78072 365778 78124
rect 449802 78072 449808 78124
rect 449860 78112 449866 78124
rect 575658 78112 575664 78124
rect 449860 78084 575664 78112
rect 449860 78072 449866 78084
rect 575658 78072 575664 78084
rect 575716 78072 575722 78124
rect 13722 78004 13728 78056
rect 13780 78044 13786 78056
rect 144914 78044 144920 78056
rect 13780 78016 144920 78044
rect 13780 78004 13786 78016
rect 144914 78004 144920 78016
rect 144972 78004 144978 78056
rect 264974 78004 264980 78056
rect 265032 78044 265038 78056
rect 289078 78044 289084 78056
rect 265032 78016 289084 78044
rect 265032 78004 265038 78016
rect 289078 78004 289084 78016
rect 289136 78004 289142 78056
rect 290550 78004 290556 78056
rect 290608 78044 290614 78056
rect 385034 78044 385040 78056
rect 290608 78016 385040 78044
rect 290608 78004 290614 78016
rect 385034 78004 385040 78016
rect 385092 78004 385098 78056
rect 420730 78004 420736 78056
rect 420788 78044 420794 78056
rect 578234 78044 578240 78056
rect 420788 78016 578240 78044
rect 420788 78004 420794 78016
rect 578234 78004 578240 78016
rect 578292 78004 578298 78056
rect 14734 77936 14740 77988
rect 14792 77976 14798 77988
rect 151906 77976 151912 77988
rect 14792 77948 151912 77976
rect 14792 77936 14798 77948
rect 151906 77936 151912 77948
rect 151964 77936 151970 77988
rect 269114 77936 269120 77988
rect 269172 77976 269178 77988
rect 300118 77976 300124 77988
rect 269172 77948 300124 77976
rect 269172 77936 269178 77948
rect 300118 77936 300124 77948
rect 300176 77936 300182 77988
rect 310422 77936 310428 77988
rect 310480 77976 310486 77988
rect 580442 77976 580448 77988
rect 310480 77948 580448 77976
rect 310480 77936 310486 77948
rect 580442 77936 580448 77948
rect 580500 77936 580506 77988
rect 144914 77256 144920 77308
rect 144972 77296 144978 77308
rect 145926 77296 145932 77308
rect 144972 77268 145932 77296
rect 144972 77256 144978 77268
rect 145926 77256 145932 77268
rect 145984 77256 145990 77308
rect 419534 77256 419540 77308
rect 419592 77296 419598 77308
rect 420270 77296 420276 77308
rect 419592 77268 420276 77296
rect 419592 77256 419598 77268
rect 420270 77256 420276 77268
rect 420328 77256 420334 77308
rect 448514 77256 448520 77308
rect 448572 77296 448578 77308
rect 449250 77296 449256 77308
rect 448572 77268 449256 77296
rect 448572 77256 448578 77268
rect 449250 77256 449256 77268
rect 449308 77256 449314 77308
rect 75914 77052 75920 77104
rect 75972 77092 75978 77104
rect 76696 77092 76702 77104
rect 75972 77064 76702 77092
rect 75972 77052 75978 77064
rect 76696 77052 76702 77064
rect 76754 77052 76760 77104
rect 295242 76848 295248 76900
rect 295300 76888 295306 76900
rect 398834 76888 398840 76900
rect 295300 76860 398840 76888
rect 295300 76848 295306 76860
rect 398834 76848 398840 76860
rect 398892 76848 398898 76900
rect 390554 76780 390560 76832
rect 390612 76820 390618 76832
rect 568942 76820 568948 76832
rect 390612 76792 568948 76820
rect 390612 76780 390618 76792
rect 568942 76780 568948 76792
rect 569000 76780 569006 76832
rect 393314 76712 393320 76764
rect 393372 76752 393378 76764
rect 571334 76752 571340 76764
rect 393372 76724 571340 76752
rect 393372 76712 393378 76724
rect 571334 76712 571340 76724
rect 571392 76712 571398 76764
rect 295978 76644 295984 76696
rect 296036 76684 296042 76696
rect 382274 76684 382280 76696
rect 296036 76656 382280 76684
rect 296036 76644 296042 76656
rect 382274 76644 382280 76656
rect 382332 76644 382338 76696
rect 394694 76644 394700 76696
rect 394752 76684 394758 76696
rect 572990 76684 572996 76696
rect 394752 76656 572996 76684
rect 394752 76644 394758 76656
rect 572990 76644 572996 76656
rect 573048 76644 573054 76696
rect 266354 76576 266360 76628
rect 266412 76616 266418 76628
rect 290458 76616 290464 76628
rect 266412 76588 290464 76616
rect 266412 76576 266418 76588
rect 290458 76576 290464 76588
rect 290516 76576 290522 76628
rect 376754 76576 376760 76628
rect 376812 76616 376818 76628
rect 572806 76616 572812 76628
rect 376812 76588 572812 76616
rect 376812 76576 376818 76588
rect 572806 76576 572812 76588
rect 572864 76576 572870 76628
rect 13538 76508 13544 76560
rect 13596 76548 13602 76560
rect 183462 76548 183468 76560
rect 13596 76520 183468 76548
rect 13596 76508 13602 76520
rect 183462 76508 183468 76520
rect 183520 76508 183526 76560
rect 252554 76508 252560 76560
rect 252612 76548 252618 76560
rect 297634 76548 297640 76560
rect 252612 76520 297640 76548
rect 252612 76508 252618 76520
rect 297634 76508 297640 76520
rect 297692 76508 297698 76560
rect 299198 76508 299204 76560
rect 299256 76548 299262 76560
rect 333238 76548 333244 76560
rect 299256 76520 333244 76548
rect 299256 76508 299262 76520
rect 333238 76508 333244 76520
rect 333296 76508 333302 76560
rect 372614 76508 372620 76560
rect 372672 76548 372678 76560
rect 572714 76548 572720 76560
rect 372672 76520 572720 76548
rect 372672 76508 372678 76520
rect 572714 76508 572720 76520
rect 572772 76508 572778 76560
rect 19058 76032 19064 76084
rect 19116 76072 19122 76084
rect 75914 76072 75920 76084
rect 19116 76044 75920 76072
rect 19116 76032 19122 76044
rect 75914 76032 75920 76044
rect 75972 76032 75978 76084
rect 20254 75964 20260 76016
rect 20312 76004 20318 76016
rect 82170 76004 82176 76016
rect 20312 75976 82176 76004
rect 20312 75964 20318 75976
rect 82170 75964 82176 75976
rect 82228 76004 82234 76016
rect 82538 76004 82544 76016
rect 82228 75976 82544 76004
rect 82228 75964 82234 75976
rect 82538 75964 82544 75976
rect 82596 75964 82602 76016
rect 15010 75896 15016 75948
rect 15068 75936 15074 75948
rect 163682 75936 163688 75948
rect 15068 75908 163688 75936
rect 15068 75896 15074 75908
rect 163682 75896 163688 75908
rect 163740 75896 163746 75948
rect 4798 75828 4804 75880
rect 4856 75868 4862 75880
rect 30006 75868 30012 75880
rect 4856 75840 30012 75868
rect 4856 75828 4862 75840
rect 30006 75828 30012 75840
rect 30064 75828 30070 75880
rect 82814 75828 82820 75880
rect 82872 75868 82878 75880
rect 180978 75868 180984 75880
rect 82872 75840 180984 75868
rect 82872 75828 82878 75840
rect 180978 75828 180984 75840
rect 181036 75868 181042 75880
rect 181438 75868 181444 75880
rect 181036 75840 181444 75868
rect 181036 75828 181042 75840
rect 181438 75828 181444 75840
rect 181496 75828 181502 75880
rect 183462 75828 183468 75880
rect 183520 75868 183526 75880
rect 186498 75868 186504 75880
rect 183520 75840 186504 75868
rect 183520 75828 183526 75840
rect 186498 75828 186504 75840
rect 186556 75868 186562 75880
rect 186958 75868 186964 75880
rect 186556 75840 186964 75868
rect 186556 75828 186562 75840
rect 186958 75828 186964 75840
rect 187016 75828 187022 75880
rect 313274 75828 313280 75880
rect 313332 75868 313338 75880
rect 321922 75868 321928 75880
rect 313332 75840 321928 75868
rect 313332 75828 313338 75840
rect 321922 75828 321928 75840
rect 321980 75828 321986 75880
rect 323578 75828 323584 75880
rect 323636 75868 323642 75880
rect 324314 75868 324320 75880
rect 323636 75840 324320 75868
rect 323636 75828 323642 75840
rect 324314 75828 324320 75840
rect 324372 75868 324378 75880
rect 327718 75868 327724 75880
rect 324372 75840 327724 75868
rect 324372 75828 324378 75840
rect 327718 75828 327724 75840
rect 327776 75828 327782 75880
rect 333238 75828 333244 75880
rect 333296 75868 333302 75880
rect 339310 75868 339316 75880
rect 333296 75840 339316 75868
rect 333296 75828 333302 75840
rect 339310 75828 339316 75840
rect 339368 75828 339374 75880
rect 408862 75828 408868 75880
rect 408920 75868 408926 75880
rect 414658 75868 414664 75880
rect 408920 75840 414664 75868
rect 408920 75828 408926 75840
rect 414658 75828 414664 75840
rect 414716 75828 414722 75880
rect 467098 75828 467104 75880
rect 467156 75868 467162 75880
rect 575474 75868 575480 75880
rect 467156 75840 575480 75868
rect 467156 75828 467162 75840
rect 575474 75828 575480 75840
rect 575532 75828 575538 75880
rect 17770 75760 17776 75812
rect 17828 75800 17834 75812
rect 105722 75800 105728 75812
rect 17828 75772 105728 75800
rect 17828 75760 17834 75772
rect 105722 75760 105728 75772
rect 105780 75760 105786 75812
rect 129182 75760 129188 75812
rect 129240 75800 129246 75812
rect 134518 75800 134524 75812
rect 129240 75772 134524 75800
rect 129240 75760 129246 75772
rect 134518 75760 134524 75772
rect 134576 75760 134582 75812
rect 483658 75760 483664 75812
rect 483716 75800 483722 75812
rect 570138 75800 570144 75812
rect 483716 75772 570144 75800
rect 483716 75760 483722 75772
rect 570138 75760 570144 75772
rect 570196 75760 570202 75812
rect 16298 75692 16304 75744
rect 16356 75732 16362 75744
rect 100202 75732 100208 75744
rect 16356 75704 100208 75732
rect 16356 75692 16362 75704
rect 100202 75692 100208 75704
rect 100260 75692 100266 75744
rect 491202 75692 491208 75744
rect 491260 75732 491266 75744
rect 574186 75732 574192 75744
rect 491260 75704 574192 75732
rect 491260 75692 491266 75704
rect 574186 75692 574192 75704
rect 574244 75692 574250 75744
rect 19242 75624 19248 75676
rect 19300 75664 19306 75676
rect 94038 75664 94044 75676
rect 19300 75636 94044 75664
rect 19300 75624 19306 75636
rect 94038 75624 94044 75636
rect 94096 75624 94102 75676
rect 327718 75624 327724 75676
rect 327776 75664 327782 75676
rect 328454 75664 328460 75676
rect 327776 75636 328460 75664
rect 327776 75624 327782 75636
rect 328454 75624 328460 75636
rect 328512 75624 328518 75676
rect 496078 75624 496084 75676
rect 496136 75664 496142 75676
rect 571518 75664 571524 75676
rect 496136 75636 571524 75664
rect 496136 75624 496142 75636
rect 571518 75624 571524 75636
rect 571576 75624 571582 75676
rect 20346 75556 20352 75608
rect 20404 75596 20410 75608
rect 65058 75596 65064 75608
rect 20404 75568 65064 75596
rect 20404 75556 20410 75568
rect 65058 75556 65064 75568
rect 65116 75596 65122 75608
rect 65518 75596 65524 75608
rect 65116 75568 65524 75596
rect 65116 75556 65122 75568
rect 65518 75556 65524 75568
rect 65576 75556 65582 75608
rect 501598 75556 501604 75608
rect 501656 75596 501662 75608
rect 574462 75596 574468 75608
rect 501656 75568 574468 75596
rect 501656 75556 501662 75568
rect 574462 75556 574468 75568
rect 574520 75556 574526 75608
rect 17494 75488 17500 75540
rect 17552 75528 17558 75540
rect 88242 75528 88248 75540
rect 17552 75500 88248 75528
rect 17552 75488 17558 75500
rect 88242 75488 88248 75500
rect 88300 75488 88306 75540
rect 513190 75488 513196 75540
rect 513248 75528 513254 75540
rect 568758 75528 568764 75540
rect 513248 75500 568764 75528
rect 513248 75488 513254 75500
rect 568758 75488 568764 75500
rect 568816 75488 568822 75540
rect 4890 75420 4896 75472
rect 4948 75460 4954 75472
rect 24210 75460 24216 75472
rect 4948 75432 24216 75460
rect 4948 75420 4954 75432
rect 24210 75420 24216 75432
rect 24268 75420 24274 75472
rect 221918 75352 221924 75404
rect 221976 75392 221982 75404
rect 284202 75392 284208 75404
rect 221976 75364 284208 75392
rect 221976 75352 221982 75364
rect 284202 75352 284208 75364
rect 284260 75352 284266 75404
rect 204162 75284 204168 75336
rect 204220 75324 204226 75336
rect 221458 75324 221464 75336
rect 204220 75296 221464 75324
rect 204220 75284 204226 75296
rect 221458 75284 221464 75296
rect 221516 75284 221522 75336
rect 273254 75284 273260 75336
rect 273312 75324 273318 75336
rect 490006 75324 490012 75336
rect 273312 75296 490012 75324
rect 273312 75284 273318 75296
rect 490006 75284 490012 75296
rect 490064 75324 490070 75336
rect 491202 75324 491208 75336
rect 490064 75296 491208 75324
rect 490064 75284 490070 75296
rect 491202 75284 491208 75296
rect 491260 75284 491266 75336
rect 210326 75216 210332 75268
rect 210384 75256 210390 75268
rect 274542 75256 274548 75268
rect 210384 75228 274548 75256
rect 210384 75216 210390 75228
rect 274542 75216 274548 75228
rect 274600 75216 274606 75268
rect 277394 75216 277400 75268
rect 277452 75256 277458 75268
rect 501598 75256 501604 75268
rect 277452 75228 501604 75256
rect 277452 75216 277458 75228
rect 501598 75216 501604 75228
rect 501656 75216 501662 75268
rect 59262 75148 59268 75200
rect 59320 75188 59326 75200
rect 123478 75188 123484 75200
rect 59320 75160 123484 75188
rect 59320 75148 59326 75160
rect 123478 75148 123484 75160
rect 123536 75148 123542 75200
rect 216122 75148 216128 75200
rect 216180 75188 216186 75200
rect 278866 75188 278872 75200
rect 216180 75160 278872 75188
rect 216180 75148 216186 75160
rect 278866 75148 278872 75160
rect 278924 75148 278930 75200
rect 280154 75148 280160 75200
rect 280212 75188 280218 75200
rect 513190 75188 513196 75200
rect 280212 75160 513196 75188
rect 280212 75148 280218 75160
rect 513190 75148 513196 75160
rect 513248 75148 513254 75200
rect 338758 74536 338764 74588
rect 338816 74576 338822 74588
rect 345106 74576 345112 74588
rect 338816 74548 345112 74576
rect 338816 74536 338822 74548
rect 345106 74536 345112 74548
rect 345164 74536 345170 74588
rect 19150 74468 19156 74520
rect 19208 74508 19214 74520
rect 123018 74508 123024 74520
rect 19208 74480 123024 74508
rect 19208 74468 19214 74480
rect 123018 74468 123024 74480
rect 123076 74508 123082 74520
rect 124122 74508 124128 74520
rect 123076 74480 124128 74508
rect 123076 74468 123082 74480
rect 124122 74468 124128 74480
rect 124180 74468 124186 74520
rect 250806 74468 250812 74520
rect 250864 74508 250870 74520
rect 291470 74508 291476 74520
rect 250864 74480 291476 74508
rect 250864 74468 250870 74480
rect 291470 74468 291476 74480
rect 291528 74468 291534 74520
rect 524782 74468 524788 74520
rect 524840 74508 524846 74520
rect 572898 74508 572904 74520
rect 524840 74480 572904 74508
rect 524840 74468 524846 74480
rect 572898 74468 572904 74480
rect 572956 74468 572962 74520
rect 16390 74400 16396 74452
rect 16448 74440 16454 74452
rect 116946 74440 116952 74452
rect 16448 74412 116952 74440
rect 16448 74400 16454 74412
rect 116946 74400 116952 74412
rect 117004 74400 117010 74452
rect 530578 74400 530584 74452
rect 530636 74440 530642 74452
rect 571426 74440 571432 74452
rect 530636 74412 571432 74440
rect 530636 74400 530642 74412
rect 571426 74400 571432 74412
rect 571484 74400 571490 74452
rect 22002 74332 22008 74384
rect 22060 74372 22066 74384
rect 53558 74372 53564 74384
rect 22060 74344 53564 74372
rect 22060 74332 22066 74344
rect 53558 74332 53564 74344
rect 53616 74332 53622 74384
rect 536098 74332 536104 74384
rect 536156 74372 536162 74384
rect 568666 74372 568672 74384
rect 536156 74344 568672 74372
rect 536156 74332 536162 74344
rect 568666 74332 568672 74344
rect 568724 74332 568730 74384
rect 20438 74264 20444 74316
rect 20496 74304 20502 74316
rect 47762 74304 47768 74316
rect 20496 74276 47768 74304
rect 20496 74264 20502 74276
rect 47762 74264 47768 74276
rect 47820 74264 47826 74316
rect 542170 74264 542176 74316
rect 542228 74304 542234 74316
rect 570046 74304 570052 74316
rect 542228 74276 570052 74304
rect 542228 74264 542234 74276
rect 570046 74264 570052 74276
rect 570104 74264 570110 74316
rect 20622 74196 20628 74248
rect 20680 74236 20686 74248
rect 41874 74236 41880 74248
rect 20680 74208 41880 74236
rect 20680 74196 20686 74208
rect 41874 74196 41880 74208
rect 41932 74196 41938 74248
rect 547874 74196 547880 74248
rect 547932 74236 547938 74248
rect 569954 74236 569960 74248
rect 547932 74208 569960 74236
rect 547932 74196 547938 74208
rect 569954 74196 569960 74208
rect 570012 74196 570018 74248
rect 20530 74128 20536 74180
rect 20588 74168 20594 74180
rect 36078 74168 36084 74180
rect 20588 74140 36084 74168
rect 20588 74128 20594 74140
rect 35866 73828 35894 74140
rect 36078 74128 36084 74140
rect 36136 74128 36142 74180
rect 559558 74128 559564 74180
rect 559616 74168 559622 74180
rect 571610 74168 571616 74180
rect 559616 74140 571616 74168
rect 559616 74128 559622 74140
rect 571610 74128 571616 74140
rect 571668 74128 571674 74180
rect 284202 74060 284208 74112
rect 284260 74100 284266 74112
rect 287146 74100 287152 74112
rect 284260 74072 287152 74100
rect 284260 74060 284266 74072
rect 287146 74060 287152 74072
rect 287204 74100 287210 74112
rect 295334 74100 295340 74112
rect 287204 74072 295340 74100
rect 287204 74060 287210 74072
rect 295334 74060 295340 74072
rect 295392 74060 295398 74112
rect 278866 73992 278872 74044
rect 278924 74032 278930 74044
rect 285674 74032 285680 74044
rect 278924 74004 285680 74032
rect 278924 73992 278930 74004
rect 285674 73992 285680 74004
rect 285732 74032 285738 74044
rect 291378 74032 291384 74044
rect 285732 74004 291384 74032
rect 285732 73992 285738 74004
rect 291378 73992 291384 74004
rect 291436 73992 291442 74044
rect 291470 73992 291476 74044
rect 291528 74032 291534 74044
rect 305362 74032 305368 74044
rect 291528 74004 305368 74032
rect 291528 73992 291534 74004
rect 305362 73992 305368 74004
rect 305420 73992 305426 74044
rect 329742 73992 329748 74044
rect 329800 74032 329806 74044
rect 374086 74032 374092 74044
rect 329800 74004 374092 74032
rect 329800 73992 329806 74004
rect 374086 73992 374092 74004
rect 374144 73992 374150 74044
rect 175182 73924 175188 73976
rect 175240 73964 175246 73976
rect 231854 73964 231860 73976
rect 175240 73936 231860 73964
rect 175240 73924 175246 73936
rect 231854 73924 231860 73936
rect 231912 73964 231918 73976
rect 235258 73964 235264 73976
rect 231912 73936 235264 73964
rect 231912 73924 231918 73936
rect 235258 73924 235264 73936
rect 235316 73924 235322 73976
rect 274542 73924 274548 73976
rect 274600 73964 274606 73976
rect 283834 73964 283840 73976
rect 274600 73936 283840 73964
rect 274600 73924 274606 73936
rect 283834 73924 283840 73936
rect 283892 73964 283898 73976
rect 294138 73964 294144 73976
rect 283892 73936 294144 73964
rect 283892 73924 283898 73936
rect 294138 73924 294144 73936
rect 294196 73924 294202 73976
rect 295426 73924 295432 73976
rect 295484 73964 295490 73976
rect 530578 73964 530584 73976
rect 295484 73936 530584 73964
rect 295484 73924 295490 73936
rect 530578 73924 530584 73936
rect 530636 73924 530642 73976
rect 124122 73856 124128 73908
rect 124180 73896 124186 73908
rect 363322 73896 363328 73908
rect 124180 73868 363328 73896
rect 124180 73856 124186 73868
rect 363322 73856 363328 73868
rect 363380 73856 363386 73908
rect 338482 73828 338488 73840
rect 35866 73800 338488 73828
rect 338482 73788 338488 73800
rect 338540 73788 338546 73840
rect 378226 73788 378232 73840
rect 378284 73828 378290 73840
rect 571702 73828 571708 73840
rect 378284 73800 571708 73828
rect 378284 73788 378290 73800
rect 571702 73788 571708 73800
rect 571760 73788 571766 73840
rect 13630 73108 13636 73160
rect 13688 73148 13694 73160
rect 140038 73148 140044 73160
rect 13688 73120 140044 73148
rect 13688 73108 13694 73120
rect 140038 73108 140044 73120
rect 140096 73108 140102 73160
rect 245010 73108 245016 73160
rect 245068 73148 245074 73160
rect 291654 73148 291660 73160
rect 245068 73120 291660 73148
rect 245068 73108 245074 73120
rect 291654 73108 291660 73120
rect 291712 73108 291718 73160
rect 296530 73108 296536 73160
rect 296588 73148 296594 73160
rect 328546 73148 328552 73160
rect 296588 73120 328552 73148
rect 296588 73108 296594 73120
rect 328546 73108 328552 73120
rect 328604 73148 328610 73160
rect 329742 73148 329748 73160
rect 328604 73120 329748 73148
rect 328604 73108 328610 73120
rect 329742 73108 329748 73120
rect 329800 73108 329806 73160
rect 461026 73108 461032 73160
rect 461084 73148 461090 73160
rect 575750 73148 575756 73160
rect 461084 73120 575756 73148
rect 461084 73108 461090 73120
rect 575750 73108 575756 73120
rect 575808 73108 575814 73160
rect 291654 72700 291660 72752
rect 291712 72740 291718 72752
rect 303706 72740 303712 72752
rect 291712 72712 303712 72740
rect 291712 72700 291718 72712
rect 303706 72700 303712 72712
rect 303764 72700 303770 72752
rect 299290 72632 299296 72684
rect 299348 72672 299354 72684
rect 322934 72672 322940 72684
rect 299348 72644 322940 72672
rect 299348 72632 299354 72644
rect 322934 72632 322940 72644
rect 322992 72672 322998 72684
rect 356698 72672 356704 72684
rect 322992 72644 356704 72672
rect 322992 72632 322998 72644
rect 356698 72632 356704 72644
rect 356756 72632 356762 72684
rect 169662 72564 169668 72616
rect 169720 72604 169726 72616
rect 231302 72604 231308 72616
rect 169720 72576 231308 72604
rect 169720 72564 169726 72576
rect 231302 72564 231308 72576
rect 231360 72564 231366 72616
rect 293954 72564 293960 72616
rect 294012 72604 294018 72616
rect 524782 72604 524788 72616
rect 294012 72576 524788 72604
rect 294012 72564 294018 72576
rect 524782 72564 524788 72576
rect 524840 72564 524846 72616
rect 94038 72496 94044 72548
rect 94096 72536 94102 72548
rect 355042 72536 355048 72548
rect 94096 72508 355048 72536
rect 94096 72496 94102 72508
rect 355042 72496 355048 72508
rect 355100 72496 355106 72548
rect 41874 72428 41880 72480
rect 41932 72468 41938 72480
rect 340138 72468 340144 72480
rect 41932 72440 340144 72468
rect 41932 72428 41938 72440
rect 340138 72428 340144 72440
rect 340196 72428 340202 72480
rect 461026 72292 461032 72344
rect 461084 72332 461090 72344
rect 461578 72332 461584 72344
rect 461084 72304 461584 72332
rect 461084 72292 461090 72304
rect 461578 72292 461584 72304
rect 461636 72292 461642 72344
rect 230842 71680 230848 71732
rect 230900 71720 230906 71732
rect 231302 71720 231308 71732
rect 230900 71692 231308 71720
rect 230900 71680 230906 71692
rect 231302 71680 231308 71692
rect 231360 71720 231366 71732
rect 287698 71720 287704 71732
rect 231360 71692 287704 71720
rect 231360 71680 231366 71692
rect 287698 71680 287704 71692
rect 287756 71680 287762 71732
rect 438118 71680 438124 71732
rect 438176 71720 438182 71732
rect 576854 71720 576860 71732
rect 438176 71692 576860 71720
rect 438176 71680 438182 71692
rect 576854 71680 576860 71692
rect 576912 71680 576918 71732
rect 443638 71612 443644 71664
rect 443696 71652 443702 71664
rect 577130 71652 577136 71664
rect 443696 71624 577136 71652
rect 443696 71612 443702 71624
rect 577130 71612 577136 71624
rect 577188 71612 577194 71664
rect 270586 71204 270592 71256
rect 270644 71244 270650 71256
rect 408862 71244 408868 71256
rect 270644 71216 408868 71244
rect 270644 71204 270650 71216
rect 408862 71204 408868 71216
rect 408920 71204 408926 71256
rect 300394 71136 300400 71188
rect 300452 71176 300458 71188
rect 547874 71176 547880 71188
rect 300452 71148 547880 71176
rect 300452 71136 300458 71148
rect 547874 71136 547880 71148
rect 547932 71136 547938 71188
rect 111702 71068 111708 71120
rect 111760 71108 111766 71120
rect 360194 71108 360200 71120
rect 111760 71080 360200 71108
rect 111760 71068 111766 71080
rect 360194 71068 360200 71080
rect 360252 71068 360258 71120
rect 88242 71000 88248 71052
rect 88300 71040 88306 71052
rect 353386 71040 353392 71052
rect 88300 71012 353392 71040
rect 88300 71000 88306 71012
rect 353386 71000 353392 71012
rect 353444 71000 353450 71052
rect 3050 70388 3056 70440
rect 3108 70428 3114 70440
rect 199378 70428 199384 70440
rect 3108 70400 199384 70428
rect 3108 70388 3114 70400
rect 199378 70388 199384 70400
rect 199436 70388 199442 70440
rect 239306 70320 239312 70372
rect 239364 70360 239370 70372
rect 292758 70360 292764 70372
rect 239364 70332 292764 70360
rect 239364 70320 239370 70332
rect 292758 70320 292764 70332
rect 292816 70360 292822 70372
rect 293494 70360 293500 70372
rect 292816 70332 293500 70360
rect 292816 70320 292822 70332
rect 293494 70320 293500 70332
rect 293552 70320 293558 70372
rect 293494 69912 293500 69964
rect 293552 69952 293558 69964
rect 302234 69952 302240 69964
rect 293552 69924 302240 69952
rect 293552 69912 293558 69924
rect 302234 69912 302240 69924
rect 302292 69912 302298 69964
rect 298738 69844 298744 69896
rect 298796 69884 298802 69896
rect 330202 69884 330208 69896
rect 298796 69856 330208 69884
rect 298796 69844 298802 69856
rect 330202 69844 330208 69856
rect 330260 69884 330266 69896
rect 379882 69884 379888 69896
rect 330260 69856 379888 69884
rect 330260 69844 330266 69856
rect 379882 69844 379888 69856
rect 379940 69844 379946 69896
rect 163682 69776 163688 69828
rect 163740 69816 163746 69828
rect 229186 69816 229192 69828
rect 163740 69788 229192 69816
rect 163740 69776 163746 69788
rect 229186 69776 229192 69788
rect 229244 69776 229250 69828
rect 292114 69776 292120 69828
rect 292172 69816 292178 69828
rect 518986 69816 518992 69828
rect 292172 69788 518992 69816
rect 292172 69776 292178 69788
rect 518986 69776 518992 69788
rect 519044 69776 519050 69828
rect 100202 69708 100208 69760
rect 100260 69748 100266 69760
rect 356698 69748 356704 69760
rect 100260 69720 356704 69748
rect 100260 69708 100266 69720
rect 356698 69708 356704 69720
rect 356756 69708 356762 69760
rect 47762 69640 47768 69692
rect 47820 69680 47826 69692
rect 341794 69680 341800 69692
rect 47820 69652 341800 69680
rect 47820 69640 47826 69652
rect 341794 69640 341800 69652
rect 341852 69640 341858 69692
rect 256602 68960 256608 69012
rect 256660 69000 256666 69012
rect 289998 69000 290004 69012
rect 256660 68972 290004 69000
rect 256660 68960 256666 68972
rect 289998 68960 290004 68972
rect 290056 69000 290062 69012
rect 291102 69000 291108 69012
rect 290056 68972 291108 69000
rect 290056 68960 290062 68972
rect 291102 68960 291108 68972
rect 291160 68960 291166 69012
rect 291102 68552 291108 68604
rect 291160 68592 291166 68604
rect 307018 68592 307024 68604
rect 291160 68564 307024 68592
rect 291160 68552 291166 68564
rect 307018 68552 307024 68564
rect 307076 68552 307082 68604
rect 298738 68484 298744 68536
rect 298796 68524 298802 68536
rect 542170 68524 542176 68536
rect 298796 68496 542176 68524
rect 298796 68484 298802 68496
rect 542170 68484 542176 68496
rect 542228 68484 542234 68536
rect 105722 68416 105728 68468
rect 105780 68456 105786 68468
rect 358354 68456 358360 68468
rect 105780 68428 358360 68456
rect 105780 68416 105786 68428
rect 358354 68416 358360 68428
rect 358412 68416 358418 68468
rect 82538 68348 82544 68400
rect 82596 68388 82602 68400
rect 351914 68388 351920 68400
rect 82596 68360 351920 68388
rect 82596 68348 82602 68360
rect 351914 68348 351920 68360
rect 351972 68348 351978 68400
rect 53558 68280 53564 68332
rect 53616 68320 53622 68332
rect 343634 68320 343640 68332
rect 53616 68292 343640 68320
rect 53616 68280 53622 68292
rect 343634 68280 343640 68292
rect 343692 68280 343698 68332
rect 267734 67532 267740 67584
rect 267792 67572 267798 67584
rect 292574 67572 292580 67584
rect 267792 67544 292580 67572
rect 267792 67532 267798 67544
rect 292574 67532 292580 67544
rect 292632 67532 292638 67584
rect 197354 67056 197360 67108
rect 197412 67096 197418 67108
rect 221550 67096 221556 67108
rect 197412 67068 221556 67096
rect 197412 67056 197418 67068
rect 221550 67056 221556 67068
rect 221608 67056 221614 67108
rect 292574 67056 292580 67108
rect 292632 67096 292638 67108
rect 310514 67096 310520 67108
rect 292632 67068 310520 67096
rect 292632 67056 292638 67068
rect 310514 67056 310520 67068
rect 310572 67056 310578 67108
rect 336642 67056 336648 67108
rect 336700 67096 336706 67108
rect 396074 67096 396080 67108
rect 336700 67068 396080 67096
rect 336700 67056 336706 67068
rect 396074 67056 396080 67068
rect 396132 67056 396138 67108
rect 134518 66988 134524 67040
rect 134576 67028 134582 67040
rect 255682 67028 255688 67040
rect 134576 67000 255688 67028
rect 134576 66988 134582 67000
rect 255682 66988 255688 67000
rect 255740 66988 255746 67040
rect 297082 66988 297088 67040
rect 297140 67028 297146 67040
rect 536098 67028 536104 67040
rect 297140 67000 536104 67028
rect 297140 66988 297146 67000
rect 536098 66988 536104 67000
rect 536156 66988 536162 67040
rect 116946 66920 116952 66972
rect 117004 66960 117010 66972
rect 361666 66960 361672 66972
rect 117004 66932 361672 66960
rect 117004 66920 117010 66932
rect 361666 66920 361672 66932
rect 361724 66920 361730 66972
rect 220906 66852 220912 66904
rect 220964 66892 220970 66904
rect 471974 66892 471980 66904
rect 220964 66864 471980 66892
rect 220964 66852 220970 66864
rect 471974 66852 471980 66864
rect 472032 66852 472038 66904
rect 215938 65628 215944 65680
rect 215996 65668 216002 65680
rect 454034 65668 454040 65680
rect 215996 65640 454040 65668
rect 215996 65628 216002 65640
rect 454034 65628 454040 65640
rect 454092 65628 454098 65680
rect 219434 65560 219440 65612
rect 219492 65600 219498 65612
rect 467098 65600 467104 65612
rect 219492 65572 467104 65600
rect 219492 65560 219498 65572
rect 467098 65560 467104 65572
rect 467156 65560 467162 65612
rect 202874 65492 202880 65544
rect 202932 65532 202938 65544
rect 559558 65532 559564 65544
rect 202932 65504 559564 65532
rect 202932 65492 202938 65504
rect 559558 65492 559564 65504
rect 559616 65492 559622 65544
rect 302326 64812 302332 64864
rect 302384 64852 302390 64864
rect 431954 64852 431960 64864
rect 302384 64824 431960 64852
rect 302384 64812 302390 64824
rect 431954 64812 431960 64824
rect 432012 64812 432018 64864
rect 209314 64336 209320 64388
rect 209372 64376 209378 64388
rect 302326 64376 302332 64388
rect 209372 64348 302332 64376
rect 209372 64336 209378 64348
rect 302326 64336 302332 64348
rect 302384 64336 302390 64388
rect 272518 64268 272524 64320
rect 272576 64308 272582 64320
rect 477494 64308 477500 64320
rect 272576 64280 477500 64308
rect 272576 64268 272582 64280
rect 477494 64268 477500 64280
rect 477552 64268 477558 64320
rect 212626 64200 212632 64252
rect 212684 64240 212690 64252
rect 443638 64240 443644 64252
rect 212684 64212 443644 64240
rect 212684 64200 212690 64212
rect 443638 64200 443644 64212
rect 443696 64200 443702 64252
rect 8938 64132 8944 64184
rect 8996 64172 9002 64184
rect 57606 64172 57612 64184
rect 8996 64144 57612 64172
rect 8996 64132 9002 64144
rect 57606 64132 57612 64144
rect 57664 64132 57670 64184
rect 217594 64132 217600 64184
rect 217652 64172 217658 64184
rect 461578 64172 461584 64184
rect 217652 64144 461584 64172
rect 217652 64132 217658 64144
rect 461578 64132 461584 64144
rect 461636 64132 461642 64184
rect 123478 62976 123484 63028
rect 123536 63016 123542 63028
rect 345106 63016 345112 63028
rect 123536 62988 345112 63016
rect 123536 62976 123542 62988
rect 345106 62976 345112 62988
rect 345164 62976 345170 63028
rect 75914 62908 75920 62960
rect 75972 62948 75978 62960
rect 350074 62948 350080 62960
rect 75972 62920 350080 62948
rect 75972 62908 75978 62920
rect 350074 62908 350080 62920
rect 350132 62908 350138 62960
rect 71038 62840 71044 62892
rect 71096 62880 71102 62892
rect 348418 62880 348424 62892
rect 71096 62852 348424 62880
rect 71096 62840 71102 62852
rect 348418 62840 348424 62852
rect 348476 62840 348482 62892
rect 65518 62772 65524 62824
rect 65576 62812 65582 62824
rect 346762 62812 346768 62824
rect 65576 62784 346768 62812
rect 65576 62772 65582 62784
rect 346762 62772 346768 62784
rect 346820 62772 346826 62824
rect 379882 62772 379888 62824
rect 379940 62812 379946 62824
rect 553394 62812 553400 62824
rect 379940 62784 553400 62812
rect 379940 62772 379946 62784
rect 553394 62772 553400 62784
rect 553452 62772 553458 62824
rect 226334 62024 226340 62076
rect 226392 62064 226398 62076
rect 288526 62064 288532 62076
rect 226392 62036 288532 62064
rect 226392 62024 226398 62036
rect 288526 62024 288532 62036
rect 288584 62064 288590 62076
rect 288802 62064 288808 62076
rect 288584 62036 288808 62064
rect 288584 62024 288590 62036
rect 288802 62024 288808 62036
rect 288860 62024 288866 62076
rect 303798 62024 303804 62076
rect 303856 62064 303862 62076
rect 425054 62064 425060 62076
rect 303856 62036 425060 62064
rect 303856 62024 303862 62036
rect 425054 62024 425060 62036
rect 425112 62024 425118 62076
rect 186958 61548 186964 61600
rect 187016 61588 187022 61600
rect 235994 61588 236000 61600
rect 187016 61560 236000 61588
rect 187016 61548 187022 61560
rect 235994 61548 236000 61560
rect 236052 61548 236058 61600
rect 315298 61548 315304 61600
rect 315356 61588 315362 61600
rect 323578 61588 323584 61600
rect 315356 61560 323584 61588
rect 315356 61548 315362 61560
rect 323578 61548 323584 61560
rect 323636 61548 323642 61600
rect 144914 61480 144920 61532
rect 144972 61520 144978 61532
rect 221734 61520 221740 61532
rect 144972 61492 221740 61520
rect 144972 61480 144978 61492
rect 221734 61480 221740 61492
rect 221792 61480 221798 61532
rect 300762 61480 300768 61532
rect 300820 61520 300826 61532
rect 325234 61520 325240 61532
rect 300820 61492 325240 61520
rect 300820 61480 300826 61492
rect 325234 61480 325240 61492
rect 325292 61520 325298 61532
rect 361574 61520 361580 61532
rect 325292 61492 361580 61520
rect 325292 61480 325298 61492
rect 361574 61480 361580 61492
rect 361632 61480 361638 61532
rect 140038 61412 140044 61464
rect 140096 61452 140102 61464
rect 222562 61452 222568 61464
rect 140096 61424 222568 61452
rect 140096 61412 140102 61424
rect 222562 61412 222568 61424
rect 222620 61412 222626 61464
rect 284294 61412 284300 61464
rect 284352 61452 284358 61464
rect 381538 61452 381544 61464
rect 284352 61424 381544 61452
rect 284352 61412 284358 61424
rect 381538 61412 381544 61424
rect 381596 61412 381602 61464
rect 222102 61344 222108 61396
rect 222160 61384 222166 61396
rect 438118 61384 438124 61396
rect 222160 61356 438124 61384
rect 222160 61344 222166 61356
rect 438118 61344 438124 61356
rect 438176 61344 438182 61396
rect 318794 60324 318800 60376
rect 318852 60364 318858 60376
rect 333238 60364 333244 60376
rect 318852 60336 333244 60364
rect 318852 60324 318858 60336
rect 333238 60324 333244 60336
rect 333296 60324 333302 60376
rect 321922 60256 321928 60308
rect 321980 60296 321986 60308
rect 350534 60296 350540 60308
rect 321980 60268 350540 60296
rect 321980 60256 321986 60268
rect 350534 60256 350540 60268
rect 350592 60256 350598 60308
rect 191834 60188 191840 60240
rect 191892 60228 191898 60240
rect 237374 60228 237380 60240
rect 191892 60200 237380 60228
rect 191892 60188 191898 60200
rect 237374 60188 237380 60200
rect 237432 60188 237438 60240
rect 273346 60188 273352 60240
rect 273404 60228 273410 60240
rect 320082 60228 320088 60240
rect 273404 60200 320088 60228
rect 273404 60188 273410 60200
rect 320082 60188 320088 60200
rect 320140 60188 320146 60240
rect 331858 60228 331864 60240
rect 325666 60200 331864 60228
rect 181438 60120 181444 60172
rect 181496 60160 181502 60172
rect 234154 60160 234160 60172
rect 181496 60132 234160 60160
rect 181496 60120 181502 60132
rect 234154 60120 234160 60132
rect 234212 60120 234218 60172
rect 242434 60120 242440 60172
rect 242492 60160 242498 60172
rect 289814 60160 289820 60172
rect 242492 60132 289820 60160
rect 242492 60120 242498 60132
rect 289814 60120 289820 60132
rect 289872 60120 289878 60172
rect 296438 60120 296444 60172
rect 296496 60160 296502 60172
rect 325666 60160 325694 60200
rect 331858 60188 331864 60200
rect 331916 60228 331922 60240
rect 385126 60228 385132 60240
rect 331916 60200 385132 60228
rect 331916 60188 331922 60200
rect 385126 60188 385132 60200
rect 385184 60188 385190 60240
rect 296496 60132 325694 60160
rect 296496 60120 296502 60132
rect 332962 60120 332968 60172
rect 333020 60160 333026 60172
rect 390646 60160 390652 60172
rect 333020 60132 390652 60160
rect 333020 60120 333026 60132
rect 390646 60120 390652 60132
rect 390704 60120 390710 60172
rect 221458 60052 221464 60104
rect 221516 60092 221522 60104
rect 282178 60092 282184 60104
rect 221516 60064 282184 60092
rect 221516 60052 221522 60064
rect 282178 60052 282184 60064
rect 282236 60092 282242 60104
rect 292850 60092 292856 60104
rect 282236 60064 292856 60092
rect 282236 60052 282242 60064
rect 292850 60052 292856 60064
rect 292908 60052 292914 60104
rect 294598 60052 294604 60104
rect 294656 60092 294662 60104
rect 371602 60092 371608 60104
rect 294656 60064 371608 60092
rect 294656 60052 294662 60064
rect 371602 60052 371608 60064
rect 371660 60052 371666 60104
rect 206002 59984 206008 60036
rect 206060 60024 206066 60036
rect 419534 60024 419540 60036
rect 206060 59996 419540 60024
rect 206060 59984 206066 59996
rect 419534 59984 419540 59996
rect 419592 59984 419598 60036
rect 237374 59304 237380 59356
rect 237432 59344 237438 59356
rect 294046 59344 294052 59356
rect 237432 59316 294052 59344
rect 237432 59304 237438 59316
rect 294046 59304 294052 59316
rect 294104 59304 294110 59356
rect 296622 59304 296628 59356
rect 296680 59344 296686 59356
rect 332962 59344 332968 59356
rect 296680 59316 332968 59344
rect 296680 59304 296686 59316
rect 332962 59304 332968 59316
rect 333020 59344 333026 59356
rect 333514 59344 333520 59356
rect 333020 59316 333520 59344
rect 333020 59304 333026 59316
rect 333514 59304 333520 59316
rect 333572 59304 333578 59356
rect 260834 59236 260840 59288
rect 260892 59276 260898 59288
rect 292574 59276 292580 59288
rect 260892 59248 292580 59276
rect 260892 59236 260898 59248
rect 292574 59236 292580 59248
rect 292632 59276 292638 59288
rect 292942 59276 292948 59288
rect 292632 59248 292948 59276
rect 292632 59236 292638 59248
rect 292942 59236 292948 59248
rect 293000 59236 293006 59288
rect 316954 58896 316960 58948
rect 317012 58936 317018 58948
rect 327718 58936 327724 58948
rect 317012 58908 327724 58936
rect 317012 58896 317018 58908
rect 327718 58896 327724 58908
rect 327776 58896 327782 58948
rect 220722 58828 220728 58880
rect 220780 58868 220786 58880
rect 278774 58868 278780 58880
rect 220780 58840 278780 58868
rect 220780 58828 220786 58840
rect 278774 58828 278780 58840
rect 278832 58828 278838 58880
rect 320818 58828 320824 58880
rect 320876 58868 320882 58880
rect 338758 58868 338764 58880
rect 320876 58840 338764 58868
rect 320876 58828 320882 58840
rect 338758 58828 338764 58840
rect 338816 58828 338822 58880
rect 157978 58760 157984 58812
rect 158036 58800 158042 58812
rect 227714 58800 227720 58812
rect 158036 58772 227720 58800
rect 158036 58760 158042 58772
rect 227714 58760 227720 58772
rect 227772 58760 227778 58812
rect 298002 58760 298008 58812
rect 298060 58800 298066 58812
rect 336826 58800 336832 58812
rect 298060 58772 336832 58800
rect 298060 58760 298066 58772
rect 336826 58760 336832 58772
rect 336884 58800 336890 58812
rect 402974 58800 402980 58812
rect 336884 58772 402980 58800
rect 336884 58760 336890 58772
rect 402974 58760 402980 58772
rect 403032 58760 403038 58812
rect 151814 58692 151820 58744
rect 151872 58732 151878 58744
rect 225874 58732 225880 58744
rect 151872 58704 225880 58732
rect 151872 58692 151878 58704
rect 225874 58692 225880 58704
rect 225932 58692 225938 58744
rect 231946 58692 231952 58744
rect 232004 58732 232010 58744
rect 261570 58732 261576 58744
rect 232004 58704 261576 58732
rect 232004 58692 232010 58704
rect 261570 58692 261576 58704
rect 261628 58692 261634 58744
rect 328362 58692 328368 58744
rect 328420 58732 328426 58744
rect 367094 58732 367100 58744
rect 328420 58704 367100 58732
rect 328420 58692 328426 58704
rect 367094 58692 367100 58704
rect 367152 58692 367158 58744
rect 396442 58692 396448 58744
rect 396500 58732 396506 58744
rect 564434 58732 564440 58744
rect 396500 58704 564440 58732
rect 396500 58692 396506 58704
rect 564434 58692 564440 58704
rect 564492 58692 564498 58744
rect 214282 58624 214288 58676
rect 214340 58664 214346 58676
rect 448514 58664 448520 58676
rect 214340 58636 448520 58664
rect 214340 58624 214346 58636
rect 448514 58624 448520 58636
rect 448572 58624 448578 58676
rect 102134 57944 102140 57996
rect 102192 57984 102198 57996
rect 104158 57984 104164 57996
rect 102192 57956 104164 57984
rect 102192 57944 102198 57956
rect 104158 57944 104164 57956
rect 104216 57944 104222 57996
rect 221734 57876 221740 57928
rect 221792 57916 221798 57928
rect 224586 57916 224592 57928
rect 221792 57888 224592 57916
rect 221792 57876 221798 57888
rect 224586 57876 224592 57888
rect 224644 57876 224650 57928
rect 299382 57876 299388 57928
rect 299440 57916 299446 57928
rect 320818 57916 320824 57928
rect 299440 57888 320824 57916
rect 299440 57876 299446 57888
rect 320818 57876 320824 57888
rect 320876 57876 320882 57928
rect 261570 57604 261576 57656
rect 261628 57644 261634 57656
rect 291102 57644 291108 57656
rect 261628 57616 291108 57644
rect 261628 57604 261634 57616
rect 291102 57604 291108 57616
rect 291160 57604 291166 57656
rect 259362 57536 259368 57588
rect 259420 57576 259426 57588
rect 288434 57576 288440 57588
rect 259420 57548 288440 57576
rect 259420 57536 259426 57548
rect 288434 57536 288440 57548
rect 288492 57536 288498 57588
rect 292574 57536 292580 57588
rect 292632 57576 292638 57588
rect 309042 57576 309048 57588
rect 292632 57548 309048 57576
rect 292632 57536 292638 57548
rect 309042 57536 309048 57548
rect 309100 57536 309106 57588
rect 320082 57536 320088 57588
rect 320140 57576 320146 57588
rect 365346 57576 365352 57588
rect 320140 57548 365352 57576
rect 320140 57536 320146 57548
rect 365346 57536 365352 57548
rect 365404 57536 365410 57588
rect 251082 57468 251088 57520
rect 251140 57508 251146 57520
rect 297450 57508 297456 57520
rect 251140 57480 297456 57508
rect 251140 57468 251146 57480
rect 297450 57468 297456 57480
rect 297508 57468 297514 57520
rect 297542 57468 297548 57520
rect 297600 57508 297606 57520
rect 368658 57508 368664 57520
rect 297600 57480 368664 57508
rect 297600 57468 297606 57480
rect 368658 57468 368664 57480
rect 368716 57468 368722 57520
rect 257706 57400 257712 57452
rect 257764 57440 257770 57452
rect 289906 57440 289912 57452
rect 257764 57412 289912 57440
rect 257764 57400 257770 57412
rect 289906 57400 289912 57412
rect 289964 57400 289970 57452
rect 294690 57400 294696 57452
rect 294748 57440 294754 57452
rect 370314 57440 370320 57452
rect 294748 57412 370320 57440
rect 294748 57400 294754 57412
rect 370314 57400 370320 57412
rect 370372 57400 370378 57452
rect 211338 57332 211344 57384
rect 211396 57372 211402 57384
rect 222102 57372 222108 57384
rect 211396 57344 222108 57372
rect 211396 57332 211402 57344
rect 222102 57332 222108 57344
rect 222160 57332 222166 57384
rect 272610 57332 272616 57384
rect 272668 57372 272674 57384
rect 483658 57372 483664 57384
rect 272668 57344 483664 57372
rect 272668 57332 272674 57344
rect 483658 57332 483664 57344
rect 483716 57332 483722 57384
rect 208026 57264 208032 57316
rect 208084 57304 208090 57316
rect 218054 57304 218060 57316
rect 208084 57276 218060 57304
rect 208084 57264 208090 57276
rect 218054 57264 218060 57276
rect 218112 57264 218118 57316
rect 275922 57264 275928 57316
rect 275980 57304 275986 57316
rect 496078 57304 496084 57316
rect 275980 57276 496084 57304
rect 275980 57264 275986 57276
rect 496078 57264 496084 57276
rect 496136 57264 496142 57316
rect 204714 57196 204720 57248
rect 204772 57236 204778 57248
rect 220722 57236 220728 57248
rect 204772 57208 220728 57236
rect 204772 57196 204778 57208
rect 220722 57196 220728 57208
rect 220780 57196 220786 57248
rect 221550 57196 221556 57248
rect 221608 57236 221614 57248
rect 239490 57236 239496 57248
rect 221608 57208 239496 57236
rect 221608 57196 221614 57208
rect 239490 57196 239496 57208
rect 239548 57196 239554 57248
rect 254394 57196 254400 57248
rect 254452 57236 254458 57248
rect 272518 57236 272524 57248
rect 254452 57208 272524 57236
rect 254452 57196 254458 57208
rect 272518 57196 272524 57208
rect 272576 57196 272582 57248
rect 279234 57196 279240 57248
rect 279292 57236 279298 57248
rect 507118 57236 507124 57248
rect 279292 57208 507124 57236
rect 279292 57196 279298 57208
rect 507118 57196 507124 57208
rect 507176 57196 507182 57248
rect 312354 56584 312360 56636
rect 312412 56624 312418 56636
rect 316034 56624 316040 56636
rect 312412 56596 316040 56624
rect 312412 56584 312418 56596
rect 316034 56584 316040 56596
rect 316092 56584 316098 56636
rect 5166 56516 5172 56568
rect 5224 56556 5230 56568
rect 57514 56556 57520 56568
rect 5224 56528 57520 56556
rect 5224 56516 5230 56528
rect 57514 56516 57520 56528
rect 57572 56516 57578 56568
rect 102134 53796 102140 53848
rect 102192 53836 102198 53848
rect 109034 53836 109040 53848
rect 102192 53808 109040 53836
rect 102192 53796 102198 53808
rect 109034 53796 109040 53808
rect 109092 53796 109098 53848
rect 102134 52640 102140 52692
rect 102192 52680 102198 52692
rect 103882 52680 103888 52692
rect 102192 52652 103888 52680
rect 102192 52640 102198 52652
rect 103882 52640 103888 52652
rect 103940 52640 103946 52692
rect 102134 52436 102140 52488
rect 102192 52476 102198 52488
rect 196158 52476 196164 52488
rect 102192 52448 196164 52476
rect 102192 52436 102198 52448
rect 196158 52436 196164 52448
rect 196216 52436 196222 52488
rect 5074 52368 5080 52420
rect 5132 52408 5138 52420
rect 57054 52408 57060 52420
rect 5132 52380 57060 52408
rect 5132 52368 5138 52380
rect 57054 52368 57060 52380
rect 57112 52368 57118 52420
rect 102778 52368 102784 52420
rect 102836 52408 102842 52420
rect 195974 52408 195980 52420
rect 102836 52380 195980 52408
rect 102836 52368 102842 52380
rect 195974 52368 195980 52380
rect 196032 52368 196038 52420
rect 102870 52300 102876 52352
rect 102928 52340 102934 52352
rect 196066 52340 196072 52352
rect 102928 52312 196072 52340
rect 102928 52300 102934 52312
rect 196066 52300 196072 52312
rect 196124 52300 196130 52352
rect 102962 51008 102968 51060
rect 103020 51048 103026 51060
rect 195974 51048 195980 51060
rect 103020 51020 195980 51048
rect 103020 51008 103026 51020
rect 195974 51008 195980 51020
rect 196032 51008 196038 51060
rect 102134 49784 102140 49836
rect 102192 49824 102198 49836
rect 104434 49824 104440 49836
rect 102192 49796 104440 49824
rect 102192 49784 102198 49796
rect 104434 49784 104440 49796
rect 104492 49784 104498 49836
rect 102594 49648 102600 49700
rect 102652 49688 102658 49700
rect 196066 49688 196072 49700
rect 102652 49660 196072 49688
rect 102652 49648 102658 49660
rect 196066 49648 196072 49660
rect 196124 49648 196130 49700
rect 104158 49580 104164 49632
rect 104216 49620 104222 49632
rect 195974 49620 195980 49632
rect 104216 49592 195980 49620
rect 104216 49580 104222 49592
rect 195974 49580 195980 49592
rect 196032 49580 196038 49632
rect 102134 48832 102140 48884
rect 102192 48872 102198 48884
rect 104342 48872 104348 48884
rect 102192 48844 104348 48872
rect 102192 48832 102198 48844
rect 104342 48832 104348 48844
rect 104400 48832 104406 48884
rect 103054 48220 103060 48272
rect 103112 48260 103118 48272
rect 195974 48260 195980 48272
rect 103112 48232 195980 48260
rect 103112 48220 103118 48232
rect 195974 48220 195980 48232
rect 196032 48220 196038 48272
rect 109034 48152 109040 48204
rect 109092 48192 109098 48204
rect 196066 48192 196072 48204
rect 109092 48164 196072 48192
rect 109092 48152 109098 48164
rect 196066 48152 196072 48164
rect 196124 48152 196130 48204
rect 6178 46860 6184 46912
rect 6236 46900 6242 46912
rect 57514 46900 57520 46912
rect 6236 46872 57520 46900
rect 6236 46860 6242 46872
rect 57514 46860 57520 46872
rect 57572 46860 57578 46912
rect 103882 46860 103888 46912
rect 103940 46900 103946 46912
rect 195974 46900 195980 46912
rect 103940 46872 195980 46900
rect 103940 46860 103946 46872
rect 195974 46860 195980 46872
rect 196032 46860 196038 46912
rect 103238 45500 103244 45552
rect 103296 45540 103302 45552
rect 195974 45540 195980 45552
rect 103296 45512 195980 45540
rect 103296 45500 103302 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 104434 44820 104440 44872
rect 104492 44860 104498 44872
rect 196066 44860 196072 44872
rect 104492 44832 196072 44860
rect 104492 44820 104498 44832
rect 196066 44820 196072 44832
rect 196124 44820 196130 44872
rect 3326 44140 3332 44192
rect 3384 44180 3390 44192
rect 59998 44180 60004 44192
rect 3384 44152 60004 44180
rect 3384 44140 3390 44152
rect 59998 44140 60004 44152
rect 60056 44140 60062 44192
rect 104342 44072 104348 44124
rect 104400 44112 104406 44124
rect 195974 44112 195980 44124
rect 104400 44084 195980 44112
rect 104400 44072 104406 44084
rect 195974 44072 195980 44084
rect 196032 44072 196038 44124
rect 3510 42712 3516 42764
rect 3568 42752 3574 42764
rect 57146 42752 57152 42764
rect 3568 42724 57152 42752
rect 3568 42712 3574 42724
rect 57146 42712 57152 42724
rect 57204 42712 57210 42764
rect 102962 42712 102968 42764
rect 103020 42752 103026 42764
rect 195974 42752 195980 42764
rect 103020 42724 195980 42752
rect 103020 42712 103026 42724
rect 195974 42712 195980 42724
rect 196032 42712 196038 42764
rect 102594 42644 102600 42696
rect 102652 42684 102658 42696
rect 196066 42684 196072 42696
rect 102652 42656 196072 42684
rect 102652 42644 102658 42656
rect 196066 42644 196072 42656
rect 196124 42644 196130 42696
rect 102870 41352 102876 41404
rect 102928 41392 102934 41404
rect 195974 41392 195980 41404
rect 102928 41364 195980 41392
rect 102928 41352 102934 41364
rect 195974 41352 195980 41364
rect 196032 41352 196038 41404
rect 102134 40672 102140 40724
rect 102192 40712 102198 40724
rect 196158 40712 196164 40724
rect 102192 40684 196164 40712
rect 102192 40672 102198 40684
rect 196158 40672 196164 40684
rect 196216 40672 196222 40724
rect 102318 39992 102324 40044
rect 102376 40032 102382 40044
rect 196066 40032 196072 40044
rect 102376 40004 196072 40032
rect 102376 39992 102382 40004
rect 196066 39992 196072 40004
rect 196124 39992 196130 40044
rect 103514 39924 103520 39976
rect 103572 39964 103578 39976
rect 195974 39964 195980 39976
rect 103572 39936 195980 39964
rect 103572 39924 103578 39936
rect 195974 39924 195980 39936
rect 196032 39924 196038 39976
rect 102226 38564 102232 38616
rect 102284 38604 102290 38616
rect 195974 38604 195980 38616
rect 102284 38576 195980 38604
rect 102284 38564 102290 38576
rect 195974 38564 195980 38576
rect 196032 38564 196038 38616
rect 6270 37204 6276 37256
rect 6328 37244 6334 37256
rect 57054 37244 57060 37256
rect 6328 37216 57060 37244
rect 6328 37204 6334 37216
rect 57054 37204 57060 37216
rect 57112 37204 57118 37256
rect 102134 37204 102140 37256
rect 102192 37244 102198 37256
rect 195974 37244 195980 37256
rect 102192 37216 195980 37244
rect 102192 37204 102198 37216
rect 195974 37204 195980 37216
rect 196032 37204 196038 37256
rect 102778 35844 102784 35896
rect 102836 35884 102842 35896
rect 195974 35884 195980 35896
rect 102836 35856 195980 35884
rect 102836 35844 102842 35856
rect 195974 35844 195980 35856
rect 196032 35844 196038 35896
rect 102686 35776 102692 35828
rect 102744 35816 102750 35828
rect 196066 35816 196072 35828
rect 102744 35788 196072 35816
rect 102744 35776 102750 35788
rect 196066 35776 196072 35788
rect 196124 35776 196130 35828
rect 102870 34416 102876 34468
rect 102928 34456 102934 34468
rect 195974 34456 195980 34468
rect 102928 34428 195980 34456
rect 102928 34416 102934 34428
rect 195974 34416 195980 34428
rect 196032 34416 196038 34468
rect 102594 34348 102600 34400
rect 102652 34388 102658 34400
rect 196066 34388 196072 34400
rect 102652 34360 196072 34388
rect 102652 34348 102658 34360
rect 196066 34348 196072 34360
rect 196124 34348 196130 34400
rect 102134 33056 102140 33108
rect 102192 33096 102198 33108
rect 195974 33096 195980 33108
rect 102192 33068 195980 33096
rect 102192 33056 102198 33068
rect 195974 33056 195980 33068
rect 196032 33056 196038 33108
rect 4982 31696 4988 31748
rect 5040 31736 5046 31748
rect 57606 31736 57612 31748
rect 5040 31708 57612 31736
rect 5040 31696 5046 31708
rect 57606 31696 57612 31708
rect 57664 31696 57670 31748
rect 102318 31696 102324 31748
rect 102376 31736 102382 31748
rect 195974 31736 195980 31748
rect 102376 31708 195980 31736
rect 102376 31696 102382 31708
rect 195974 31696 195980 31708
rect 196032 31696 196038 31748
rect 102134 31628 102140 31680
rect 102192 31668 102198 31680
rect 196066 31668 196072 31680
rect 102192 31640 196072 31668
rect 102192 31628 102198 31640
rect 196066 31628 196072 31640
rect 196124 31628 196130 31680
rect 102226 30268 102232 30320
rect 102284 30308 102290 30320
rect 195974 30308 195980 30320
rect 102284 30280 195980 30308
rect 102284 30268 102290 30280
rect 195974 30268 195980 30280
rect 196032 30268 196038 30320
rect 102134 30200 102140 30252
rect 102192 30240 102198 30252
rect 196066 30240 196072 30252
rect 102192 30212 196072 30240
rect 102192 30200 102198 30212
rect 196066 30200 196072 30212
rect 196124 30200 196130 30252
rect 102134 28908 102140 28960
rect 102192 28948 102198 28960
rect 195974 28948 195980 28960
rect 102192 28920 195980 28948
rect 102192 28908 102198 28920
rect 195974 28908 195980 28920
rect 196032 28908 196038 28960
rect 102134 28228 102140 28280
rect 102192 28268 102198 28280
rect 195974 28268 195980 28280
rect 102192 28240 195980 28268
rect 102192 28228 102198 28240
rect 195974 28228 195980 28240
rect 196032 28228 196038 28280
rect 17218 27548 17224 27600
rect 17276 27588 17282 27600
rect 57238 27588 57244 27600
rect 17276 27560 57244 27588
rect 17276 27548 17282 27560
rect 57238 27548 57244 27560
rect 57296 27548 57302 27600
rect 102134 27548 102140 27600
rect 102192 27588 102198 27600
rect 195974 27588 195980 27600
rect 102192 27560 195980 27588
rect 102192 27548 102198 27560
rect 195974 27548 195980 27560
rect 196032 27548 196038 27600
rect 102778 26188 102784 26240
rect 102836 26228 102842 26240
rect 195974 26228 195980 26240
rect 102836 26200 195980 26228
rect 102836 26188 102842 26200
rect 195974 26188 195980 26200
rect 196032 26188 196038 26240
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 356974 24256 356980 24268
rect 18656 24228 356980 24256
rect 18656 24216 18662 24228
rect 356974 24216 356980 24228
rect 357032 24216 357038 24268
rect 7558 24148 7564 24200
rect 7616 24188 7622 24200
rect 364426 24188 364432 24200
rect 7616 24160 364432 24188
rect 7616 24148 7622 24160
rect 364426 24148 364432 24160
rect 364484 24148 364490 24200
rect 382826 24148 382832 24200
rect 382884 24188 382890 24200
rect 398834 24188 398840 24200
rect 382884 24160 398840 24188
rect 382884 24148 382890 24160
rect 398834 24148 398840 24160
rect 398892 24148 398898 24200
rect 16482 24080 16488 24132
rect 16540 24120 16546 24132
rect 375006 24120 375012 24132
rect 16540 24092 375012 24120
rect 16540 24080 16546 24092
rect 375006 24080 375012 24092
rect 375064 24080 375070 24132
rect 393314 24080 393320 24132
rect 393372 24120 393378 24132
rect 569218 24120 569224 24132
rect 393372 24092 569224 24120
rect 393372 24080 393378 24092
rect 569218 24080 569224 24092
rect 569276 24080 569282 24132
rect 85482 23468 85488 23520
rect 85540 23508 85546 23520
rect 266354 23508 266360 23520
rect 85540 23480 266360 23508
rect 85540 23468 85546 23480
rect 266354 23468 266360 23480
rect 266412 23508 266418 23520
rect 267366 23508 267372 23520
rect 266412 23480 267372 23508
rect 266412 23468 266418 23480
rect 267366 23468 267372 23480
rect 267424 23468 267430 23520
rect 59998 22244 60004 22296
rect 60056 22284 60062 22296
rect 353754 22284 353760 22296
rect 60056 22256 353760 22284
rect 60056 22244 60062 22256
rect 353754 22244 353760 22256
rect 353812 22244 353818 22296
rect 3510 22176 3516 22228
rect 3568 22216 3574 22228
rect 335814 22216 335820 22228
rect 3568 22188 335820 22216
rect 3568 22176 3574 22188
rect 335814 22176 335820 22188
rect 335872 22176 335878 22228
rect 3602 22108 3608 22160
rect 3660 22148 3666 22160
rect 346578 22148 346584 22160
rect 3660 22120 346584 22148
rect 3660 22108 3666 22120
rect 346578 22108 346584 22120
rect 346636 22108 346642 22160
rect 62298 22040 62304 22092
rect 62356 22080 62362 22092
rect 85482 22080 85488 22092
rect 62356 22052 85488 22080
rect 62356 22040 62362 22052
rect 85482 22040 85488 22052
rect 85540 22040 85546 22092
rect 199378 22040 199384 22092
rect 199436 22080 199442 22092
rect 350166 22080 350172 22092
rect 199436 22052 350172 22080
rect 199436 22040 199442 22052
rect 350166 22040 350172 22052
rect 350224 22040 350230 22092
rect 386046 22040 386052 22092
rect 386104 22080 386110 22092
rect 574094 22080 574100 22092
rect 386104 22052 574100 22080
rect 386104 22040 386110 22052
rect 574094 22040 574100 22052
rect 574152 22040 574158 22092
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 371694 22012 371700 22024
rect 3476 21984 371700 22012
rect 3476 21972 3482 21984
rect 371694 21972 371700 21984
rect 371752 21972 371758 22024
rect 396810 21972 396816 22024
rect 396868 22012 396874 22024
rect 570598 22012 570604 22024
rect 396868 21984 570604 22012
rect 396868 21972 396874 21984
rect 570598 21972 570604 21984
rect 570656 21972 570662 22024
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 360930 21944 360936 21956
rect 18748 21916 360936 21944
rect 18748 21904 18754 21916
rect 360930 21904 360936 21916
rect 360988 21904 360994 21956
rect 378870 21904 378876 21956
rect 378928 21944 378934 21956
rect 400214 21944 400220 21956
rect 378928 21916 400220 21944
rect 378928 21904 378934 21916
rect 400214 21904 400220 21916
rect 400272 21904 400278 21956
rect 175458 21496 175464 21548
rect 175516 21536 175522 21548
rect 285582 21536 285588 21548
rect 175516 21508 285588 21536
rect 175516 21496 175522 21508
rect 285582 21496 285588 21508
rect 285640 21496 285646 21548
rect 187694 21428 187700 21480
rect 187752 21468 187758 21480
rect 299934 21468 299940 21480
rect 187752 21440 299940 21468
rect 187752 21428 187758 21440
rect 299934 21428 299940 21440
rect 299992 21428 299998 21480
rect 152458 21360 152464 21412
rect 152516 21400 152522 21412
rect 292758 21400 292764 21412
rect 152516 21372 292764 21400
rect 152516 21360 152522 21372
rect 292758 21360 292764 21372
rect 292816 21360 292822 21412
rect 178034 20068 178040 20120
rect 178092 20108 178098 20120
rect 256878 20108 256884 20120
rect 178092 20080 256884 20108
rect 178092 20068 178098 20080
rect 256878 20068 256884 20080
rect 256936 20068 256942 20120
rect 162854 20000 162860 20052
rect 162912 20040 162918 20052
rect 307110 20040 307116 20052
rect 162912 20012 307116 20040
rect 162912 20000 162918 20012
rect 307110 20000 307116 20012
rect 307168 20000 307174 20052
rect 138014 19932 138020 19984
rect 138072 19972 138078 19984
rect 281994 19972 282000 19984
rect 138072 19944 282000 19972
rect 138072 19932 138078 19944
rect 281994 19932 282000 19944
rect 282052 19932 282058 19984
rect 155954 18776 155960 18828
rect 156012 18816 156018 18828
rect 187694 18816 187700 18828
rect 156012 18788 187700 18816
rect 156012 18776 156018 18788
rect 187694 18776 187700 18788
rect 187752 18776 187758 18828
rect 175274 18708 175280 18760
rect 175332 18748 175338 18760
rect 253290 18748 253296 18760
rect 175332 18720 253296 18748
rect 175332 18708 175338 18720
rect 253290 18708 253296 18720
rect 253348 18708 253354 18760
rect 150434 18640 150440 18692
rect 150492 18680 150498 18692
rect 228174 18680 228180 18692
rect 150492 18652 228180 18680
rect 150492 18640 150498 18652
rect 228174 18640 228180 18652
rect 228232 18640 228238 18692
rect 142154 18572 142160 18624
rect 142212 18612 142218 18624
rect 175458 18612 175464 18624
rect 142212 18584 175464 18612
rect 142212 18572 142218 18584
rect 175458 18572 175464 18584
rect 175516 18572 175522 18624
rect 184934 18572 184940 18624
rect 184992 18612 184998 18624
rect 328638 18612 328644 18624
rect 184992 18584 328644 18612
rect 184992 18572 184998 18584
rect 328638 18572 328644 18584
rect 328696 18572 328702 18624
rect 171134 17348 171140 17400
rect 171192 17388 171198 17400
rect 249702 17388 249708 17400
rect 171192 17360 249708 17388
rect 171192 17348 171198 17360
rect 249702 17348 249708 17360
rect 249760 17348 249766 17400
rect 131114 17280 131120 17332
rect 131172 17320 131178 17332
rect 274818 17320 274824 17332
rect 131172 17292 274824 17320
rect 131172 17280 131178 17292
rect 274818 17280 274824 17292
rect 274876 17280 274882 17332
rect 71130 17212 71136 17264
rect 71188 17252 71194 17264
rect 242894 17252 242900 17264
rect 71188 17224 242900 17252
rect 71188 17212 71194 17224
rect 242894 17212 242900 17224
rect 242952 17212 242958 17264
rect 168374 15988 168380 16040
rect 168432 16028 168438 16040
rect 245654 16028 245660 16040
rect 168432 16000 245660 16028
rect 168432 15988 168438 16000
rect 245654 15988 245660 16000
rect 245712 15988 245718 16040
rect 135254 15920 135260 15972
rect 135312 15960 135318 15972
rect 277394 15960 277400 15972
rect 135312 15932 277400 15960
rect 135312 15920 135318 15932
rect 277394 15920 277400 15932
rect 277452 15920 277458 15972
rect 74534 15852 74540 15904
rect 74592 15892 74598 15904
rect 245930 15892 245936 15904
rect 74592 15864 245936 15892
rect 74592 15852 74598 15864
rect 245930 15852 245936 15864
rect 245988 15852 245994 15904
rect 136450 14560 136456 14612
rect 136508 14600 136514 14612
rect 212534 14600 212540 14612
rect 136508 14572 212540 14600
rect 136508 14560 136514 14572
rect 212534 14560 212540 14572
rect 212592 14560 212598 14612
rect 164418 14492 164424 14544
rect 164476 14532 164482 14544
rect 241514 14532 241520 14544
rect 164476 14504 241520 14532
rect 164476 14492 164482 14504
rect 241514 14492 241520 14504
rect 241572 14492 241578 14544
rect 170306 14424 170312 14476
rect 170364 14464 170370 14476
rect 313274 14464 313280 14476
rect 170364 14436 313280 14464
rect 170364 14424 170370 14436
rect 313274 14424 313280 14436
rect 313332 14424 313338 14476
rect 139578 13200 139584 13252
rect 139636 13240 139642 13252
rect 216674 13240 216680 13252
rect 139636 13212 216680 13240
rect 139636 13200 139642 13212
rect 216674 13200 216680 13212
rect 216732 13200 216738 13252
rect 160094 13132 160100 13184
rect 160152 13172 160158 13184
rect 238754 13172 238760 13184
rect 160152 13144 238760 13172
rect 160152 13132 160158 13144
rect 238754 13132 238760 13144
rect 238812 13132 238818 13184
rect 176654 13064 176660 13116
rect 176712 13104 176718 13116
rect 320174 13104 320180 13116
rect 176712 13076 320180 13104
rect 176712 13064 176718 13076
rect 320174 13064 320180 13076
rect 320232 13064 320238 13116
rect 153746 11908 153752 11960
rect 153804 11948 153810 11960
rect 230474 11948 230480 11960
rect 153804 11920 230480 11948
rect 153804 11908 153810 11920
rect 230474 11908 230480 11920
rect 230532 11908 230538 11960
rect 125594 11840 125600 11892
rect 125652 11880 125658 11892
rect 202874 11880 202880 11892
rect 125652 11852 202880 11880
rect 125652 11840 125658 11852
rect 202874 11840 202880 11852
rect 202932 11840 202938 11892
rect 186130 11772 186136 11824
rect 186188 11812 186194 11824
rect 263594 11812 263600 11824
rect 186188 11784 263600 11812
rect 186188 11772 186194 11784
rect 263594 11772 263600 11784
rect 263652 11772 263658 11824
rect 151814 11704 151820 11756
rect 151872 11744 151878 11756
rect 295334 11744 295340 11756
rect 151872 11716 295340 11744
rect 151872 11704 151878 11716
rect 295334 11704 295340 11716
rect 295392 11704 295398 11756
rect 156598 10412 156604 10464
rect 156656 10452 156662 10464
rect 209774 10452 209780 10464
rect 156656 10424 209780 10452
rect 156656 10412 156662 10424
rect 209774 10412 209780 10424
rect 209832 10412 209838 10464
rect 147122 10344 147128 10396
rect 147180 10384 147186 10396
rect 223574 10384 223580 10396
rect 147180 10356 223580 10384
rect 147180 10344 147186 10356
rect 223574 10344 223580 10356
rect 223632 10344 223638 10396
rect 3418 10276 3424 10328
rect 3476 10316 3482 10328
rect 338114 10316 338120 10328
rect 3476 10288 338120 10316
rect 3476 10276 3482 10288
rect 338114 10276 338120 10288
rect 338172 10276 338178 10328
rect 174262 9052 174268 9104
rect 174320 9092 174326 9104
rect 317414 9092 317420 9104
rect 174320 9064 317420 9092
rect 174320 9052 174326 9064
rect 317414 9052 317420 9064
rect 317472 9052 317478 9104
rect 167178 8984 167184 9036
rect 167236 9024 167242 9036
rect 310514 9024 310520 9036
rect 167236 8996 310520 9024
rect 167236 8984 167242 8996
rect 310514 8984 310520 8996
rect 310572 8984 310578 9036
rect 84194 8916 84200 8968
rect 84252 8956 84258 8968
rect 241698 8956 241704 8968
rect 84252 8928 241704 8956
rect 84252 8916 84258 8928
rect 241698 8916 241704 8928
rect 241756 8916 241762 8968
rect 157794 7692 157800 7744
rect 157852 7732 157858 7744
rect 234614 7732 234620 7744
rect 157852 7704 234620 7732
rect 157852 7692 157858 7704
rect 234614 7692 234620 7704
rect 234672 7692 234678 7744
rect 235902 7692 235908 7744
rect 235960 7732 235966 7744
rect 288434 7732 288440 7744
rect 235960 7704 288440 7732
rect 235960 7692 235966 7704
rect 288434 7692 288440 7704
rect 288492 7692 288498 7744
rect 128170 7624 128176 7676
rect 128228 7664 128234 7676
rect 270494 7664 270500 7676
rect 128228 7636 270500 7664
rect 128228 7624 128234 7636
rect 270494 7624 270500 7636
rect 270552 7624 270558 7676
rect 88334 7556 88340 7608
rect 88392 7596 88398 7608
rect 245194 7596 245200 7608
rect 88392 7568 245200 7596
rect 88392 7556 88398 7568
rect 245194 7556 245200 7568
rect 245252 7556 245258 7608
rect 143534 6332 143540 6384
rect 143592 6372 143598 6384
rect 220814 6372 220820 6384
rect 143592 6344 220820 6372
rect 143592 6332 143598 6344
rect 220814 6332 220820 6344
rect 220872 6332 220878 6384
rect 181438 6264 181444 6316
rect 181496 6304 181502 6316
rect 324314 6304 324320 6316
rect 181496 6276 324320 6304
rect 181496 6264 181502 6276
rect 324314 6264 324320 6276
rect 324372 6264 324378 6316
rect 92474 6196 92480 6248
rect 92532 6236 92538 6248
rect 248782 6236 248788 6248
rect 92532 6208 248788 6236
rect 92532 6196 92538 6208
rect 248782 6196 248788 6208
rect 248840 6196 248846 6248
rect 78674 6128 78680 6180
rect 78732 6168 78738 6180
rect 249978 6168 249984 6180
rect 78732 6140 249984 6168
rect 78732 6128 78738 6140
rect 249978 6128 249984 6140
rect 250036 6128 250042 6180
rect 182542 4972 182548 5024
rect 182600 5012 182606 5024
rect 259454 5012 259460 5024
rect 182600 4984 259460 5012
rect 182600 4972 182606 4984
rect 259454 4972 259460 4984
rect 259512 4972 259518 5024
rect 129366 4904 129372 4956
rect 129424 4944 129430 4956
rect 205634 4944 205640 4956
rect 129424 4916 205640 4944
rect 129424 4904 129430 4916
rect 205634 4904 205640 4916
rect 205692 4904 205698 4956
rect 188522 4836 188528 4888
rect 188580 4876 188586 4888
rect 331214 4876 331220 4888
rect 188580 4848 331220 4876
rect 188580 4836 188586 4848
rect 331214 4836 331220 4848
rect 331272 4836 331278 4888
rect 96614 4768 96620 4820
rect 96672 4808 96678 4820
rect 252370 4808 252376 4820
rect 96672 4780 252376 4808
rect 96672 4768 96678 4780
rect 252370 4768 252376 4780
rect 252428 4768 252434 4820
rect 149514 3816 149520 3868
rect 149572 3856 149578 3868
rect 152458 3856 152464 3868
rect 149572 3828 152464 3856
rect 149572 3816 149578 3828
rect 152458 3816 152464 3828
rect 152516 3816 152522 3868
rect 145926 3544 145932 3596
rect 145984 3584 145990 3596
rect 235902 3584 235908 3596
rect 145984 3556 235908 3584
rect 145984 3544 145990 3556
rect 235902 3544 235908 3556
rect 235960 3544 235966 3596
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 156598 3516 156604 3528
rect 133012 3488 156604 3516
rect 133012 3476 133018 3488
rect 156598 3476 156604 3488
rect 156656 3476 156662 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 161382 3476 161388 3528
rect 161440 3516 161446 3528
rect 302234 3516 302240 3528
rect 161440 3488 302240 3516
rect 161440 3476 161446 3488
rect 302234 3476 302240 3488
rect 302292 3476 302298 3528
rect 66254 3408 66260 3460
rect 66312 3448 66318 3460
rect 239306 3448 239312 3460
rect 66312 3420 239312 3448
rect 66312 3408 66318 3420
rect 239306 3408 239312 3420
rect 239364 3408 239370 3460
rect 266354 3408 266360 3460
rect 266412 3448 266418 3460
rect 579798 3448 579804 3460
rect 266412 3420 579804 3448
rect 266412 3408 266418 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 151814 3340 151820 3392
rect 151872 3380 151878 3392
rect 153010 3380 153016 3392
rect 151872 3352 153016 3380
rect 151872 3340 151878 3352
rect 153010 3340 153016 3352
rect 153068 3340 153074 3392
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 177850 3380 177856 3392
rect 176712 3352 177856 3380
rect 176712 3340 176718 3352
rect 177850 3340 177856 3352
rect 177908 3340 177914 3392
rect 160094 2796 160100 2848
rect 160152 2836 160158 2848
rect 161382 2836 161388 2848
rect 160152 2808 161388 2836
rect 160152 2796 160158 2808
rect 161382 2796 161388 2808
rect 161440 2796 161446 2848
<< via1 >>
rect 137836 700952 137888 701004
rect 202788 700952 202840 701004
rect 397460 700952 397512 701004
rect 462320 700952 462372 701004
rect 8116 700476 8168 700528
rect 16488 700476 16540 700528
rect 72976 700476 73028 700528
rect 295248 700476 295300 700528
rect 397460 700476 397512 700528
rect 20628 700408 20680 700460
rect 89168 700408 89220 700460
rect 300584 700408 300636 700460
rect 413652 700408 413704 700460
rect 20444 700340 20496 700392
rect 154120 700340 154172 700392
rect 300676 700340 300728 700392
rect 478512 700340 478564 700392
rect 20352 700272 20404 700324
rect 218980 700272 219032 700324
rect 300768 700272 300820 700324
rect 543464 700272 543516 700324
rect 20536 699660 20588 699712
rect 24308 699660 24360 699712
rect 527180 697552 527232 697604
rect 574100 697552 574152 697604
rect 574100 696940 574152 696992
rect 580172 696940 580224 696992
rect 3424 671032 3476 671084
rect 7656 671032 7708 671084
rect 2872 618876 2924 618928
rect 4988 618876 5040 618928
rect 300584 588616 300636 588668
rect 304172 588616 304224 588668
rect 300676 586508 300728 586560
rect 310336 586508 310388 586560
rect 20444 586440 20496 586492
rect 24216 586440 24268 586492
rect 129188 586440 129240 586492
rect 134340 586440 134392 586492
rect 198648 586440 198700 586492
rect 292580 586440 292632 586492
rect 408868 586440 408920 586492
rect 414664 586440 414716 586492
rect 20352 586372 20404 586424
rect 30012 586372 30064 586424
rect 559564 586168 559616 586220
rect 569960 586168 570012 586220
rect 22008 586100 22060 586152
rect 47400 586100 47452 586152
rect 300492 586100 300544 586152
rect 316132 586100 316184 586152
rect 553768 586100 553820 586152
rect 572720 586100 572772 586152
rect 20444 586032 20496 586084
rect 53196 586032 53248 586084
rect 279884 586032 279936 586084
rect 290004 586032 290056 586084
rect 300676 586032 300728 586084
rect 321928 586032 321980 586084
rect 547972 586032 548024 586084
rect 570144 586032 570196 586084
rect 17868 585964 17920 586016
rect 58992 585964 59044 586016
rect 268292 585964 268344 586016
rect 289912 585964 289964 586016
rect 302148 585964 302200 586016
rect 327724 585964 327776 586016
rect 542176 585964 542228 586016
rect 570052 585964 570104 586016
rect 20352 585896 20404 585948
rect 35900 585896 35952 585948
rect 37924 585896 37976 585948
rect 105360 585896 105412 585948
rect 262128 585896 262180 585948
rect 289820 585896 289872 585948
rect 300584 585896 300636 585948
rect 333520 585896 333572 585948
rect 536380 585896 536432 585948
rect 568580 585896 568632 585948
rect 31024 585828 31076 585880
rect 99564 585828 99616 585880
rect 256608 585828 256660 585880
rect 288440 585828 288492 585880
rect 297824 585828 297876 585880
rect 339316 585828 339368 585880
rect 524788 585828 524840 585880
rect 569316 585828 569368 585880
rect 20260 585760 20312 585812
rect 41604 585760 41656 585812
rect 43444 585760 43496 585812
rect 116952 585760 117004 585812
rect 250904 585760 250956 585812
rect 288624 585760 288676 585812
rect 299388 585760 299440 585812
rect 345112 585760 345164 585812
rect 507400 585760 507452 585812
rect 568672 585760 568724 585812
rect 17684 583380 17736 583432
rect 76380 583380 76432 583432
rect 233148 583380 233200 583432
rect 291292 583380 291344 583432
rect 17776 583312 17828 583364
rect 87972 583312 88024 583364
rect 221924 583312 221976 583364
rect 292764 583312 292816 583364
rect 513196 583312 513248 583364
rect 571524 583312 571576 583364
rect 19156 583244 19208 583296
rect 93860 583244 93912 583296
rect 216128 583244 216180 583296
rect 291200 583244 291252 583296
rect 297732 583244 297784 583296
rect 356704 583244 356756 583296
rect 501604 583244 501656 583296
rect 571432 583244 571484 583296
rect 15016 583176 15068 583228
rect 111156 583176 111208 583228
rect 210332 583176 210384 583228
rect 292580 583176 292632 583228
rect 298836 583176 298888 583228
rect 368296 583176 368348 583228
rect 490012 583176 490064 583228
rect 574192 583176 574244 583228
rect 19064 583108 19116 583160
rect 122840 583108 122892 583160
rect 204168 583108 204220 583160
rect 291384 583108 291436 583160
rect 299204 583108 299256 583160
rect 374092 583108 374144 583160
rect 484216 583108 484268 583160
rect 571616 583108 571668 583160
rect 15108 583040 15160 583092
rect 140136 583040 140188 583092
rect 192944 583040 192996 583092
rect 293960 583040 294012 583092
rect 297916 583040 297968 583092
rect 379888 583040 379940 583092
rect 472624 583040 472676 583092
rect 572812 583040 572864 583092
rect 16396 582972 16448 583024
rect 151820 582972 151872 583024
rect 175188 582972 175240 583024
rect 291844 582972 291896 583024
rect 296628 582972 296680 583024
rect 391480 582972 391532 583024
rect 455236 582972 455288 583024
rect 571340 582972 571392 583024
rect 296536 580524 296588 580576
rect 397276 580524 397328 580576
rect 300400 580456 300452 580508
rect 403072 580456 403124 580508
rect 181352 580388 181404 580440
rect 293224 580388 293276 580440
rect 296444 580388 296496 580440
rect 420460 580388 420512 580440
rect 158168 580320 158220 580372
rect 288532 580320 288584 580372
rect 298008 580320 298060 580372
rect 426256 580320 426308 580372
rect 14924 580252 14976 580304
rect 145932 580252 145984 580304
rect 163964 580252 164016 580304
rect 294052 580252 294104 580304
rect 299112 580252 299164 580304
rect 432052 580252 432104 580304
rect 449440 580252 449492 580304
rect 572904 580252 572956 580304
rect 273260 572160 273312 572212
rect 294604 572160 294656 572212
rect 529940 572160 529992 572212
rect 570236 572160 570288 572212
rect 18604 572092 18656 572144
rect 31024 572092 31076 572144
rect 244280 572092 244332 572144
rect 290096 572092 290148 572144
rect 495440 572092 495492 572144
rect 571708 572092 571760 572144
rect 17592 572024 17644 572076
rect 37924 572024 37976 572076
rect 186320 572024 186372 572076
rect 290188 572024 290240 572076
rect 460940 572024 460992 572076
rect 572996 572024 573048 572076
rect 18696 571956 18748 572008
rect 43444 571956 43496 572008
rect 168380 571956 168432 572008
rect 293316 571956 293368 572008
rect 443000 571956 443052 572008
rect 575572 571956 575624 572008
rect 569224 485052 569276 485104
rect 580540 485052 580592 485104
rect 580908 485052 580960 485104
rect 19064 463360 19116 463412
rect 23388 463360 23440 463412
rect 291844 462544 291896 462596
rect 292948 462544 293000 462596
rect 2780 462408 2832 462460
rect 4804 462408 4856 462460
rect 24860 462408 24912 462460
rect 140136 462408 140188 462460
rect 296628 462408 296680 462460
rect 391204 462408 391256 462460
rect 438216 462408 438268 462460
rect 568764 462408 568816 462460
rect 575480 462408 575532 462460
rect 14832 462272 14884 462324
rect 15016 462272 15068 462324
rect 16396 462272 16448 462324
rect 151912 462340 151964 462392
rect 292580 462340 292632 462392
rect 293224 462340 293276 462392
rect 296720 462340 296772 462392
rect 300124 462340 300176 462392
rect 402888 462340 402940 462392
rect 443736 462340 443788 462392
rect 575572 462340 575624 462392
rect 288256 462272 288308 462324
rect 288532 462272 288584 462324
rect 291476 462272 291528 462324
rect 294052 462272 294104 462324
rect 297824 462272 297876 462324
rect 300216 462272 300268 462324
rect 300768 462272 300820 462324
rect 304172 462272 304224 462324
rect 570328 462272 570380 462324
rect 571616 462272 571668 462324
rect 20536 462204 20588 462256
rect 24216 462204 24268 462256
rect 297732 462204 297784 462256
rect 298744 462204 298796 462256
rect 300676 462204 300728 462256
rect 302148 462204 302200 462256
rect 300308 461864 300360 461916
rect 300584 461864 300636 461916
rect 15108 461592 15160 461644
rect 17408 461592 17460 461644
rect 24860 461592 24912 461644
rect 291292 461320 291344 461372
rect 291568 461320 291620 461372
rect 455328 461320 455380 461372
rect 567108 461320 567160 461372
rect 571340 461320 571392 461372
rect 158168 461252 158220 461304
rect 288256 461252 288308 461304
rect 233332 461184 233384 461236
rect 513288 461252 513340 461304
rect 571524 461252 571576 461304
rect 300216 461184 300268 461236
rect 336740 461184 336792 461236
rect 507768 461184 507820 461236
rect 567752 461184 567804 461236
rect 568672 461184 568724 461236
rect 181352 461116 181404 461168
rect 292580 461116 292632 461168
rect 299296 461116 299348 461168
rect 302056 461116 302108 461168
rect 327356 461116 327408 461168
rect 501880 461116 501932 461168
rect 571432 461116 571484 461168
rect 574652 461116 574704 461168
rect 175234 461048 175286 461100
rect 291844 461048 291896 461100
rect 300308 461048 300360 461100
rect 333520 461048 333572 461100
rect 484216 461048 484268 461100
rect 570328 461048 570380 461100
rect 14832 460980 14884 461032
rect 26240 460980 26292 461032
rect 163642 460980 163694 461032
rect 291476 460980 291528 461032
rect 303528 460980 303580 461032
rect 350908 460980 350960 461032
rect 561588 460980 561640 461032
rect 574192 460980 574244 461032
rect 14924 460844 14976 460896
rect 145932 460912 145984 460964
rect 280712 460912 280764 460964
rect 292488 460912 292540 460964
rect 298744 460912 298796 460964
rect 356704 460912 356756 460964
rect 449440 460912 449492 460964
rect 572904 460912 572956 460964
rect 192944 460844 192996 460896
rect 293960 460844 294012 460896
rect 296536 460844 296588 460896
rect 397276 460844 397328 460896
rect 461032 460844 461084 460896
rect 572996 460844 573048 460896
rect 15016 459620 15068 459672
rect 18696 459620 18748 459672
rect 16304 459552 16356 459604
rect 18604 459552 18656 459604
rect 20260 459552 20312 459604
rect 20628 459484 20680 459536
rect 30012 459484 30064 459536
rect 293960 459552 294012 459604
rect 295432 459552 295484 459604
rect 569316 459552 569368 459604
rect 571616 459552 571668 459604
rect 572996 459552 573048 459604
rect 574284 459552 574336 459604
rect 41604 459484 41656 459536
rect 129188 459484 129240 459536
rect 134340 459484 134392 459536
rect 187148 459484 187200 459536
rect 290280 459484 290332 459536
rect 318800 459484 318852 459536
rect 321928 459484 321980 459536
rect 336740 459484 336792 459536
rect 339316 459484 339368 459536
rect 408868 459484 408920 459536
rect 414664 459484 414716 459536
rect 466828 459484 466880 459536
rect 567936 459484 567988 459536
rect 568488 459484 568540 459536
rect 204168 459416 204220 459468
rect 291384 459416 291436 459468
rect 297824 459416 297876 459468
rect 379888 459416 379940 459468
rect 559564 459416 559616 459468
rect 569960 459416 570012 459468
rect 18604 459348 18656 459400
rect 99564 459348 99616 459400
rect 216128 459348 216180 459400
rect 291200 459348 291252 459400
rect 299020 459348 299072 459400
rect 374092 459348 374144 459400
rect 524788 459348 524840 459400
rect 569316 459348 569368 459400
rect 17776 459280 17828 459332
rect 87972 459280 88024 459332
rect 221924 459280 221976 459332
rect 292764 459280 292816 459332
rect 299388 459280 299440 459332
rect 345112 459280 345164 459332
rect 530584 459280 530636 459332
rect 570236 459280 570288 459332
rect 18696 459212 18748 459264
rect 116952 459212 117004 459264
rect 210332 459212 210384 459264
rect 280712 459212 280764 459264
rect 305000 459212 305052 459264
rect 316132 459212 316184 459264
rect 547972 459212 548024 459264
rect 570144 459212 570196 459264
rect 17592 459144 17644 459196
rect 105360 459144 105412 459196
rect 279884 459144 279936 459196
rect 290004 459144 290056 459196
rect 299204 459144 299256 459196
rect 385684 459144 385736 459196
rect 490012 459144 490064 459196
rect 561588 459144 561640 459196
rect 30932 459008 30984 459060
rect 35900 459008 35952 459060
rect 274088 458872 274140 458924
rect 294696 458872 294748 458924
rect 300400 458872 300452 458924
rect 368296 458872 368348 458924
rect 19248 458668 19300 458720
rect 20536 458668 20588 458720
rect 64880 458804 64932 458856
rect 268292 458804 268344 458856
rect 280068 458804 280120 458856
rect 289084 458804 289136 458856
rect 408868 458804 408920 458856
rect 495808 458804 495860 458856
rect 569316 458804 569368 458856
rect 571708 458804 571760 458856
rect 298836 458668 298888 458720
rect 300400 458668 300452 458720
rect 569960 458532 570012 458584
rect 570420 458532 570472 458584
rect 569960 458396 570012 458448
rect 570144 458396 570196 458448
rect 291200 458260 291252 458312
rect 292856 458260 292908 458312
rect 17500 458192 17552 458244
rect 17776 458192 17828 458244
rect 291384 458192 291436 458244
rect 292672 458192 292724 458244
rect 293316 458192 293368 458244
rect 293960 458192 294012 458244
rect 299112 458192 299164 458244
rect 299388 458192 299440 458244
rect 565360 458192 565412 458244
rect 568948 458192 569000 458244
rect 570236 458192 570288 458244
rect 571524 458192 571576 458244
rect 26240 458124 26292 458176
rect 111156 458124 111208 458176
rect 169668 458124 169720 458176
rect 518992 458124 519044 458176
rect 565820 458124 565872 458176
rect 570420 458124 570472 458176
rect 571708 458124 571760 458176
rect 19156 458056 19208 458108
rect 93860 458056 93912 458108
rect 245108 458056 245160 458108
rect 290096 458056 290148 458108
rect 536380 458056 536432 458108
rect 568672 458056 568724 458108
rect 17684 457988 17736 458040
rect 76380 457988 76432 458040
rect 250904 457988 250956 458040
rect 288624 457988 288676 458040
rect 291384 457988 291436 458040
rect 542176 457988 542228 458040
rect 570052 457988 570104 458040
rect 20444 457920 20496 457972
rect 53196 457920 53248 457972
rect 256608 457920 256660 457972
rect 287612 457920 287664 457972
rect 288440 457920 288492 457972
rect 21916 457852 21968 457904
rect 47400 457852 47452 457904
rect 262128 457852 262180 457904
rect 289820 457852 289872 457904
rect 280068 457444 280120 457496
rect 289176 457444 289228 457496
rect 289912 457444 289964 457496
rect 305000 457444 305052 457496
rect 426440 457444 426492 457496
rect 55956 456832 56008 456884
rect 58992 456832 59044 456884
rect 306380 456696 306432 456748
rect 420460 456696 420512 456748
rect 298008 456492 298060 456544
rect 299204 456492 299256 456544
rect 305000 456492 305052 456544
rect 288256 456288 288308 456340
rect 290188 456288 290240 456340
rect 17868 456016 17920 456068
rect 19156 456016 19208 456068
rect 55956 456016 56008 456068
rect 307668 456016 307720 456068
rect 432052 456016 432104 456068
rect 297916 455336 297968 455388
rect 302240 455336 302292 455388
rect 307668 455336 307720 455388
rect 471980 444320 472032 444372
rect 572812 444320 572864 444372
rect 284300 443640 284352 443692
rect 297364 443640 297416 443692
rect 567108 443640 567160 443692
rect 570236 443640 570288 443692
rect 19064 443368 19116 443420
rect 23480 443368 23532 443420
rect 2872 409912 2924 409964
rect 4896 409912 4948 409964
rect 2780 398692 2832 398744
rect 7564 398692 7616 398744
rect 570604 378768 570656 378820
rect 580448 378768 580500 378820
rect 580908 378768 580960 378820
rect 3332 357416 3384 357468
rect 18604 357416 18656 357468
rect 3332 345040 3384 345092
rect 18696 345040 18748 345092
rect 14924 333956 14976 334008
rect 27528 333956 27580 334008
rect 292488 333956 292540 334008
rect 295616 333956 295668 334008
rect 19156 333276 19208 333328
rect 21824 333276 21876 333328
rect 17408 333208 17460 333260
rect 26240 333208 26292 333260
rect 286968 333276 287020 333328
rect 291476 333276 291528 333328
rect 291752 333276 291804 333328
rect 292856 333276 292908 333328
rect 281448 333208 281500 333260
rect 290280 333208 290332 333260
rect 296628 333208 296680 333260
rect 306380 333208 306432 333260
rect 567108 333208 567160 333260
rect 570328 333208 570380 333260
rect 300216 333140 300268 333192
rect 300768 333140 300820 333192
rect 56508 332936 56560 332988
rect 250904 332936 250956 332988
rect 291292 332936 291344 332988
rect 300768 332936 300820 332988
rect 338948 332936 339000 332988
rect 19064 332868 19116 332920
rect 122748 332868 122800 332920
rect 239312 332868 239364 332920
rect 282184 332868 282236 332920
rect 299112 332868 299164 332920
rect 342260 332868 342312 332920
rect 22008 332800 22060 332852
rect 82176 332800 82228 332852
rect 169760 332800 169812 332852
rect 294052 332800 294104 332852
rect 299020 332800 299072 332852
rect 373908 332800 373960 332852
rect 16304 332732 16356 332784
rect 99564 332732 99616 332784
rect 216128 332732 216180 332784
rect 291752 332732 291804 332784
rect 302056 332732 302108 332784
rect 368296 332732 368348 332784
rect 513196 332732 513248 332784
rect 571340 332868 571392 332920
rect 4988 332664 5040 332716
rect 24216 332664 24268 332716
rect 27528 332664 27580 332716
rect 111156 332664 111208 332716
rect 210332 332664 210384 332716
rect 292488 332664 292540 332716
rect 296260 332664 296312 332716
rect 297824 332664 297876 332716
rect 379888 332664 379940 332716
rect 472624 332664 472676 332716
rect 572812 332732 572864 332784
rect 574560 332732 574612 332784
rect 571340 332664 571392 332716
rect 572996 332664 573048 332716
rect 17592 332596 17644 332648
rect 105360 332596 105412 332648
rect 181352 332596 181404 332648
rect 292580 332596 292632 332648
rect 296720 332596 296772 332648
rect 298836 332596 298888 332648
rect 299020 332596 299072 332648
rect 304540 332596 304592 332648
rect 580356 332596 580408 332648
rect 7656 332528 7708 332580
rect 30012 332528 30064 332580
rect 21916 332460 21968 332512
rect 31024 332528 31076 332580
rect 56508 332528 56560 332580
rect 58992 332528 59044 332580
rect 129188 332528 129240 332580
rect 134984 332528 135036 332580
rect 256608 332528 256660 332580
rect 287796 332528 287848 332580
rect 342260 332528 342312 332580
rect 345112 332528 345164 332580
rect 408868 332528 408920 332580
rect 414664 332528 414716 332580
rect 524788 332528 524840 332580
rect 571616 332528 571668 332580
rect 20536 332392 20588 332444
rect 64972 332460 65024 332512
rect 262128 332460 262180 332512
rect 289820 332460 289872 332512
rect 300308 332460 300360 332512
rect 333520 332460 333572 332512
rect 518992 332460 519044 332512
rect 565820 332460 565872 332512
rect 20444 332324 20496 332376
rect 53196 332392 53248 332444
rect 268292 332392 268344 332444
rect 289176 332392 289228 332444
rect 293040 332392 293092 332444
rect 299296 332392 299348 332444
rect 327724 332392 327776 332444
rect 536380 332392 536432 332444
rect 568672 332392 568724 332444
rect 31024 332324 31076 332376
rect 47400 332324 47452 332376
rect 279884 332324 279936 332376
rect 290004 332324 290056 332376
rect 302148 332324 302200 332376
rect 321928 332324 321980 332376
rect 542176 332324 542228 332376
rect 570052 332324 570104 332376
rect 20260 332256 20312 332308
rect 41604 332256 41656 332308
rect 300584 332256 300636 332308
rect 316132 332256 316184 332308
rect 547972 332256 548024 332308
rect 569960 332256 570012 332308
rect 20352 332188 20404 332240
rect 35992 332188 36044 332240
rect 303528 332188 303580 332240
rect 350908 332188 350960 332240
rect 559564 332188 559616 332240
rect 571892 332188 571944 332240
rect 23388 332120 23440 332172
rect 70584 332120 70636 332172
rect 289820 332052 289872 332104
rect 293960 332052 294012 332104
rect 285588 331984 285640 332036
rect 290556 331984 290608 332036
rect 198648 331916 198700 331968
rect 289820 331916 289872 331968
rect 290464 331916 290516 331968
rect 408868 331916 408920 331968
rect 443644 331916 443696 331968
rect 561588 331916 561640 331968
rect 134984 331848 135036 331900
rect 288440 331848 288492 331900
rect 297456 331848 297508 331900
rect 478420 331848 478472 331900
rect 565360 331848 565412 331900
rect 571340 331848 571392 331900
rect 282184 331712 282236 331764
rect 285588 331712 285640 331764
rect 20076 331372 20128 331424
rect 20444 331372 20496 331424
rect 20168 331304 20220 331356
rect 20536 331304 20588 331356
rect 20444 331236 20496 331288
rect 21916 331236 21968 331288
rect 245108 331236 245160 331288
rect 246304 331236 246356 331288
rect 299020 331236 299072 331288
rect 299296 331236 299348 331288
rect 453948 331236 454000 331288
rect 455236 331236 455288 331288
rect 482928 331236 482980 331288
rect 484216 331236 484268 331288
rect 571616 331236 571668 331288
rect 573088 331236 573140 331288
rect 192944 331168 192996 331220
rect 295432 331168 295484 331220
rect 561588 331168 561640 331220
rect 575572 331168 575624 331220
rect 576216 331168 576268 331220
rect 221924 331100 221976 331152
rect 292764 331100 292816 331152
rect 24860 330488 24912 330540
rect 145932 330488 145984 330540
rect 204168 330488 204220 330540
rect 289728 330488 289780 330540
rect 292672 330488 292724 330540
rect 299204 330488 299256 330540
rect 307668 330488 307720 330540
rect 576216 330352 576268 330404
rect 576860 330352 576912 330404
rect 15016 329740 15068 329792
rect 116952 329740 117004 329792
rect 307668 329740 307720 329792
rect 425704 329740 425756 329792
rect 426256 329740 426308 329792
rect 461032 329740 461084 329792
rect 574284 329740 574336 329792
rect 574468 329740 574520 329792
rect 575664 329740 575716 329792
rect 17500 329672 17552 329724
rect 87972 329672 88024 329724
rect 490012 329672 490064 329724
rect 15108 329604 15160 329656
rect 24860 329604 24912 329656
rect 3332 318792 3384 318844
rect 17224 318792 17276 318844
rect 437480 318112 437532 318164
rect 562324 318112 562376 318164
rect 307668 318044 307720 318096
rect 431960 318044 432012 318096
rect 578240 318044 578292 318096
rect 298744 317432 298796 317484
rect 305000 317432 305052 317484
rect 297916 317364 297968 317416
rect 307668 317364 307720 317416
rect 562324 317364 562376 317416
rect 575480 317364 575532 317416
rect 425704 316684 425756 316736
rect 565820 316684 565872 316736
rect 281448 316004 281500 316056
rect 295524 316004 295576 316056
rect 26332 315936 26384 315988
rect 139400 315936 139452 315988
rect 157340 315936 157392 315988
rect 280804 315936 280856 315988
rect 19248 315868 19300 315920
rect 93860 315868 93912 315920
rect 186228 315868 186280 315920
rect 305000 315936 305052 315988
rect 419540 315936 419592 315988
rect 448520 315936 448572 315988
rect 572904 315936 572956 315988
rect 300124 315868 300176 315920
rect 402980 315868 403032 315920
rect 482928 315868 482980 315920
rect 567108 315868 567160 315920
rect 226340 315800 226392 315852
rect 288532 315800 288584 315852
rect 296352 315800 296404 315852
rect 396080 315800 396132 315852
rect 495440 315800 495492 315852
rect 569316 315800 569368 315852
rect 231860 315732 231912 315784
rect 291568 315732 291620 315784
rect 307668 315732 307720 315784
rect 390560 315732 390612 315784
rect 500868 315732 500920 315784
rect 574652 315732 574704 315784
rect 246304 315664 246356 315716
rect 290096 315664 290148 315716
rect 302056 315664 302108 315716
rect 361580 315664 361632 315716
rect 506480 315664 506532 315716
rect 567476 315664 567528 315716
rect 298928 315596 298980 315648
rect 356060 315596 356112 315648
rect 529940 315596 529992 315648
rect 571800 315596 571852 315648
rect 14832 315392 14884 315444
rect 26332 315392 26384 315444
rect 27528 315324 27580 315376
rect 151820 315324 151872 315376
rect 285588 315324 285640 315376
rect 292948 315324 293000 315376
rect 298008 315324 298060 315376
rect 306380 315324 306432 315376
rect 307668 315324 307720 315376
rect 17592 315256 17644 315308
rect 157340 315256 157392 315308
rect 273260 315256 273312 315308
rect 297548 315256 297600 315308
rect 298100 315256 298152 315308
rect 385040 315256 385092 315308
rect 466460 315256 466512 315308
rect 571432 315256 571484 315308
rect 300124 315052 300176 315104
rect 300400 315052 300452 315104
rect 572904 314712 572956 314764
rect 576952 314712 577004 314764
rect 290096 314644 290148 314696
rect 291200 314644 291252 314696
rect 291568 314644 291620 314696
rect 292856 314644 292908 314696
rect 298928 314644 298980 314696
rect 299296 314644 299348 314696
rect 567108 314644 567160 314696
rect 568856 314644 568908 314696
rect 569316 314644 569368 314696
rect 571524 314644 571576 314696
rect 574192 314644 574244 314696
rect 574652 314644 574704 314696
rect 16396 314576 16448 314628
rect 27528 314576 27580 314628
rect 162860 314576 162912 314628
rect 285772 314576 285824 314628
rect 453948 314576 454000 314628
rect 568488 314576 568540 314628
rect 571708 314576 571760 314628
rect 285772 313896 285824 313948
rect 286968 313896 287020 313948
rect 296720 313896 296772 313948
rect 565820 313896 565872 313948
rect 575480 313896 575532 313948
rect 289728 313284 289780 313336
rect 289912 313284 289964 313336
rect 571248 313284 571300 313336
rect 571432 313284 571484 313336
rect 2780 292612 2832 292664
rect 4988 292612 5040 292664
rect 3148 266432 3200 266484
rect 6184 266432 6236 266484
rect 2780 240184 2832 240236
rect 5080 240184 5132 240236
rect 2964 213936 3016 213988
rect 6276 213936 6328 213988
rect 300400 206592 300452 206644
rect 307024 206592 307076 206644
rect 560208 206320 560260 206372
rect 571708 206320 571760 206372
rect 14924 206252 14976 206304
rect 24952 206252 25004 206304
rect 495440 206252 495492 206304
rect 575480 206252 575532 206304
rect 298008 205708 298060 205760
rect 305000 205708 305052 205760
rect 302884 205640 302936 205692
rect 310428 205640 310480 205692
rect 283288 204960 283340 205012
rect 290004 204960 290056 205012
rect 293132 204960 293184 205012
rect 540888 204960 540940 205012
rect 578240 204960 578292 205012
rect 14832 204892 14884 204944
rect 24860 204892 24912 204944
rect 289176 204892 289228 204944
rect 295524 204892 295576 204944
rect 296536 204892 296588 204944
rect 298836 204892 298888 204944
rect 374000 204892 374052 204944
rect 467104 204892 467156 204944
rect 571248 204892 571300 204944
rect 575480 204892 575532 204944
rect 292764 204756 292816 204808
rect 295340 204756 295392 204808
rect 571432 204756 571484 204808
rect 571800 204756 571852 204808
rect 17500 204688 17552 204740
rect 17684 204688 17736 204740
rect 245108 204552 245160 204604
rect 291200 204552 291252 204604
rect 291660 204552 291712 204604
rect 221924 204484 221976 204536
rect 292764 204484 292816 204536
rect 530952 204484 531004 204536
rect 571432 204484 571484 204536
rect 204168 204416 204220 204468
rect 288256 204416 288308 204468
rect 289912 204416 289964 204468
rect 299388 204416 299440 204468
rect 340880 204416 340932 204468
rect 192944 204348 192996 204400
rect 288348 204348 288400 204400
rect 295432 204348 295484 204400
rect 302056 204348 302108 204400
rect 366272 204348 366324 204400
rect 17500 204280 17552 204332
rect 87972 204280 88024 204332
rect 175188 204280 175240 204332
rect 287336 204280 287388 204332
rect 291476 204280 291528 204332
rect 304264 204280 304316 204332
rect 305000 204280 305052 204332
rect 391480 204280 391532 204332
rect 3516 204212 3568 204264
rect 30012 204212 30064 204264
rect 33140 204212 33192 204264
rect 35992 204212 36044 204264
rect 129188 204212 129240 204264
rect 134984 204212 135036 204264
rect 279884 204212 279936 204264
rect 283288 204212 283340 204264
rect 291200 204212 291252 204264
rect 292856 204212 292908 204264
rect 299204 204212 299256 204264
rect 300768 204212 300820 204264
rect 339316 204212 339368 204264
rect 340880 204212 340932 204264
rect 345112 204212 345164 204264
rect 366272 204212 366324 204264
rect 368296 204212 368348 204264
rect 408868 204212 408920 204264
rect 414664 204212 414716 204264
rect 495808 204212 495860 204264
rect 571524 204416 571576 204468
rect 513196 204348 513248 204400
rect 568764 204348 568816 204400
rect 572996 204348 573048 204400
rect 507400 204280 507452 204332
rect 567292 204280 567344 204332
rect 542176 204212 542228 204264
rect 570052 204212 570104 204264
rect 24124 204144 24176 204196
rect 25044 204144 25096 204196
rect 105360 204144 105412 204196
rect 227628 204144 227680 204196
rect 288532 204144 288584 204196
rect 300308 204144 300360 204196
rect 333520 204144 333572 204196
rect 426256 204144 426308 204196
rect 495440 204144 495492 204196
rect 524788 204144 524840 204196
rect 572904 204144 572956 204196
rect 3608 204076 3660 204128
rect 24216 204076 24268 204128
rect 24952 204076 25004 204128
rect 111156 204076 111208 204128
rect 239312 204076 239364 204128
rect 16304 204008 16356 204060
rect 99564 204008 99616 204060
rect 268292 204008 268344 204060
rect 280068 204008 280120 204060
rect 291384 204076 291436 204128
rect 291752 204076 291804 204128
rect 299020 204076 299072 204128
rect 327724 204076 327776 204128
rect 536380 204076 536432 204128
rect 568672 204076 568724 204128
rect 292764 204008 292816 204060
rect 302148 204008 302200 204060
rect 321928 204008 321980 204060
rect 432052 204008 432104 204060
rect 540888 204008 540940 204060
rect 547972 204008 548024 204060
rect 569960 204008 570012 204060
rect 19248 203940 19300 203992
rect 93952 203940 94004 203992
rect 216128 203940 216180 203992
rect 291384 203940 291436 203992
rect 300584 203940 300636 203992
rect 316132 203940 316184 203992
rect 559564 203940 559616 203992
rect 571616 203940 571668 203992
rect 21824 203872 21876 203924
rect 58992 203872 59044 203924
rect 24860 203804 24912 203856
rect 25504 203804 25556 203856
rect 140136 203804 140188 203856
rect 17776 203736 17828 203788
rect 25044 203736 25096 203788
rect 285588 203736 285640 203788
rect 295984 203736 296036 203788
rect 274088 203668 274140 203720
rect 300216 203668 300268 203720
rect 233148 203600 233200 203652
rect 291200 203600 291252 203652
rect 300124 203600 300176 203652
rect 408868 203600 408920 203652
rect 565360 203600 565412 203652
rect 572996 203600 573048 203652
rect 134984 203532 135036 203584
rect 289912 203532 289964 203584
rect 297640 203532 297692 203584
rect 478420 203532 478472 203584
rect 553768 203532 553820 203584
rect 571708 203532 571760 203584
rect 471888 202852 471940 202904
rect 472624 202852 472676 202904
rect 17868 202784 17920 202836
rect 19064 202784 19116 202836
rect 20076 202784 20128 202836
rect 22008 202784 22060 202836
rect 23388 202784 23440 202836
rect 70584 202784 70636 202836
rect 250904 202784 250956 202836
rect 291476 202784 291528 202836
rect 292948 202784 293000 202836
rect 293960 202784 294012 202836
rect 310428 202784 310480 202836
rect 426256 202784 426308 202836
rect 20352 202716 20404 202768
rect 64972 202716 65024 202768
rect 256608 202716 256660 202768
rect 287888 202716 287940 202768
rect 20444 202648 20496 202700
rect 47400 202648 47452 202700
rect 22008 202172 22060 202224
rect 53196 202172 53248 202224
rect 19064 202104 19116 202156
rect 76380 202104 76432 202156
rect 262128 202104 262180 202156
rect 292948 202104 293000 202156
rect 303712 202104 303764 202156
rect 432052 202104 432104 202156
rect 181444 201424 181496 201476
rect 292580 201424 292632 201476
rect 303528 201424 303580 201476
rect 350908 201424 350960 201476
rect 501604 201424 501656 201476
rect 574192 201424 574244 201476
rect 574468 201424 574520 201476
rect 574284 201356 574336 201408
rect 575664 201356 575716 201408
rect 490012 200744 490064 200796
rect 574284 200744 574336 200796
rect 19156 199384 19208 199436
rect 22100 199384 22152 199436
rect 122748 199384 122800 199436
rect 162860 188980 162912 189032
rect 296720 188980 296772 189032
rect 298560 188980 298612 189032
rect 396080 188980 396132 189032
rect 437480 188980 437532 189032
rect 575572 188980 575624 189032
rect 168380 188912 168432 188964
rect 276664 188912 276716 188964
rect 296444 188912 296496 188964
rect 298100 188912 298152 188964
rect 385040 188912 385092 188964
rect 442908 188912 442960 188964
rect 576860 188912 576912 188964
rect 577136 188912 577188 188964
rect 186320 188844 186372 188896
rect 289176 188844 289228 188896
rect 460940 188844 460992 188896
rect 574376 188844 574428 188896
rect 454040 188776 454092 188828
rect 560208 188776 560260 188828
rect 471888 188708 471940 188760
rect 574560 188708 574612 188760
rect 483020 188640 483072 188692
rect 568856 188640 568908 188692
rect 575572 188572 575624 188624
rect 576860 188572 576912 188624
rect 103980 188368 104032 188420
rect 162860 188368 162912 188420
rect 296260 188368 296312 188420
rect 298744 188368 298796 188420
rect 379520 188368 379572 188420
rect 560208 188368 560260 188420
rect 577044 188368 577096 188420
rect 14924 188300 14976 188352
rect 181444 188300 181496 188352
rect 307024 188300 307076 188352
rect 308036 188300 308088 188352
rect 402980 188300 403032 188352
rect 448520 188300 448572 188352
rect 575664 188300 575716 188352
rect 576952 188300 577004 188352
rect 574284 187892 574336 187944
rect 574560 187892 574612 187944
rect 568856 187688 568908 187740
rect 570144 187688 570196 187740
rect 574376 187688 574428 187740
rect 575756 187688 575808 187740
rect 300768 187620 300820 187672
rect 361580 187620 361632 187672
rect 299296 187552 299348 187604
rect 356060 187552 356112 187604
rect 13636 187076 13688 187128
rect 25504 187076 25556 187128
rect 15016 187008 15068 187060
rect 103980 187008 104032 187060
rect 296628 187008 296680 187060
rect 304264 187008 304316 187060
rect 13544 186940 13596 186992
rect 186320 186940 186372 186992
rect 298008 186940 298060 186992
rect 308036 186940 308088 186992
rect 419540 186940 419592 186992
rect 578240 186940 578292 186992
rect 288256 186872 288308 186924
rect 292856 186872 292908 186924
rect 17684 186396 17736 186448
rect 24124 186396 24176 186448
rect 19156 186328 19208 186380
rect 22100 186328 22152 186380
rect 288348 186328 288400 186380
rect 294052 186328 294104 186380
rect 276664 185852 276716 185904
rect 291568 185852 291620 185904
rect 2780 149472 2832 149524
rect 5172 149472 5224 149524
rect 3332 136688 3384 136740
rect 8944 136688 8996 136740
rect 302148 78344 302200 78396
rect 313280 78344 313332 78396
rect 300584 78276 300636 78328
rect 315948 78276 316000 78328
rect 299112 78208 299164 78260
rect 324320 78208 324372 78260
rect 471980 78208 472032 78260
rect 472992 78208 473044 78260
rect 574284 78208 574336 78260
rect 14924 78140 14976 78192
rect 82820 78140 82872 78192
rect 300492 78140 300544 78192
rect 328460 78140 328512 78192
rect 333244 78140 333296 78192
rect 454040 78140 454092 78192
rect 455328 78140 455380 78192
rect 577044 78140 577096 78192
rect 17684 78072 17736 78124
rect 111156 78072 111208 78124
rect 278780 78072 278832 78124
rect 279884 78072 279936 78124
rect 293132 78072 293184 78124
rect 300216 78072 300268 78124
rect 365720 78072 365772 78124
rect 449808 78072 449860 78124
rect 575664 78072 575716 78124
rect 13728 78004 13780 78056
rect 144920 78004 144972 78056
rect 264980 78004 265032 78056
rect 289084 78004 289136 78056
rect 290556 78004 290608 78056
rect 385040 78004 385092 78056
rect 420736 78004 420788 78056
rect 578240 78004 578292 78056
rect 14740 77936 14792 77988
rect 151912 77936 151964 77988
rect 269120 77936 269172 77988
rect 300124 77936 300176 77988
rect 310428 77936 310480 77988
rect 580448 77936 580500 77988
rect 144920 77256 144972 77308
rect 145932 77256 145984 77308
rect 419540 77256 419592 77308
rect 420276 77256 420328 77308
rect 448520 77256 448572 77308
rect 449256 77256 449308 77308
rect 75920 77052 75972 77104
rect 76702 77052 76754 77104
rect 295248 76848 295300 76900
rect 398840 76848 398892 76900
rect 390560 76780 390612 76832
rect 568948 76780 569000 76832
rect 393320 76712 393372 76764
rect 571340 76712 571392 76764
rect 295984 76644 296036 76696
rect 382280 76644 382332 76696
rect 394700 76644 394752 76696
rect 572996 76644 573048 76696
rect 266360 76576 266412 76628
rect 290464 76576 290516 76628
rect 376760 76576 376812 76628
rect 572812 76576 572864 76628
rect 13544 76508 13596 76560
rect 183468 76508 183520 76560
rect 252560 76508 252612 76560
rect 297640 76508 297692 76560
rect 299204 76508 299256 76560
rect 333244 76508 333296 76560
rect 372620 76508 372672 76560
rect 572720 76508 572772 76560
rect 19064 76032 19116 76084
rect 75920 76032 75972 76084
rect 20260 75964 20312 76016
rect 82176 75964 82228 76016
rect 82544 75964 82596 76016
rect 15016 75896 15068 75948
rect 163688 75896 163740 75948
rect 4804 75828 4856 75880
rect 30012 75828 30064 75880
rect 82820 75828 82872 75880
rect 180984 75828 181036 75880
rect 181444 75828 181496 75880
rect 183468 75828 183520 75880
rect 186504 75828 186556 75880
rect 186964 75828 187016 75880
rect 313280 75828 313332 75880
rect 321928 75828 321980 75880
rect 323584 75828 323636 75880
rect 324320 75828 324372 75880
rect 327724 75828 327776 75880
rect 333244 75828 333296 75880
rect 339316 75828 339368 75880
rect 408868 75828 408920 75880
rect 414664 75828 414716 75880
rect 467104 75828 467156 75880
rect 575480 75828 575532 75880
rect 17776 75760 17828 75812
rect 105728 75760 105780 75812
rect 129188 75760 129240 75812
rect 134524 75760 134576 75812
rect 483664 75760 483716 75812
rect 570144 75760 570196 75812
rect 16304 75692 16356 75744
rect 100208 75692 100260 75744
rect 491208 75692 491260 75744
rect 574192 75692 574244 75744
rect 19248 75624 19300 75676
rect 94044 75624 94096 75676
rect 327724 75624 327776 75676
rect 328460 75624 328512 75676
rect 496084 75624 496136 75676
rect 571524 75624 571576 75676
rect 20352 75556 20404 75608
rect 65064 75556 65116 75608
rect 65524 75556 65576 75608
rect 501604 75556 501656 75608
rect 574468 75556 574520 75608
rect 17500 75488 17552 75540
rect 88248 75488 88300 75540
rect 513196 75488 513248 75540
rect 568764 75488 568816 75540
rect 4896 75420 4948 75472
rect 24216 75420 24268 75472
rect 221924 75352 221976 75404
rect 284208 75352 284260 75404
rect 204168 75284 204220 75336
rect 221464 75284 221516 75336
rect 273260 75284 273312 75336
rect 490012 75284 490064 75336
rect 491208 75284 491260 75336
rect 210332 75216 210384 75268
rect 274548 75216 274600 75268
rect 277400 75216 277452 75268
rect 501604 75216 501656 75268
rect 59268 75148 59320 75200
rect 123484 75148 123536 75200
rect 216128 75148 216180 75200
rect 278872 75148 278924 75200
rect 280160 75148 280212 75200
rect 513196 75148 513248 75200
rect 338764 74536 338816 74588
rect 345112 74536 345164 74588
rect 19156 74468 19208 74520
rect 123024 74468 123076 74520
rect 124128 74468 124180 74520
rect 250812 74468 250864 74520
rect 291476 74468 291528 74520
rect 524788 74468 524840 74520
rect 572904 74468 572956 74520
rect 16396 74400 16448 74452
rect 116952 74400 117004 74452
rect 530584 74400 530636 74452
rect 571432 74400 571484 74452
rect 22008 74332 22060 74384
rect 53564 74332 53616 74384
rect 536104 74332 536156 74384
rect 568672 74332 568724 74384
rect 20444 74264 20496 74316
rect 47768 74264 47820 74316
rect 542176 74264 542228 74316
rect 570052 74264 570104 74316
rect 20628 74196 20680 74248
rect 41880 74196 41932 74248
rect 547880 74196 547932 74248
rect 569960 74196 570012 74248
rect 20536 74128 20588 74180
rect 36084 74128 36136 74180
rect 559564 74128 559616 74180
rect 571616 74128 571668 74180
rect 284208 74060 284260 74112
rect 287152 74060 287204 74112
rect 295340 74060 295392 74112
rect 278872 73992 278924 74044
rect 285680 73992 285732 74044
rect 291384 73992 291436 74044
rect 291476 73992 291528 74044
rect 305368 73992 305420 74044
rect 329748 73992 329800 74044
rect 374092 73992 374144 74044
rect 175188 73924 175240 73976
rect 231860 73924 231912 73976
rect 235264 73924 235316 73976
rect 274548 73924 274600 73976
rect 283840 73924 283892 73976
rect 294144 73924 294196 73976
rect 295432 73924 295484 73976
rect 530584 73924 530636 73976
rect 124128 73856 124180 73908
rect 363328 73856 363380 73908
rect 338488 73788 338540 73840
rect 378232 73788 378284 73840
rect 571708 73788 571760 73840
rect 13636 73108 13688 73160
rect 140044 73108 140096 73160
rect 245016 73108 245068 73160
rect 291660 73108 291712 73160
rect 296536 73108 296588 73160
rect 328552 73108 328604 73160
rect 329748 73108 329800 73160
rect 461032 73108 461084 73160
rect 575756 73108 575808 73160
rect 291660 72700 291712 72752
rect 303712 72700 303764 72752
rect 299296 72632 299348 72684
rect 322940 72632 322992 72684
rect 356704 72632 356756 72684
rect 169668 72564 169720 72616
rect 231308 72564 231360 72616
rect 293960 72564 294012 72616
rect 524788 72564 524840 72616
rect 94044 72496 94096 72548
rect 355048 72496 355100 72548
rect 41880 72428 41932 72480
rect 340144 72428 340196 72480
rect 461032 72292 461084 72344
rect 461584 72292 461636 72344
rect 230848 71680 230900 71732
rect 231308 71680 231360 71732
rect 287704 71680 287756 71732
rect 438124 71680 438176 71732
rect 576860 71680 576912 71732
rect 443644 71612 443696 71664
rect 577136 71612 577188 71664
rect 270592 71204 270644 71256
rect 408868 71204 408920 71256
rect 300400 71136 300452 71188
rect 547880 71136 547932 71188
rect 111708 71068 111760 71120
rect 360200 71068 360252 71120
rect 88248 71000 88300 71052
rect 353392 71000 353444 71052
rect 3056 70388 3108 70440
rect 199384 70388 199436 70440
rect 239312 70320 239364 70372
rect 292764 70320 292816 70372
rect 293500 70320 293552 70372
rect 293500 69912 293552 69964
rect 302240 69912 302292 69964
rect 298744 69844 298796 69896
rect 330208 69844 330260 69896
rect 379888 69844 379940 69896
rect 163688 69776 163740 69828
rect 229192 69776 229244 69828
rect 292120 69776 292172 69828
rect 518992 69776 519044 69828
rect 100208 69708 100260 69760
rect 356704 69708 356756 69760
rect 47768 69640 47820 69692
rect 341800 69640 341852 69692
rect 256608 68960 256660 69012
rect 290004 68960 290056 69012
rect 291108 68960 291160 69012
rect 291108 68552 291160 68604
rect 307024 68552 307076 68604
rect 298744 68484 298796 68536
rect 542176 68484 542228 68536
rect 105728 68416 105780 68468
rect 358360 68416 358412 68468
rect 82544 68348 82596 68400
rect 351920 68348 351972 68400
rect 53564 68280 53616 68332
rect 343640 68280 343692 68332
rect 267740 67532 267792 67584
rect 292580 67532 292632 67584
rect 197360 67056 197412 67108
rect 221556 67056 221608 67108
rect 292580 67056 292632 67108
rect 310520 67056 310572 67108
rect 336648 67056 336700 67108
rect 396080 67056 396132 67108
rect 134524 66988 134576 67040
rect 255688 66988 255740 67040
rect 297088 66988 297140 67040
rect 536104 66988 536156 67040
rect 116952 66920 117004 66972
rect 361672 66920 361724 66972
rect 220912 66852 220964 66904
rect 471980 66852 472032 66904
rect 215944 65628 215996 65680
rect 454040 65628 454092 65680
rect 219440 65560 219492 65612
rect 467104 65560 467156 65612
rect 202880 65492 202932 65544
rect 559564 65492 559616 65544
rect 302332 64812 302384 64864
rect 431960 64812 432012 64864
rect 209320 64336 209372 64388
rect 302332 64336 302384 64388
rect 272524 64268 272576 64320
rect 477500 64268 477552 64320
rect 212632 64200 212684 64252
rect 443644 64200 443696 64252
rect 8944 64132 8996 64184
rect 57612 64132 57664 64184
rect 217600 64132 217652 64184
rect 461584 64132 461636 64184
rect 123484 62976 123536 63028
rect 345112 62976 345164 63028
rect 75920 62908 75972 62960
rect 350080 62908 350132 62960
rect 71044 62840 71096 62892
rect 348424 62840 348476 62892
rect 65524 62772 65576 62824
rect 346768 62772 346820 62824
rect 379888 62772 379940 62824
rect 553400 62772 553452 62824
rect 226340 62024 226392 62076
rect 288532 62024 288584 62076
rect 288808 62024 288860 62076
rect 303804 62024 303856 62076
rect 425060 62024 425112 62076
rect 186964 61548 187016 61600
rect 236000 61548 236052 61600
rect 315304 61548 315356 61600
rect 323584 61548 323636 61600
rect 144920 61480 144972 61532
rect 221740 61480 221792 61532
rect 300768 61480 300820 61532
rect 325240 61480 325292 61532
rect 361580 61480 361632 61532
rect 140044 61412 140096 61464
rect 222568 61412 222620 61464
rect 284300 61412 284352 61464
rect 381544 61412 381596 61464
rect 222108 61344 222160 61396
rect 438124 61344 438176 61396
rect 318800 60324 318852 60376
rect 333244 60324 333296 60376
rect 321928 60256 321980 60308
rect 350540 60256 350592 60308
rect 191840 60188 191892 60240
rect 237380 60188 237432 60240
rect 273352 60188 273404 60240
rect 320088 60188 320140 60240
rect 181444 60120 181496 60172
rect 234160 60120 234212 60172
rect 242440 60120 242492 60172
rect 289820 60120 289872 60172
rect 296444 60120 296496 60172
rect 331864 60188 331916 60240
rect 385132 60188 385184 60240
rect 332968 60120 333020 60172
rect 390652 60120 390704 60172
rect 221464 60052 221516 60104
rect 282184 60052 282236 60104
rect 292856 60052 292908 60104
rect 294604 60052 294656 60104
rect 371608 60052 371660 60104
rect 206008 59984 206060 60036
rect 419540 59984 419592 60036
rect 237380 59304 237432 59356
rect 294052 59304 294104 59356
rect 296628 59304 296680 59356
rect 332968 59304 333020 59356
rect 333520 59304 333572 59356
rect 260840 59236 260892 59288
rect 292580 59236 292632 59288
rect 292948 59236 293000 59288
rect 316960 58896 317012 58948
rect 327724 58896 327776 58948
rect 220728 58828 220780 58880
rect 278780 58828 278832 58880
rect 320824 58828 320876 58880
rect 338764 58828 338816 58880
rect 157984 58760 158036 58812
rect 227720 58760 227772 58812
rect 298008 58760 298060 58812
rect 336832 58760 336884 58812
rect 402980 58760 403032 58812
rect 151820 58692 151872 58744
rect 225880 58692 225932 58744
rect 231952 58692 232004 58744
rect 261576 58692 261628 58744
rect 328368 58692 328420 58744
rect 367100 58692 367152 58744
rect 396448 58692 396500 58744
rect 564440 58692 564492 58744
rect 214288 58624 214340 58676
rect 448520 58624 448572 58676
rect 102140 57944 102192 57996
rect 104164 57944 104216 57996
rect 221740 57876 221792 57928
rect 224592 57876 224644 57928
rect 299388 57876 299440 57928
rect 320824 57876 320876 57928
rect 261576 57604 261628 57656
rect 291108 57604 291160 57656
rect 259368 57536 259420 57588
rect 288440 57536 288492 57588
rect 292580 57536 292632 57588
rect 309048 57536 309100 57588
rect 320088 57536 320140 57588
rect 365352 57536 365404 57588
rect 251088 57468 251140 57520
rect 297456 57468 297508 57520
rect 297548 57468 297600 57520
rect 368664 57468 368716 57520
rect 257712 57400 257764 57452
rect 289912 57400 289964 57452
rect 294696 57400 294748 57452
rect 370320 57400 370372 57452
rect 211344 57332 211396 57384
rect 222108 57332 222160 57384
rect 272616 57332 272668 57384
rect 483664 57332 483716 57384
rect 208032 57264 208084 57316
rect 218060 57264 218112 57316
rect 275928 57264 275980 57316
rect 496084 57264 496136 57316
rect 204720 57196 204772 57248
rect 220728 57196 220780 57248
rect 221556 57196 221608 57248
rect 239496 57196 239548 57248
rect 254400 57196 254452 57248
rect 272524 57196 272576 57248
rect 279240 57196 279292 57248
rect 507124 57196 507176 57248
rect 312360 56584 312412 56636
rect 316040 56584 316092 56636
rect 5172 56516 5224 56568
rect 57520 56516 57572 56568
rect 102140 53796 102192 53848
rect 109040 53796 109092 53848
rect 102140 52640 102192 52692
rect 103888 52640 103940 52692
rect 102140 52436 102192 52488
rect 196164 52436 196216 52488
rect 5080 52368 5132 52420
rect 57060 52368 57112 52420
rect 102784 52368 102836 52420
rect 195980 52368 196032 52420
rect 102876 52300 102928 52352
rect 196072 52300 196124 52352
rect 102968 51008 103020 51060
rect 195980 51008 196032 51060
rect 102140 49784 102192 49836
rect 104440 49784 104492 49836
rect 102600 49648 102652 49700
rect 196072 49648 196124 49700
rect 104164 49580 104216 49632
rect 195980 49580 196032 49632
rect 102140 48832 102192 48884
rect 104348 48832 104400 48884
rect 103060 48220 103112 48272
rect 195980 48220 196032 48272
rect 109040 48152 109092 48204
rect 196072 48152 196124 48204
rect 6184 46860 6236 46912
rect 57520 46860 57572 46912
rect 103888 46860 103940 46912
rect 195980 46860 196032 46912
rect 103244 45500 103296 45552
rect 195980 45500 196032 45552
rect 104440 44820 104492 44872
rect 196072 44820 196124 44872
rect 3332 44140 3384 44192
rect 60004 44140 60056 44192
rect 104348 44072 104400 44124
rect 195980 44072 196032 44124
rect 3516 42712 3568 42764
rect 57152 42712 57204 42764
rect 102968 42712 103020 42764
rect 195980 42712 196032 42764
rect 102600 42644 102652 42696
rect 196072 42644 196124 42696
rect 102876 41352 102928 41404
rect 195980 41352 196032 41404
rect 102140 40672 102192 40724
rect 196164 40672 196216 40724
rect 102324 39992 102376 40044
rect 196072 39992 196124 40044
rect 103520 39924 103572 39976
rect 195980 39924 196032 39976
rect 102232 38564 102284 38616
rect 195980 38564 196032 38616
rect 6276 37204 6328 37256
rect 57060 37204 57112 37256
rect 102140 37204 102192 37256
rect 195980 37204 196032 37256
rect 102784 35844 102836 35896
rect 195980 35844 196032 35896
rect 102692 35776 102744 35828
rect 196072 35776 196124 35828
rect 102876 34416 102928 34468
rect 195980 34416 196032 34468
rect 102600 34348 102652 34400
rect 196072 34348 196124 34400
rect 102140 33056 102192 33108
rect 195980 33056 196032 33108
rect 4988 31696 5040 31748
rect 57612 31696 57664 31748
rect 102324 31696 102376 31748
rect 195980 31696 196032 31748
rect 102140 31628 102192 31680
rect 196072 31628 196124 31680
rect 102232 30268 102284 30320
rect 195980 30268 196032 30320
rect 102140 30200 102192 30252
rect 196072 30200 196124 30252
rect 102140 28908 102192 28960
rect 195980 28908 196032 28960
rect 102140 28228 102192 28280
rect 195980 28228 196032 28280
rect 17224 27548 17276 27600
rect 57244 27548 57296 27600
rect 102140 27548 102192 27600
rect 195980 27548 196032 27600
rect 102784 26188 102836 26240
rect 195980 26188 196032 26240
rect 18604 24216 18656 24268
rect 356980 24216 357032 24268
rect 7564 24148 7616 24200
rect 364432 24148 364484 24200
rect 382832 24148 382884 24200
rect 398840 24148 398892 24200
rect 16488 24080 16540 24132
rect 375012 24080 375064 24132
rect 393320 24080 393372 24132
rect 569224 24080 569276 24132
rect 85488 23468 85540 23520
rect 266360 23468 266412 23520
rect 267372 23468 267424 23520
rect 60004 22244 60056 22296
rect 353760 22244 353812 22296
rect 3516 22176 3568 22228
rect 335820 22176 335872 22228
rect 3608 22108 3660 22160
rect 346584 22108 346636 22160
rect 62304 22040 62356 22092
rect 85488 22040 85540 22092
rect 199384 22040 199436 22092
rect 350172 22040 350224 22092
rect 386052 22040 386104 22092
rect 574100 22040 574152 22092
rect 3424 21972 3476 22024
rect 371700 21972 371752 22024
rect 396816 21972 396868 22024
rect 570604 21972 570656 22024
rect 18696 21904 18748 21956
rect 360936 21904 360988 21956
rect 378876 21904 378928 21956
rect 400220 21904 400272 21956
rect 175464 21496 175516 21548
rect 285588 21496 285640 21548
rect 187700 21428 187752 21480
rect 299940 21428 299992 21480
rect 152464 21360 152516 21412
rect 292764 21360 292816 21412
rect 178040 20068 178092 20120
rect 256884 20068 256936 20120
rect 162860 20000 162912 20052
rect 307116 20000 307168 20052
rect 138020 19932 138072 19984
rect 282000 19932 282052 19984
rect 155960 18776 156012 18828
rect 187700 18776 187752 18828
rect 175280 18708 175332 18760
rect 253296 18708 253348 18760
rect 150440 18640 150492 18692
rect 228180 18640 228232 18692
rect 142160 18572 142212 18624
rect 175464 18572 175516 18624
rect 184940 18572 184992 18624
rect 328644 18572 328696 18624
rect 171140 17348 171192 17400
rect 249708 17348 249760 17400
rect 131120 17280 131172 17332
rect 274824 17280 274876 17332
rect 71136 17212 71188 17264
rect 242900 17212 242952 17264
rect 168380 15988 168432 16040
rect 245660 15988 245712 16040
rect 135260 15920 135312 15972
rect 277400 15920 277452 15972
rect 74540 15852 74592 15904
rect 245936 15852 245988 15904
rect 136456 14560 136508 14612
rect 212540 14560 212592 14612
rect 164424 14492 164476 14544
rect 241520 14492 241572 14544
rect 170312 14424 170364 14476
rect 313280 14424 313332 14476
rect 139584 13200 139636 13252
rect 216680 13200 216732 13252
rect 160100 13132 160152 13184
rect 238760 13132 238812 13184
rect 176660 13064 176712 13116
rect 320180 13064 320232 13116
rect 153752 11908 153804 11960
rect 230480 11908 230532 11960
rect 125600 11840 125652 11892
rect 202880 11840 202932 11892
rect 186136 11772 186188 11824
rect 263600 11772 263652 11824
rect 151820 11704 151872 11756
rect 295340 11704 295392 11756
rect 156604 10412 156656 10464
rect 209780 10412 209832 10464
rect 147128 10344 147180 10396
rect 223580 10344 223632 10396
rect 3424 10276 3476 10328
rect 338120 10276 338172 10328
rect 174268 9052 174320 9104
rect 317420 9052 317472 9104
rect 167184 8984 167236 9036
rect 310520 8984 310572 9036
rect 84200 8916 84252 8968
rect 241704 8916 241756 8968
rect 157800 7692 157852 7744
rect 234620 7692 234672 7744
rect 235908 7692 235960 7744
rect 288440 7692 288492 7744
rect 128176 7624 128228 7676
rect 270500 7624 270552 7676
rect 88340 7556 88392 7608
rect 245200 7556 245252 7608
rect 143540 6332 143592 6384
rect 220820 6332 220872 6384
rect 181444 6264 181496 6316
rect 324320 6264 324372 6316
rect 92480 6196 92532 6248
rect 248788 6196 248840 6248
rect 78680 6128 78732 6180
rect 249984 6128 250036 6180
rect 182548 4972 182600 5024
rect 259460 4972 259512 5024
rect 129372 4904 129424 4956
rect 205640 4904 205692 4956
rect 188528 4836 188580 4888
rect 331220 4836 331272 4888
rect 96620 4768 96672 4820
rect 252376 4768 252428 4820
rect 149520 3816 149572 3868
rect 152464 3816 152516 3868
rect 145932 3544 145984 3596
rect 235908 3544 235960 3596
rect 132960 3476 133012 3528
rect 156604 3476 156656 3528
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 161388 3476 161440 3528
rect 302240 3476 302292 3528
rect 66260 3408 66312 3460
rect 239312 3408 239364 3460
rect 266360 3408 266412 3460
rect 579804 3408 579856 3460
rect 151820 3340 151872 3392
rect 153016 3340 153068 3392
rect 176660 3340 176712 3392
rect 177856 3340 177908 3392
rect 160100 2796 160152 2848
rect 161388 2796 161440 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700534 8156 703520
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 16488 700528 16540 700534
rect 16488 700470 16540 700476
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 671090 3464 671191
rect 3424 671084 3476 671090
rect 3424 671026 3476 671032
rect 7656 671084 7708 671090
rect 7656 671026 7708 671032
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 607209 2820 658135
rect 2870 619168 2926 619177
rect 2870 619103 2926 619112
rect 2884 618934 2912 619103
rect 2872 618928 2924 618934
rect 2872 618870 2924 618876
rect 4988 618928 5040 618934
rect 4988 618870 5040 618876
rect 2778 607200 2834 607209
rect 2778 607135 2834 607144
rect 3422 607200 3478 607209
rect 3422 607135 3478 607144
rect 3436 606121 3464 607135
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 2778 462632 2834 462641
rect 2778 462567 2834 462576
rect 2792 462466 2820 462567
rect 2780 462460 2832 462466
rect 2780 462402 2832 462408
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 398750 2820 449511
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409970 2912 410479
rect 2872 409964 2924 409970
rect 2872 409906 2924 409912
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292670 2820 293111
rect 2780 292664 2832 292670
rect 2780 292606 2832 292612
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3160 266490 3188 267135
rect 3148 266484 3200 266490
rect 3148 266426 3200 266432
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 2962 214976 3018 214985
rect 2962 214911 3018 214920
rect 2976 213994 3004 214911
rect 2964 213988 3016 213994
rect 2964 213930 3016 213936
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 2792 149530 2820 149767
rect 2780 149524 2832 149530
rect 2780 149466 2832 149472
rect 3330 136776 3386 136785
rect 3330 136711 3332 136720
rect 3384 136711 3386 136720
rect 3332 136682 3384 136688
rect 3054 71632 3110 71641
rect 3054 71567 3110 71576
rect 3068 70446 3096 71567
rect 3056 70440 3108 70446
rect 3056 70382 3108 70388
rect 3330 45520 3386 45529
rect 3330 45455 3386 45464
rect 3344 44198 3372 45455
rect 3332 44192 3384 44198
rect 3332 44134 3384 44140
rect 3436 22030 3464 606047
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 204270 3556 566879
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3516 204264 3568 204270
rect 3516 204206 3568 204212
rect 3620 204134 3648 514791
rect 3712 502489 3740 553823
rect 3698 502480 3754 502489
rect 3698 502415 3754 502424
rect 3712 501809 3740 502415
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 4804 462460 4856 462466
rect 4804 462402 4856 462408
rect 3608 204128 3660 204134
rect 3608 204070 3660 204076
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3528 42770 3556 188799
rect 3606 84688 3662 84697
rect 3606 84623 3662 84632
rect 3516 42764 3568 42770
rect 3516 42706 3568 42712
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3528 22234 3556 32399
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3620 22166 3648 84623
rect 4816 75886 4844 462402
rect 4896 409964 4948 409970
rect 4896 409906 4948 409912
rect 4804 75880 4856 75886
rect 4804 75822 4856 75828
rect 4908 75478 4936 409906
rect 5000 332722 5028 618870
rect 7564 398744 7616 398750
rect 7564 398686 7616 398692
rect 4988 332716 5040 332722
rect 4988 332658 5040 332664
rect 4988 292664 5040 292670
rect 4988 292606 5040 292612
rect 4896 75472 4948 75478
rect 4896 75414 4948 75420
rect 5000 31754 5028 292606
rect 6184 266484 6236 266490
rect 6184 266426 6236 266432
rect 5080 240236 5132 240242
rect 5080 240178 5132 240184
rect 5092 52426 5120 240178
rect 5172 149524 5224 149530
rect 5172 149466 5224 149472
rect 5184 56574 5212 149466
rect 5172 56568 5224 56574
rect 5172 56510 5224 56516
rect 5080 52420 5132 52426
rect 5080 52362 5132 52368
rect 6196 46918 6224 266426
rect 6276 213988 6328 213994
rect 6276 213930 6328 213936
rect 6184 46912 6236 46918
rect 6184 46854 6236 46860
rect 6288 37262 6316 213930
rect 6276 37256 6328 37262
rect 6276 37198 6328 37204
rect 4988 31748 5040 31754
rect 4988 31690 5040 31696
rect 7576 24206 7604 398686
rect 7668 332586 7696 671026
rect 15016 583228 15068 583234
rect 15016 583170 15068 583176
rect 14924 580304 14976 580310
rect 14924 580246 14976 580252
rect 14832 462324 14884 462330
rect 14832 462266 14884 462272
rect 14844 461038 14872 462266
rect 14832 461032 14884 461038
rect 14832 460974 14884 460980
rect 14844 345014 14872 460974
rect 14936 460902 14964 580246
rect 15028 462330 15056 583170
rect 15108 583092 15160 583098
rect 15108 583034 15160 583040
rect 15016 462324 15068 462330
rect 15016 462266 15068 462272
rect 15120 461650 15148 583034
rect 16396 583024 16448 583030
rect 16396 582966 16448 582972
rect 16408 462330 16436 582966
rect 16396 462324 16448 462330
rect 16396 462266 16448 462272
rect 15108 461644 15160 461650
rect 15108 461586 15160 461592
rect 14924 460896 14976 460902
rect 14924 460838 14976 460844
rect 14936 459762 14964 460838
rect 14936 459734 15148 459762
rect 15016 459672 15068 459678
rect 15016 459614 15068 459620
rect 14844 344986 14964 345014
rect 14936 334014 14964 344986
rect 14924 334008 14976 334014
rect 14924 333950 14976 333956
rect 7656 332580 7708 332586
rect 7656 332522 7708 332528
rect 14832 315444 14884 315450
rect 14832 315386 14884 315392
rect 14738 207768 14794 207777
rect 14738 207703 14794 207712
rect 13726 207632 13782 207641
rect 13726 207567 13782 207576
rect 13636 187128 13688 187134
rect 13636 187070 13688 187076
rect 13544 186992 13596 186998
rect 13544 186934 13596 186940
rect 8944 136740 8996 136746
rect 8944 136682 8996 136688
rect 8956 64190 8984 136682
rect 13556 76566 13584 186934
rect 13544 76560 13596 76566
rect 13544 76502 13596 76508
rect 13648 73166 13676 187070
rect 13740 78062 13768 207567
rect 13728 78056 13780 78062
rect 13728 77998 13780 78004
rect 14752 77994 14780 207703
rect 14844 204950 14872 315386
rect 14936 206310 14964 333950
rect 15028 329798 15056 459614
rect 15016 329792 15068 329798
rect 15016 329734 15068 329740
rect 14924 206304 14976 206310
rect 14924 206246 14976 206252
rect 14832 204944 14884 204950
rect 14832 204886 14884 204892
rect 15028 203561 15056 329734
rect 15120 329662 15148 459734
rect 16304 459604 16356 459610
rect 16304 459546 16356 459552
rect 16316 332790 16344 459546
rect 16304 332784 16356 332790
rect 16304 332726 16356 332732
rect 15108 329656 15160 329662
rect 15108 329598 15160 329604
rect 15120 207641 15148 329598
rect 15106 207632 15162 207641
rect 15106 207567 15162 207576
rect 16316 204066 16344 332726
rect 16408 314634 16436 462266
rect 16396 314628 16448 314634
rect 16396 314570 16448 314576
rect 16408 207777 16436 314570
rect 16394 207768 16450 207777
rect 16394 207703 16450 207712
rect 16304 204060 16356 204066
rect 16304 204002 16356 204008
rect 15014 203552 15070 203561
rect 15014 203487 15070 203496
rect 14924 188352 14976 188358
rect 14924 188294 14976 188300
rect 14936 78198 14964 188294
rect 15016 187060 15068 187066
rect 15016 187002 15068 187008
rect 14924 78192 14976 78198
rect 14924 78134 14976 78140
rect 14740 77988 14792 77994
rect 14740 77930 14792 77936
rect 15028 75954 15056 187002
rect 15016 75948 15068 75954
rect 15016 75890 15068 75896
rect 16316 75750 16344 204002
rect 16394 203552 16450 203561
rect 16394 203487 16450 203496
rect 16304 75744 16356 75750
rect 16304 75686 16356 75692
rect 16408 74458 16436 203487
rect 16396 74452 16448 74458
rect 16396 74394 16448 74400
rect 13636 73160 13688 73166
rect 13636 73102 13688 73108
rect 8944 64184 8996 64190
rect 8944 64126 8996 64132
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 16500 24138 16528 700470
rect 20628 700460 20680 700466
rect 20628 700402 20680 700408
rect 20444 700392 20496 700398
rect 20444 700334 20496 700340
rect 20352 700324 20404 700330
rect 20352 700266 20404 700272
rect 20364 586430 20392 700266
rect 20456 586498 20484 700334
rect 20536 699712 20588 699718
rect 20536 699654 20588 699660
rect 20444 586492 20496 586498
rect 20444 586434 20496 586440
rect 20352 586424 20404 586430
rect 20352 586366 20404 586372
rect 20444 586084 20496 586090
rect 20444 586026 20496 586032
rect 17868 586016 17920 586022
rect 17868 585958 17920 585964
rect 19246 585984 19302 585993
rect 17684 583432 17736 583438
rect 17684 583374 17736 583380
rect 17592 572076 17644 572082
rect 17592 572018 17644 572024
rect 17408 461644 17460 461650
rect 17408 461586 17460 461592
rect 17420 333266 17448 461586
rect 17604 459202 17632 572018
rect 17592 459196 17644 459202
rect 17592 459138 17644 459144
rect 17500 458244 17552 458250
rect 17500 458186 17552 458192
rect 17408 333260 17460 333266
rect 17408 333202 17460 333208
rect 17512 329730 17540 458186
rect 17604 332654 17632 459138
rect 17696 458046 17724 583374
rect 17776 583364 17828 583370
rect 17776 583306 17828 583312
rect 17788 459338 17816 583306
rect 17776 459332 17828 459338
rect 17776 459274 17828 459280
rect 17788 458250 17816 459274
rect 17776 458244 17828 458250
rect 17776 458186 17828 458192
rect 17684 458040 17736 458046
rect 17684 457982 17736 457988
rect 17696 345014 17724 457982
rect 17880 456074 17908 585958
rect 19246 585919 19302 585928
rect 20352 585948 20404 585954
rect 19156 583296 19208 583302
rect 19156 583238 19208 583244
rect 19064 583160 19116 583166
rect 19064 583102 19116 583108
rect 18604 572144 18656 572150
rect 18604 572086 18656 572092
rect 18616 459610 18644 572086
rect 18696 572008 18748 572014
rect 18696 571950 18748 571956
rect 18708 459678 18736 571950
rect 19076 463418 19104 583102
rect 19064 463412 19116 463418
rect 19064 463354 19116 463360
rect 18696 459672 18748 459678
rect 18696 459614 18748 459620
rect 18604 459604 18656 459610
rect 18604 459546 18656 459552
rect 18616 459406 18644 459546
rect 18604 459400 18656 459406
rect 18604 459342 18656 459348
rect 18708 459270 18736 459614
rect 18696 459264 18748 459270
rect 18696 459206 18748 459212
rect 19168 458114 19196 583238
rect 19260 458726 19288 585919
rect 20352 585890 20404 585896
rect 20260 585812 20312 585818
rect 20260 585754 20312 585760
rect 20272 459610 20300 585754
rect 20260 459604 20312 459610
rect 20260 459546 20312 459552
rect 19248 458720 19300 458726
rect 19248 458662 19300 458668
rect 19156 458108 19208 458114
rect 19156 458050 19208 458056
rect 19168 456770 19196 458050
rect 19168 456742 19288 456770
rect 17868 456068 17920 456074
rect 17868 456010 17920 456016
rect 19156 456068 19208 456074
rect 19156 456010 19208 456016
rect 19064 443420 19116 443426
rect 19064 443362 19116 443368
rect 18604 357468 18656 357474
rect 18604 357410 18656 357416
rect 17696 344986 17908 345014
rect 17592 332648 17644 332654
rect 17592 332590 17644 332596
rect 17604 331242 17632 332590
rect 17880 332489 17908 344986
rect 17866 332480 17922 332489
rect 17866 332415 17922 332424
rect 17604 331214 17816 331242
rect 17500 329724 17552 329730
rect 17500 329666 17552 329672
rect 17512 325694 17540 329666
rect 17512 325666 17724 325694
rect 17224 318844 17276 318850
rect 17224 318786 17276 318792
rect 17236 27606 17264 318786
rect 17592 315308 17644 315314
rect 17592 315250 17644 315256
rect 17500 204740 17552 204746
rect 17500 204682 17552 204688
rect 17512 204338 17540 204682
rect 17500 204332 17552 204338
rect 17500 204274 17552 204280
rect 17512 75546 17540 204274
rect 17604 200025 17632 315250
rect 17696 204746 17724 325666
rect 17684 204740 17736 204746
rect 17684 204682 17736 204688
rect 17788 203794 17816 331214
rect 17776 203788 17828 203794
rect 17776 203730 17828 203736
rect 17590 200016 17646 200025
rect 17590 199951 17646 199960
rect 17684 186448 17736 186454
rect 17684 186390 17736 186396
rect 17696 78130 17724 186390
rect 17684 78124 17736 78130
rect 17684 78066 17736 78072
rect 17788 75818 17816 203730
rect 17880 202842 17908 332415
rect 17868 202836 17920 202842
rect 17868 202778 17920 202784
rect 17776 75812 17828 75818
rect 17776 75754 17828 75760
rect 17500 75540 17552 75546
rect 17500 75482 17552 75488
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 18616 24274 18644 357410
rect 18696 345092 18748 345098
rect 18696 345034 18748 345040
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 16488 24132 16540 24138
rect 16488 24074 16540 24080
rect 3608 22160 3660 22166
rect 3608 22102 3660 22108
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 18708 21962 18736 345034
rect 19076 332926 19104 443362
rect 19168 333334 19196 456010
rect 19156 333328 19208 333334
rect 19156 333270 19208 333276
rect 19064 332920 19116 332926
rect 19064 332862 19116 332868
rect 19076 325694 19104 332862
rect 19076 325666 19196 325694
rect 19064 202836 19116 202842
rect 19064 202778 19116 202784
rect 19076 202162 19104 202778
rect 19064 202156 19116 202162
rect 19064 202098 19116 202104
rect 19076 76090 19104 202098
rect 19168 199442 19196 325666
rect 19260 315926 19288 456742
rect 20272 332314 20300 459546
rect 20364 458969 20392 585890
rect 20350 458960 20406 458969
rect 20350 458895 20406 458904
rect 20260 332308 20312 332314
rect 20260 332250 20312 332256
rect 20076 331424 20128 331430
rect 20076 331366 20128 331372
rect 19248 315920 19300 315926
rect 19248 315862 19300 315868
rect 19260 203998 19288 315862
rect 19248 203992 19300 203998
rect 19248 203934 19300 203940
rect 19156 199436 19208 199442
rect 19156 199378 19208 199384
rect 19156 186380 19208 186386
rect 19156 186322 19208 186328
rect 19064 76084 19116 76090
rect 19064 76026 19116 76032
rect 19168 74526 19196 186322
rect 19260 75682 19288 203934
rect 20088 202842 20116 331366
rect 20168 331356 20220 331362
rect 20168 331298 20220 331304
rect 20180 203946 20208 331298
rect 20272 204105 20300 332250
rect 20364 332246 20392 458895
rect 20456 457978 20484 586026
rect 20548 462262 20576 699654
rect 20536 462256 20588 462262
rect 20536 462198 20588 462204
rect 20640 459542 20668 700402
rect 24320 699718 24348 703520
rect 72988 700534 73016 703520
rect 72976 700528 73028 700534
rect 72976 700470 73028 700476
rect 89180 700466 89208 703520
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 154132 700398 154160 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 154120 700392 154172 700398
rect 202800 700369 202828 700946
rect 154120 700334 154172 700340
rect 202786 700360 202842 700369
rect 218992 700330 219020 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 397472 700534 397500 700946
rect 295248 700528 295300 700534
rect 295248 700470 295300 700476
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 202786 700295 202842 700304
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24228 587302 24564 587330
rect 30024 587302 30360 587330
rect 35912 587302 36156 587330
rect 41616 587302 41952 587330
rect 47412 587302 47748 587330
rect 53208 587302 53544 587330
rect 59004 587302 59340 587330
rect 64892 587302 65136 587330
rect 70596 587302 70932 587330
rect 76392 587302 76728 587330
rect 82188 587302 82524 587330
rect 87984 587302 88320 587330
rect 93872 587302 94116 587330
rect 99576 587302 99912 587330
rect 105372 587302 105708 587330
rect 111168 587302 111504 587330
rect 116964 587302 117300 587330
rect 122852 587302 123096 587330
rect 128892 587302 129228 587330
rect 24228 586498 24256 587302
rect 24216 586492 24268 586498
rect 24216 586434 24268 586440
rect 30024 586430 30052 587302
rect 30012 586424 30064 586430
rect 30012 586366 30064 586372
rect 22008 586152 22060 586158
rect 22008 586094 22060 586100
rect 22020 460934 22048 586094
rect 35912 585954 35940 587302
rect 35900 585948 35952 585954
rect 35900 585890 35952 585896
rect 37924 585948 37976 585954
rect 37924 585890 37976 585896
rect 31024 585880 31076 585886
rect 31024 585822 31076 585828
rect 31036 572150 31064 585822
rect 31024 572144 31076 572150
rect 31024 572086 31076 572092
rect 37936 572082 37964 585890
rect 41616 585818 41644 587302
rect 47412 586158 47440 587302
rect 47400 586152 47452 586158
rect 47400 586094 47452 586100
rect 53208 586090 53236 587302
rect 53196 586084 53248 586090
rect 53196 586026 53248 586032
rect 59004 586022 59032 587302
rect 58992 586016 59044 586022
rect 64892 585993 64920 587302
rect 58992 585958 59044 585964
rect 64878 585984 64934 585993
rect 64878 585919 64934 585928
rect 70596 585857 70624 587302
rect 70582 585848 70638 585857
rect 41604 585812 41656 585818
rect 41604 585754 41656 585760
rect 43444 585812 43496 585818
rect 70582 585783 70638 585792
rect 43444 585754 43496 585760
rect 37924 572076 37976 572082
rect 37924 572018 37976 572024
rect 43456 572014 43484 585754
rect 76392 583438 76420 587302
rect 82188 585721 82216 587302
rect 82174 585712 82230 585721
rect 82174 585647 82230 585656
rect 76380 583432 76432 583438
rect 76380 583374 76432 583380
rect 87984 583370 88012 587302
rect 87972 583364 88024 583370
rect 87972 583306 88024 583312
rect 93872 583302 93900 587302
rect 99576 585886 99604 587302
rect 105372 585954 105400 587302
rect 105360 585948 105412 585954
rect 105360 585890 105412 585896
rect 99564 585880 99616 585886
rect 99564 585822 99616 585828
rect 93860 583296 93912 583302
rect 93860 583238 93912 583244
rect 111168 583234 111196 587302
rect 116964 585818 116992 587302
rect 116952 585812 117004 585818
rect 116952 585754 117004 585760
rect 111156 583228 111208 583234
rect 111156 583170 111208 583176
rect 122852 583166 122880 587302
rect 129200 586498 129228 587302
rect 134352 587302 134688 587330
rect 140148 587302 140484 587330
rect 145944 587302 146280 587330
rect 151832 587302 152076 587330
rect 157872 587302 158208 587330
rect 163668 587302 164004 587330
rect 134352 586498 134380 587302
rect 129188 586492 129240 586498
rect 129188 586434 129240 586440
rect 134340 586492 134392 586498
rect 134340 586434 134392 586440
rect 134352 585721 134380 586434
rect 134338 585712 134394 585721
rect 134338 585647 134394 585656
rect 122840 583160 122892 583166
rect 122840 583102 122892 583108
rect 140148 583098 140176 587302
rect 140136 583092 140188 583098
rect 140136 583034 140188 583040
rect 145944 580310 145972 587302
rect 151832 583030 151860 587302
rect 151820 583024 151872 583030
rect 151820 582966 151872 582972
rect 158180 580378 158208 587302
rect 158168 580372 158220 580378
rect 158168 580314 158220 580320
rect 163976 580310 164004 587302
rect 168392 587302 169464 587330
rect 175200 587302 175260 587330
rect 181056 587302 181392 587330
rect 145932 580304 145984 580310
rect 145932 580246 145984 580252
rect 163964 580304 164016 580310
rect 163964 580246 164016 580252
rect 168392 572014 168420 587302
rect 175200 583030 175228 587302
rect 175188 583024 175240 583030
rect 175188 582966 175240 582972
rect 181364 580446 181392 587302
rect 186332 587302 186852 587330
rect 192648 587302 192984 587330
rect 198444 587302 198688 587330
rect 181352 580440 181404 580446
rect 181352 580382 181404 580388
rect 186332 572082 186360 587302
rect 192956 583098 192984 587302
rect 198660 586498 198688 587302
rect 204180 587302 204240 587330
rect 210036 587302 210372 587330
rect 215832 587302 216168 587330
rect 221628 587302 221964 587330
rect 227424 587302 227668 587330
rect 198648 586492 198700 586498
rect 198648 586434 198700 586440
rect 204180 583166 204208 587302
rect 210344 583234 210372 587302
rect 216140 583302 216168 587302
rect 221936 583370 221964 587302
rect 227640 585857 227668 587302
rect 233160 587302 233220 587330
rect 239016 587302 239352 587330
rect 227626 585848 227682 585857
rect 227626 585783 227682 585792
rect 233160 583438 233188 587302
rect 239324 585993 239352 587302
rect 244292 587302 244812 587330
rect 250608 587302 250944 587330
rect 256404 587302 256648 587330
rect 239310 585984 239366 585993
rect 239310 585919 239366 585928
rect 233148 583432 233200 583438
rect 233148 583374 233200 583380
rect 221924 583364 221976 583370
rect 221924 583306 221976 583312
rect 216128 583296 216180 583302
rect 216128 583238 216180 583244
rect 210332 583228 210384 583234
rect 210332 583170 210384 583176
rect 204168 583160 204220 583166
rect 204168 583102 204220 583108
rect 192944 583092 192996 583098
rect 192944 583034 192996 583040
rect 244292 572150 244320 587302
rect 250916 585818 250944 587302
rect 256620 585886 256648 587302
rect 262140 587302 262200 587330
rect 267996 587302 268332 587330
rect 262140 585954 262168 587302
rect 268304 586022 268332 587302
rect 273272 587302 273792 587330
rect 279588 587302 279924 587330
rect 268292 586016 268344 586022
rect 268292 585958 268344 585964
rect 262128 585948 262180 585954
rect 262128 585890 262180 585896
rect 256608 585880 256660 585886
rect 256608 585822 256660 585828
rect 250904 585812 250956 585818
rect 250904 585754 250956 585760
rect 273272 572218 273300 587302
rect 279896 586090 279924 587302
rect 284312 587302 285384 587330
rect 279884 586084 279936 586090
rect 279884 586026 279936 586032
rect 273260 572212 273312 572218
rect 273260 572154 273312 572160
rect 244280 572144 244332 572150
rect 244280 572086 244332 572092
rect 186320 572076 186372 572082
rect 186320 572018 186372 572024
rect 43444 572008 43496 572014
rect 43444 571950 43496 571956
rect 168380 572008 168432 572014
rect 284312 571985 284340 587302
rect 292580 586492 292632 586498
rect 292580 586434 292632 586440
rect 292592 586401 292620 586434
rect 292578 586392 292634 586401
rect 292578 586327 292634 586336
rect 290004 586084 290056 586090
rect 290004 586026 290056 586032
rect 289912 586016 289964 586022
rect 289912 585958 289964 585964
rect 289820 585948 289872 585954
rect 289820 585890 289872 585896
rect 288440 585880 288492 585886
rect 288440 585822 288492 585828
rect 168380 571950 168432 571956
rect 284298 571976 284354 571985
rect 284298 571911 284354 571920
rect 23388 463412 23440 463418
rect 23388 463354 23440 463360
rect 21928 460906 22048 460934
rect 20628 459536 20680 459542
rect 20628 459478 20680 459484
rect 20536 458720 20588 458726
rect 20536 458662 20588 458668
rect 20444 457972 20496 457978
rect 20444 457914 20496 457920
rect 20456 332382 20484 457914
rect 20548 332450 20576 458662
rect 21928 457910 21956 460906
rect 23400 458833 23428 463354
rect 140148 462466 140484 462482
rect 24860 462460 24912 462466
rect 24860 462402 24912 462408
rect 140136 462460 140484 462466
rect 140188 462454 140484 462460
rect 140136 462402 140188 462408
rect 24216 462256 24268 462262
rect 24268 462204 24564 462210
rect 24216 462198 24564 462204
rect 24228 462182 24564 462198
rect 24872 461650 24900 462402
rect 151912 462392 151964 462398
rect 151964 462340 152076 462346
rect 151912 462334 152076 462340
rect 151924 462318 152076 462334
rect 288256 462324 288308 462330
rect 288256 462266 288308 462272
rect 24860 461644 24912 461650
rect 24860 461586 24912 461592
rect 288268 461310 288296 462266
rect 158168 461304 158220 461310
rect 30024 461230 30360 461258
rect 35912 461230 36156 461258
rect 41616 461230 41952 461258
rect 47412 461230 47748 461258
rect 53208 461230 53544 461258
rect 59004 461230 59340 461258
rect 64892 461230 65136 461258
rect 70596 461230 70932 461258
rect 76392 461230 76728 461258
rect 82188 461230 82524 461258
rect 87984 461230 88320 461258
rect 93872 461230 94116 461258
rect 99576 461230 99912 461258
rect 105372 461230 105708 461258
rect 111168 461230 111504 461258
rect 116964 461230 117300 461258
rect 122852 461230 123096 461258
rect 128892 461230 129228 461258
rect 26240 461032 26292 461038
rect 26240 460974 26292 460980
rect 23386 458824 23442 458833
rect 23386 458759 23442 458768
rect 23400 458266 23428 458759
rect 23400 458238 23520 458266
rect 21916 457904 21968 457910
rect 21916 457846 21968 457852
rect 21824 333328 21876 333334
rect 21824 333270 21876 333276
rect 20536 332444 20588 332450
rect 20536 332386 20588 332392
rect 20444 332376 20496 332382
rect 20444 332318 20496 332324
rect 20352 332240 20404 332246
rect 20352 332182 20404 332188
rect 20364 204241 20392 332182
rect 20456 331430 20484 332318
rect 20444 331424 20496 331430
rect 20444 331366 20496 331372
rect 20548 331362 20576 332386
rect 20536 331356 20588 331362
rect 20536 331298 20588 331304
rect 20444 331288 20496 331294
rect 20444 331230 20496 331236
rect 20350 204232 20406 204241
rect 20350 204167 20406 204176
rect 20258 204096 20314 204105
rect 20258 204031 20314 204040
rect 20180 203918 20392 203946
rect 20258 202872 20314 202881
rect 20076 202836 20128 202842
rect 20258 202807 20314 202816
rect 20076 202778 20128 202784
rect 20272 76022 20300 202807
rect 20364 202774 20392 203918
rect 20352 202768 20404 202774
rect 20352 202710 20404 202716
rect 20260 76016 20312 76022
rect 20260 75958 20312 75964
rect 19248 75676 19300 75682
rect 19248 75618 19300 75624
rect 20364 75614 20392 202710
rect 20456 202706 20484 331230
rect 20534 204232 20590 204241
rect 20534 204167 20590 204176
rect 20548 203697 20576 204167
rect 20626 204096 20682 204105
rect 20626 204031 20682 204040
rect 20534 203688 20590 203697
rect 20534 203623 20590 203632
rect 20444 202700 20496 202706
rect 20444 202642 20496 202648
rect 20352 75608 20404 75614
rect 20352 75550 20404 75556
rect 19156 74520 19208 74526
rect 19156 74462 19208 74468
rect 20456 74322 20484 202642
rect 20444 74316 20496 74322
rect 20444 74258 20496 74264
rect 20548 74186 20576 203623
rect 20640 74254 20668 204031
rect 21836 203930 21864 333270
rect 21928 332518 21956 457846
rect 23492 443426 23520 458238
rect 26252 458182 26280 460974
rect 30024 459542 30052 461230
rect 30012 459536 30064 459542
rect 30012 459478 30064 459484
rect 35912 459066 35940 461230
rect 41616 459542 41644 461230
rect 41604 459536 41656 459542
rect 41604 459478 41656 459484
rect 30932 459060 30984 459066
rect 30932 459002 30984 459008
rect 35900 459060 35952 459066
rect 35900 459002 35952 459008
rect 30944 458969 30972 459002
rect 30930 458960 30986 458969
rect 30930 458895 30986 458904
rect 26240 458176 26292 458182
rect 26240 458118 26292 458124
rect 47412 457910 47440 461230
rect 53208 457978 53236 461230
rect 53196 457972 53248 457978
rect 53196 457914 53248 457920
rect 47400 457904 47452 457910
rect 47400 457846 47452 457852
rect 59004 456890 59032 461230
rect 64892 458862 64920 461230
rect 64880 458856 64932 458862
rect 64880 458798 64932 458804
rect 70596 458153 70624 461230
rect 70582 458144 70638 458153
rect 70582 458079 70638 458088
rect 76392 458046 76420 461230
rect 82188 459513 82216 461230
rect 82174 459504 82230 459513
rect 82174 459439 82230 459448
rect 87984 459338 88012 461230
rect 87972 459332 88024 459338
rect 87972 459274 88024 459280
rect 93872 458114 93900 461230
rect 99576 459406 99604 461230
rect 99564 459400 99616 459406
rect 99564 459342 99616 459348
rect 105372 459202 105400 461230
rect 105360 459196 105412 459202
rect 105360 459138 105412 459144
rect 111168 458182 111196 461230
rect 116964 459270 116992 461230
rect 116952 459264 117004 459270
rect 116952 459206 117004 459212
rect 122852 458833 122880 461230
rect 129200 459542 129228 461230
rect 134352 461230 134688 461258
rect 145944 461230 146280 461258
rect 157872 461252 158168 461258
rect 288256 461304 288308 461310
rect 157872 461246 158220 461252
rect 157872 461230 158208 461246
rect 134352 459542 134380 461230
rect 145944 460970 145972 461230
rect 163654 461038 163682 461244
rect 169464 461230 169708 461258
rect 163642 461032 163694 461038
rect 163642 460974 163694 460980
rect 145932 460964 145984 460970
rect 145932 460906 145984 460912
rect 129188 459536 129240 459542
rect 129188 459478 129240 459484
rect 134340 459536 134392 459542
rect 134340 459478 134392 459484
rect 134352 458833 134380 459478
rect 122838 458824 122894 458833
rect 122838 458759 122894 458768
rect 134338 458824 134394 458833
rect 134338 458759 134394 458768
rect 169680 458182 169708 461230
rect 175246 461106 175274 461244
rect 181056 461230 181392 461258
rect 186852 461230 187188 461258
rect 192648 461230 192984 461258
rect 198444 461230 198688 461258
rect 181364 461174 181392 461230
rect 181352 461168 181404 461174
rect 181352 461110 181404 461116
rect 175234 461100 175286 461106
rect 175234 461042 175286 461048
rect 187160 459542 187188 461230
rect 192956 460902 192984 461230
rect 192944 460896 192996 460902
rect 192944 460838 192996 460844
rect 187148 459536 187200 459542
rect 187148 459478 187200 459484
rect 198660 458969 198688 461230
rect 204180 461230 204240 461258
rect 210036 461230 210372 461258
rect 215832 461230 216168 461258
rect 221628 461230 221964 461258
rect 204180 459474 204208 461230
rect 204168 459468 204220 459474
rect 204168 459410 204220 459416
rect 210344 459270 210372 461230
rect 216140 459406 216168 461230
rect 216128 459400 216180 459406
rect 216128 459342 216180 459348
rect 221936 459338 221964 461230
rect 227410 461009 227438 461244
rect 233220 461242 233372 461258
rect 233220 461236 233384 461242
rect 233220 461230 233332 461236
rect 239016 461230 239352 461258
rect 244812 461230 245148 461258
rect 250608 461230 250944 461258
rect 256404 461230 256648 461258
rect 233332 461178 233384 461184
rect 227396 461000 227452 461009
rect 227396 460935 227452 460944
rect 221924 459332 221976 459338
rect 221924 459274 221976 459280
rect 210332 459264 210384 459270
rect 210332 459206 210384 459212
rect 198646 458960 198702 458969
rect 198646 458895 198702 458904
rect 111156 458176 111208 458182
rect 111156 458118 111208 458124
rect 169668 458176 169720 458182
rect 239324 458153 239352 461230
rect 169668 458118 169720 458124
rect 239310 458144 239366 458153
rect 93860 458108 93912 458114
rect 245120 458114 245148 461230
rect 239310 458079 239366 458088
rect 245108 458108 245160 458114
rect 93860 458050 93912 458056
rect 245108 458050 245160 458056
rect 250916 458046 250944 461230
rect 76380 458040 76432 458046
rect 76380 457982 76432 457988
rect 250904 458040 250956 458046
rect 250904 457982 250956 457988
rect 256620 457978 256648 461230
rect 262140 461230 262200 461258
rect 267996 461230 268332 461258
rect 273792 461230 274128 461258
rect 279588 461230 279924 461258
rect 256608 457972 256660 457978
rect 256608 457914 256660 457920
rect 262140 457910 262168 461230
rect 268304 458862 268332 461230
rect 274100 458930 274128 461230
rect 279896 459202 279924 461230
rect 284312 461230 285384 461258
rect 288256 461246 288308 461252
rect 280712 460964 280764 460970
rect 280712 460906 280764 460912
rect 280724 459270 280752 460906
rect 280712 459264 280764 459270
rect 280712 459206 280764 459212
rect 279884 459196 279936 459202
rect 279884 459138 279936 459144
rect 274088 458924 274140 458930
rect 274088 458866 274140 458872
rect 268292 458856 268344 458862
rect 268292 458798 268344 458804
rect 280068 458856 280120 458862
rect 280068 458798 280120 458804
rect 262128 457904 262180 457910
rect 262128 457846 262180 457852
rect 280080 457502 280108 458798
rect 280068 457496 280120 457502
rect 280068 457438 280120 457444
rect 55956 456884 56008 456890
rect 55956 456826 56008 456832
rect 58992 456884 59044 456890
rect 58992 456826 59044 456832
rect 55968 456074 55996 456826
rect 55956 456068 56008 456074
rect 55956 456010 56008 456016
rect 284312 443698 284340 461230
rect 287612 457972 287664 457978
rect 287612 457914 287664 457920
rect 287624 457881 287652 457914
rect 287610 457872 287666 457881
rect 287610 457807 287666 457816
rect 288268 456346 288296 461246
rect 288452 457978 288480 585822
rect 288624 585812 288676 585818
rect 288624 585754 288676 585760
rect 288532 580372 288584 580378
rect 288532 580314 288584 580320
rect 288544 462330 288572 580314
rect 288532 462324 288584 462330
rect 288532 462266 288584 462272
rect 288530 461000 288586 461009
rect 288530 460935 288586 460944
rect 288440 457972 288492 457978
rect 288440 457914 288492 457920
rect 288256 456340 288308 456346
rect 288256 456282 288308 456288
rect 284300 443692 284352 443698
rect 284300 443634 284352 443640
rect 23480 443420 23532 443426
rect 23480 443362 23532 443368
rect 27528 334008 27580 334014
rect 27528 333950 27580 333956
rect 24228 333254 24564 333282
rect 26240 333260 26292 333266
rect 22006 332888 22062 332897
rect 22006 332823 22008 332832
rect 22060 332823 22062 332832
rect 22008 332794 22060 332800
rect 24228 332722 24256 333254
rect 26240 333202 26292 333208
rect 24216 332716 24268 332722
rect 24216 332658 24268 332664
rect 21916 332512 21968 332518
rect 21916 332454 21968 332460
rect 21928 331294 21956 332454
rect 23386 332208 23442 332217
rect 23386 332143 23388 332152
rect 23440 332143 23442 332152
rect 23388 332114 23440 332120
rect 21916 331288 21968 331294
rect 21916 331230 21968 331236
rect 24860 330540 24912 330546
rect 24860 330482 24912 330488
rect 24872 329662 24900 330482
rect 24860 329656 24912 329662
rect 24860 329598 24912 329604
rect 26252 325694 26280 333202
rect 27540 332722 27568 333950
rect 286968 333328 287020 333334
rect 280802 333296 280858 333305
rect 30024 333254 30360 333282
rect 36004 333254 36156 333282
rect 41616 333254 41952 333282
rect 47412 333254 47748 333282
rect 53208 333254 53544 333282
rect 59004 333254 59340 333282
rect 64984 333254 65136 333282
rect 70596 333254 70932 333282
rect 76392 333254 76728 333282
rect 82188 333254 82524 333282
rect 87984 333254 88320 333282
rect 93872 333254 94116 333282
rect 99576 333254 99912 333282
rect 105372 333254 105708 333282
rect 111168 333254 111504 333282
rect 116964 333254 117300 333282
rect 122760 333254 123096 333282
rect 128892 333254 129228 333282
rect 134688 333254 135024 333282
rect 27528 332716 27580 332722
rect 27528 332658 27580 332664
rect 30024 332586 30052 333254
rect 30012 332580 30064 332586
rect 30012 332522 30064 332528
rect 31024 332580 31076 332586
rect 31024 332522 31076 332528
rect 31036 332382 31064 332522
rect 31024 332376 31076 332382
rect 31024 332318 31076 332324
rect 36004 332246 36032 333254
rect 41616 332314 41644 333254
rect 47412 332382 47440 333254
rect 53208 332450 53236 333254
rect 56508 332988 56560 332994
rect 56508 332930 56560 332936
rect 56520 332586 56548 332930
rect 59004 332586 59032 333254
rect 56508 332580 56560 332586
rect 56508 332522 56560 332528
rect 58992 332580 59044 332586
rect 58992 332522 59044 332528
rect 64984 332518 65012 333254
rect 64972 332512 65024 332518
rect 64972 332454 65024 332460
rect 53196 332444 53248 332450
rect 53196 332386 53248 332392
rect 47400 332376 47452 332382
rect 47400 332318 47452 332324
rect 41604 332308 41656 332314
rect 41604 332250 41656 332256
rect 35992 332240 36044 332246
rect 35992 332182 36044 332188
rect 70596 332178 70624 333254
rect 76392 332489 76420 333254
rect 82188 332858 82216 333254
rect 82176 332852 82228 332858
rect 82176 332794 82228 332800
rect 76378 332480 76434 332489
rect 76378 332415 76434 332424
rect 70584 332172 70636 332178
rect 70584 332114 70636 332120
rect 87984 329730 88012 333254
rect 87972 329724 88024 329730
rect 87972 329666 88024 329672
rect 26252 325666 26372 325694
rect 26344 315994 26372 325666
rect 26332 315988 26384 315994
rect 26332 315930 26384 315936
rect 26344 315450 26372 315930
rect 93872 315926 93900 333254
rect 99576 332790 99604 333254
rect 99564 332784 99616 332790
rect 99564 332726 99616 332732
rect 105372 332654 105400 333254
rect 111168 332722 111196 333254
rect 111156 332716 111208 332722
rect 111156 332658 111208 332664
rect 105360 332648 105412 332654
rect 105360 332590 105412 332596
rect 116964 329798 116992 333254
rect 122760 332926 122788 333254
rect 122748 332920 122800 332926
rect 122748 332862 122800 332868
rect 129200 332586 129228 333254
rect 134996 332586 135024 333254
rect 139412 333254 140484 333282
rect 145944 333254 146280 333282
rect 151832 333254 152076 333282
rect 157352 333254 157872 333282
rect 162872 333254 163668 333282
rect 169464 333254 169800 333282
rect 129188 332580 129240 332586
rect 129188 332522 129240 332528
rect 134984 332580 135036 332586
rect 134984 332522 135036 332528
rect 134996 331906 135024 332522
rect 134984 331900 135036 331906
rect 134984 331842 135036 331848
rect 116952 329792 117004 329798
rect 116952 329734 117004 329740
rect 139412 315994 139440 333254
rect 145944 330546 145972 333254
rect 145932 330540 145984 330546
rect 145932 330482 145984 330488
rect 139400 315988 139452 315994
rect 139400 315930 139452 315936
rect 93860 315920 93912 315926
rect 93860 315862 93912 315868
rect 26332 315444 26384 315450
rect 26332 315386 26384 315392
rect 151832 315382 151860 333254
rect 157352 315994 157380 333254
rect 157340 315988 157392 315994
rect 157340 315930 157392 315936
rect 27528 315376 27580 315382
rect 27528 315318 27580 315324
rect 151820 315376 151872 315382
rect 151820 315318 151872 315324
rect 27540 314634 27568 315318
rect 157352 315314 157380 315930
rect 157340 315308 157392 315314
rect 157340 315250 157392 315256
rect 162872 314634 162900 333254
rect 169772 332858 169800 333254
rect 175200 333254 175260 333282
rect 181056 333254 181392 333282
rect 169760 332852 169812 332858
rect 169760 332794 169812 332800
rect 175200 331809 175228 333254
rect 181364 332654 181392 333254
rect 186332 333254 186852 333282
rect 192648 333254 192984 333282
rect 198444 333254 198688 333282
rect 181352 332648 181404 332654
rect 181352 332590 181404 332596
rect 175186 331800 175242 331809
rect 175186 331735 175242 331744
rect 186332 331242 186360 333254
rect 186240 331214 186360 331242
rect 192956 331226 192984 333254
rect 198660 331974 198688 333254
rect 204180 333254 204240 333282
rect 210036 333254 210372 333282
rect 215832 333254 216168 333282
rect 221628 333254 221964 333282
rect 198648 331968 198700 331974
rect 198648 331910 198700 331916
rect 192944 331220 192996 331226
rect 186240 315926 186268 331214
rect 192944 331162 192996 331168
rect 204180 330546 204208 333254
rect 210344 332722 210372 333254
rect 216140 332790 216168 333254
rect 216128 332784 216180 332790
rect 216128 332726 216180 332732
rect 210332 332716 210384 332722
rect 210332 332658 210384 332664
rect 221936 331158 221964 333254
rect 226352 333254 227424 333282
rect 231872 333254 233220 333282
rect 239016 333254 239352 333282
rect 244812 333254 245148 333282
rect 250608 333254 250944 333282
rect 256404 333254 256648 333282
rect 221924 331152 221976 331158
rect 221924 331094 221976 331100
rect 204168 330540 204220 330546
rect 204168 330482 204220 330488
rect 186228 315920 186280 315926
rect 186228 315862 186280 315868
rect 226352 315858 226380 333254
rect 226340 315852 226392 315858
rect 226340 315794 226392 315800
rect 231872 315790 231900 333254
rect 239324 332926 239352 333254
rect 239312 332920 239364 332926
rect 239312 332862 239364 332868
rect 245120 331294 245148 333254
rect 250916 332994 250944 333254
rect 250904 332988 250956 332994
rect 250904 332930 250956 332936
rect 256620 332586 256648 333254
rect 262140 333254 262200 333282
rect 267996 333254 268332 333282
rect 256608 332580 256660 332586
rect 256608 332522 256660 332528
rect 262140 332518 262168 333254
rect 262128 332512 262180 332518
rect 262128 332454 262180 332460
rect 268304 332450 268332 333254
rect 273272 333254 273792 333282
rect 279588 333254 279924 333282
rect 268292 332444 268344 332450
rect 268292 332386 268344 332392
rect 245108 331288 245160 331294
rect 245108 331230 245160 331236
rect 246304 331288 246356 331294
rect 246304 331230 246356 331236
rect 231860 315784 231912 315790
rect 231860 315726 231912 315732
rect 246316 315722 246344 331230
rect 246304 315716 246356 315722
rect 246304 315658 246356 315664
rect 273272 315314 273300 333254
rect 279896 332382 279924 333254
rect 280802 333231 280858 333240
rect 281448 333260 281500 333266
rect 279884 332376 279936 332382
rect 279884 332318 279936 332324
rect 280816 315994 280844 333231
rect 285384 333254 285628 333282
rect 286968 333270 287020 333276
rect 281448 333202 281500 333208
rect 281460 316062 281488 333202
rect 282184 332920 282236 332926
rect 282184 332862 282236 332868
rect 282196 331770 282224 332862
rect 285600 332042 285628 333254
rect 285588 332036 285640 332042
rect 285588 331978 285640 331984
rect 282184 331764 282236 331770
rect 282184 331706 282236 331712
rect 285588 331764 285640 331770
rect 285588 331706 285640 331712
rect 285600 331401 285628 331706
rect 285586 331392 285642 331401
rect 285586 331327 285642 331336
rect 281448 316056 281500 316062
rect 281448 315998 281500 316004
rect 280804 315988 280856 315994
rect 280804 315930 280856 315936
rect 285600 315382 285628 331327
rect 285588 315376 285640 315382
rect 285588 315318 285640 315324
rect 273260 315308 273312 315314
rect 273260 315250 273312 315256
rect 27528 314628 27580 314634
rect 27528 314570 27580 314576
rect 162860 314628 162912 314634
rect 162860 314570 162912 314576
rect 285772 314628 285824 314634
rect 285772 314570 285824 314576
rect 285784 313954 285812 314570
rect 286980 313954 287008 333270
rect 287796 332580 287848 332586
rect 287796 332522 287848 332528
rect 287808 332489 287836 332522
rect 287794 332480 287850 332489
rect 287794 332415 287850 332424
rect 288440 331900 288492 331906
rect 288440 331842 288492 331848
rect 285772 313948 285824 313954
rect 285772 313890 285824 313896
rect 286968 313948 287020 313954
rect 286968 313890 287020 313896
rect 145930 206408 145986 206417
rect 145986 206366 146280 206394
rect 145930 206343 145986 206352
rect 24952 206304 25004 206310
rect 24952 206246 25004 206252
rect 151910 206272 151966 206281
rect 24228 205278 24564 205306
rect 24124 204196 24176 204202
rect 24124 204138 24176 204144
rect 21824 203924 21876 203930
rect 21824 203866 21876 203872
rect 21836 203833 21864 203866
rect 21822 203824 21878 203833
rect 21822 203759 21878 203768
rect 23386 202872 23442 202881
rect 22008 202836 22060 202842
rect 23386 202807 23388 202816
rect 22008 202778 22060 202784
rect 23440 202807 23442 202816
rect 23388 202778 23440 202784
rect 22020 202230 22048 202778
rect 22008 202224 22060 202230
rect 22008 202166 22060 202172
rect 22020 74390 22048 202166
rect 22100 199436 22152 199442
rect 22100 199378 22152 199384
rect 22112 186386 22140 199378
rect 24136 186454 24164 204138
rect 24228 204134 24256 205278
rect 24860 204944 24912 204950
rect 24860 204886 24912 204892
rect 24216 204128 24268 204134
rect 24216 204070 24268 204076
rect 24872 203862 24900 204886
rect 24964 204134 24992 206246
rect 151966 206230 152076 206258
rect 151910 206207 151966 206216
rect 30024 205278 30360 205306
rect 36004 205278 36156 205306
rect 41616 205278 41952 205306
rect 47412 205278 47748 205306
rect 53208 205278 53544 205306
rect 59004 205278 59340 205306
rect 64984 205278 65136 205306
rect 70596 205278 70932 205306
rect 76392 205278 76728 205306
rect 82188 205278 82524 205306
rect 87984 205278 88320 205306
rect 93964 205278 94116 205306
rect 99576 205278 99912 205306
rect 105372 205278 105708 205306
rect 111168 205278 111504 205306
rect 116964 205278 117300 205306
rect 122852 205278 123096 205306
rect 128892 205278 129228 205306
rect 134688 205278 135024 205306
rect 30024 204270 30052 205278
rect 36004 204270 36032 205278
rect 30012 204264 30064 204270
rect 30012 204206 30064 204212
rect 33140 204264 33192 204270
rect 33140 204206 33192 204212
rect 35992 204264 36044 204270
rect 41616 204241 41644 205278
rect 35992 204206 36044 204212
rect 41602 204232 41658 204241
rect 25044 204196 25096 204202
rect 25044 204138 25096 204144
rect 24952 204128 25004 204134
rect 24952 204070 25004 204076
rect 24860 203856 24912 203862
rect 24860 203798 24912 203804
rect 25056 203794 25084 204138
rect 25504 203856 25556 203862
rect 25504 203798 25556 203804
rect 25044 203788 25096 203794
rect 25044 203730 25096 203736
rect 25516 187134 25544 203798
rect 33152 203697 33180 204206
rect 41602 204167 41658 204176
rect 33138 203688 33194 203697
rect 33138 203623 33194 203632
rect 47412 202706 47440 205278
rect 47400 202700 47452 202706
rect 47400 202642 47452 202648
rect 53208 202230 53236 205278
rect 59004 203930 59032 205278
rect 58992 203924 59044 203930
rect 58992 203866 59044 203872
rect 64984 202774 65012 205278
rect 70596 202842 70624 205278
rect 70584 202836 70636 202842
rect 70584 202778 70636 202784
rect 64972 202768 65024 202774
rect 64972 202710 65024 202716
rect 53196 202224 53248 202230
rect 53196 202166 53248 202172
rect 76392 202162 76420 205278
rect 82188 202881 82216 205278
rect 87984 204338 88012 205278
rect 87972 204332 88024 204338
rect 87972 204274 88024 204280
rect 93964 203998 93992 205278
rect 99576 204066 99604 205278
rect 105372 204202 105400 205278
rect 105360 204196 105412 204202
rect 105360 204138 105412 204144
rect 111168 204134 111196 205278
rect 111156 204128 111208 204134
rect 111156 204070 111208 204076
rect 99564 204060 99616 204066
rect 99564 204002 99616 204008
rect 93952 203992 94004 203998
rect 93952 203934 94004 203940
rect 116964 203561 116992 205278
rect 116950 203552 117006 203561
rect 116950 203487 117006 203496
rect 82174 202872 82230 202881
rect 122852 202874 122880 205278
rect 129200 204270 129228 205278
rect 134996 204270 135024 205278
rect 140148 205278 140484 205306
rect 157536 205278 157872 205306
rect 162872 205278 163668 205306
rect 168392 205278 169464 205306
rect 175200 205278 175260 205306
rect 181056 205278 181484 205306
rect 129188 204264 129240 204270
rect 129188 204206 129240 204212
rect 134984 204264 135036 204270
rect 134984 204206 135036 204212
rect 134996 203590 135024 204206
rect 140148 203862 140176 205278
rect 140136 203856 140188 203862
rect 140136 203798 140188 203804
rect 134984 203584 135036 203590
rect 134984 203526 135036 203532
rect 82174 202807 82230 202816
rect 122760 202846 122880 202874
rect 76380 202156 76432 202162
rect 76380 202098 76432 202104
rect 122760 199442 122788 202846
rect 157536 200705 157564 205278
rect 157522 200696 157578 200705
rect 157522 200631 157578 200640
rect 122748 199436 122800 199442
rect 122748 199378 122800 199384
rect 162872 189038 162900 205278
rect 162860 189032 162912 189038
rect 162860 188974 162912 188980
rect 162872 188426 162900 188974
rect 168392 188970 168420 205278
rect 175200 204338 175228 205278
rect 175188 204332 175240 204338
rect 175188 204274 175240 204280
rect 181456 201482 181484 205278
rect 186332 205278 186852 205306
rect 192648 205278 192984 205306
rect 198444 205278 198688 205306
rect 181444 201476 181496 201482
rect 181444 201418 181496 201424
rect 168380 188964 168432 188970
rect 168380 188906 168432 188912
rect 103980 188420 104032 188426
rect 103980 188362 104032 188368
rect 162860 188420 162912 188426
rect 162860 188362 162912 188368
rect 25504 187128 25556 187134
rect 25504 187070 25556 187076
rect 103992 187066 104020 188362
rect 181456 188358 181484 201418
rect 186332 188902 186360 205278
rect 192956 204406 192984 205278
rect 192944 204400 192996 204406
rect 192944 204342 192996 204348
rect 198660 203561 198688 205278
rect 204180 205278 204240 205306
rect 210036 205278 210372 205306
rect 215832 205278 216168 205306
rect 221628 205278 221964 205306
rect 227424 205278 227668 205306
rect 204180 204474 204208 205278
rect 204168 204468 204220 204474
rect 204168 204410 204220 204416
rect 210344 203697 210372 205278
rect 216140 203998 216168 205278
rect 221936 204542 221964 205278
rect 221924 204536 221976 204542
rect 221924 204478 221976 204484
rect 227640 204202 227668 205278
rect 233160 205278 233220 205306
rect 239016 205278 239352 205306
rect 244812 205278 245148 205306
rect 250608 205278 250944 205306
rect 256404 205278 256648 205306
rect 227628 204196 227680 204202
rect 227628 204138 227680 204144
rect 216128 203992 216180 203998
rect 216128 203934 216180 203940
rect 210330 203688 210386 203697
rect 233160 203658 233188 205278
rect 239324 204134 239352 205278
rect 245120 204610 245148 205278
rect 245108 204604 245160 204610
rect 245108 204546 245160 204552
rect 239312 204128 239364 204134
rect 239312 204070 239364 204076
rect 210330 203623 210386 203632
rect 233148 203652 233200 203658
rect 233148 203594 233200 203600
rect 198646 203552 198702 203561
rect 198646 203487 198702 203496
rect 250916 202842 250944 205278
rect 250904 202836 250956 202842
rect 250904 202778 250956 202784
rect 256620 202774 256648 205278
rect 262140 205278 262200 205306
rect 267996 205278 268332 205306
rect 273792 205278 274128 205306
rect 279588 205278 279924 205306
rect 285384 205278 285628 205306
rect 256608 202768 256660 202774
rect 256608 202710 256660 202716
rect 262140 202162 262168 205278
rect 268304 204066 268332 205278
rect 268292 204060 268344 204066
rect 268292 204002 268344 204008
rect 274100 203726 274128 205278
rect 276662 204912 276718 204921
rect 276662 204847 276718 204856
rect 274088 203720 274140 203726
rect 274088 203662 274140 203668
rect 262128 202156 262180 202162
rect 262128 202098 262180 202104
rect 276676 188970 276704 204847
rect 279896 204270 279924 205278
rect 283288 205012 283340 205018
rect 283288 204954 283340 204960
rect 283300 204270 283328 204954
rect 279884 204264 279936 204270
rect 279884 204206 279936 204212
rect 283288 204264 283340 204270
rect 283288 204206 283340 204212
rect 280068 204060 280120 204066
rect 280068 204002 280120 204008
rect 280080 203833 280108 204002
rect 280066 203824 280122 203833
rect 285600 203794 285628 205278
rect 288256 204468 288308 204474
rect 288256 204410 288308 204416
rect 287336 204332 287388 204338
rect 287336 204274 287388 204280
rect 280066 203759 280122 203768
rect 285588 203788 285640 203794
rect 285588 203730 285640 203736
rect 287348 202881 287376 204274
rect 287334 202872 287390 202881
rect 287334 202807 287390 202816
rect 287886 202872 287942 202881
rect 287886 202807 287942 202816
rect 287900 202774 287928 202807
rect 287888 202768 287940 202774
rect 287888 202710 287940 202716
rect 276664 188964 276716 188970
rect 276664 188906 276716 188912
rect 186320 188896 186372 188902
rect 186320 188838 186372 188844
rect 181444 188352 181496 188358
rect 181444 188294 181496 188300
rect 103980 187060 104032 187066
rect 103980 187002 104032 187008
rect 186332 186998 186360 188838
rect 186320 186992 186372 186998
rect 186320 186934 186372 186940
rect 24124 186448 24176 186454
rect 24124 186390 24176 186396
rect 22100 186380 22152 186386
rect 22100 186322 22152 186328
rect 276676 185910 276704 188906
rect 288268 186930 288296 204410
rect 288348 204400 288400 204406
rect 288348 204342 288400 204348
rect 288256 186924 288308 186930
rect 288256 186866 288308 186872
rect 288360 186386 288388 204342
rect 288348 186380 288400 186386
rect 288348 186322 288400 186328
rect 276664 185904 276716 185910
rect 276664 185846 276716 185852
rect 287702 79384 287758 79393
rect 287702 79319 287758 79328
rect 82820 78192 82872 78198
rect 82820 78134 82872 78140
rect 24228 77302 24564 77330
rect 30024 77302 30360 77330
rect 36096 77302 36156 77330
rect 41892 77302 41952 77330
rect 24228 75478 24256 77302
rect 30024 75886 30052 77302
rect 30012 75880 30064 75886
rect 30012 75822 30064 75828
rect 24216 75472 24268 75478
rect 24216 75414 24268 75420
rect 22008 74384 22060 74390
rect 22008 74326 22060 74332
rect 20628 74248 20680 74254
rect 20628 74190 20680 74196
rect 36096 74186 36124 77302
rect 41892 74254 41920 77302
rect 47734 77058 47762 77316
rect 53530 77058 53558 77316
rect 59280 77302 59340 77330
rect 65076 77302 65136 77330
rect 70932 77302 71084 77330
rect 47734 77030 47808 77058
rect 53530 77030 53604 77058
rect 47780 74322 47808 77030
rect 53576 74390 53604 77030
rect 59280 75857 59308 77302
rect 59266 75848 59322 75857
rect 59266 75783 59322 75792
rect 59280 75206 59308 75783
rect 65076 75614 65104 77302
rect 65064 75608 65116 75614
rect 65064 75550 65116 75556
rect 65524 75608 65576 75614
rect 65524 75550 65576 75556
rect 59268 75200 59320 75206
rect 59268 75142 59320 75148
rect 53564 74384 53616 74390
rect 53564 74326 53616 74332
rect 47768 74316 47820 74322
rect 47768 74258 47820 74264
rect 41880 74248 41932 74254
rect 41880 74190 41932 74196
rect 20536 74180 20588 74186
rect 20536 74122 20588 74128
rect 36084 74180 36136 74186
rect 36084 74122 36136 74128
rect 41892 72486 41920 74190
rect 41880 72480 41932 72486
rect 41880 72422 41932 72428
rect 47780 69698 47808 74258
rect 47768 69692 47820 69698
rect 47768 69634 47820 69640
rect 53576 68338 53604 74326
rect 53564 68332 53616 68338
rect 53564 68274 53616 68280
rect 57612 64184 57664 64190
rect 57612 64126 57664 64132
rect 57624 61713 57652 64126
rect 65536 62830 65564 75550
rect 71056 74361 71084 77302
rect 76714 77110 76742 77316
rect 82188 77302 82524 77330
rect 75920 77104 75972 77110
rect 75920 77046 75972 77052
rect 76702 77104 76754 77110
rect 76702 77046 76754 77052
rect 75932 76090 75960 77046
rect 75920 76084 75972 76090
rect 75920 76026 75972 76032
rect 71042 74352 71098 74361
rect 71042 74287 71098 74296
rect 71056 62898 71084 74287
rect 75932 62966 75960 76026
rect 82188 76022 82216 77302
rect 82176 76016 82228 76022
rect 82176 75958 82228 75964
rect 82544 76016 82596 76022
rect 82544 75958 82596 75964
rect 82556 68406 82584 75958
rect 82832 75886 82860 78134
rect 111168 78130 111748 78146
rect 279588 78130 279924 78146
rect 111156 78124 111748 78130
rect 111208 78118 111748 78124
rect 111156 78066 111208 78072
rect 88260 77302 88320 77330
rect 94056 77302 94116 77330
rect 99912 77302 100248 77330
rect 82820 75880 82872 75886
rect 82820 75822 82872 75828
rect 88260 75546 88288 77302
rect 94056 75682 94084 77302
rect 100220 75750 100248 77302
rect 105694 77058 105722 77316
rect 105694 77030 105768 77058
rect 105740 75818 105768 77030
rect 105728 75812 105780 75818
rect 105728 75754 105780 75760
rect 100208 75744 100260 75750
rect 100208 75686 100260 75692
rect 94044 75676 94096 75682
rect 94044 75618 94096 75624
rect 88248 75540 88300 75546
rect 88248 75482 88300 75488
rect 88260 71058 88288 75482
rect 94056 72554 94084 75618
rect 94044 72548 94096 72554
rect 94044 72490 94096 72496
rect 88248 71052 88300 71058
rect 88248 70994 88300 71000
rect 100220 69766 100248 75686
rect 100208 69760 100260 69766
rect 100208 69702 100260 69708
rect 105740 68474 105768 75754
rect 111720 71126 111748 78118
rect 278780 78124 278832 78130
rect 279588 78124 279936 78130
rect 279588 78118 279884 78124
rect 278780 78066 278832 78072
rect 279884 78066 279936 78072
rect 144920 78056 144972 78062
rect 264980 78056 265032 78062
rect 247038 78024 247094 78033
rect 144920 77998 144972 78004
rect 116964 77302 117300 77330
rect 123036 77302 123096 77330
rect 128892 77302 129228 77330
rect 116964 74458 116992 77302
rect 123036 74526 123064 77302
rect 129200 75818 129228 77302
rect 134536 77302 134688 77330
rect 140056 77302 140484 77330
rect 144932 77314 144960 77998
rect 151924 77994 152076 78010
rect 151912 77988 152076 77994
rect 151964 77982 152076 77988
rect 264980 77998 265032 78004
rect 247038 77959 247094 77968
rect 151912 77930 151964 77936
rect 151924 77330 151952 77930
rect 235262 77888 235318 77897
rect 235262 77823 235318 77832
rect 145944 77314 146280 77330
rect 144920 77308 144972 77314
rect 134536 75818 134564 77302
rect 129188 75812 129240 75818
rect 129188 75754 129240 75760
rect 134524 75812 134576 75818
rect 134524 75754 134576 75760
rect 123484 75200 123536 75206
rect 123484 75142 123536 75148
rect 123024 74520 123076 74526
rect 123024 74462 123076 74468
rect 116952 74452 117004 74458
rect 116952 74394 117004 74400
rect 111708 71120 111760 71126
rect 111708 71062 111760 71068
rect 105728 68468 105780 68474
rect 105728 68410 105780 68416
rect 82544 68400 82596 68406
rect 82544 68342 82596 68348
rect 116964 66978 116992 74394
rect 116952 66972 117004 66978
rect 116952 66914 117004 66920
rect 123496 63034 123524 75142
rect 124128 74520 124180 74526
rect 124128 74462 124180 74468
rect 124140 73914 124168 74462
rect 124128 73908 124180 73914
rect 124128 73850 124180 73856
rect 134536 67046 134564 75754
rect 140056 73166 140084 77302
rect 144920 77250 144972 77256
rect 145932 77308 146280 77314
rect 145984 77302 146280 77308
rect 151832 77302 151952 77330
rect 157872 77302 158024 77330
rect 145932 77250 145984 77256
rect 140044 73160 140096 73166
rect 140044 73102 140096 73108
rect 134524 67040 134576 67046
rect 134524 66982 134576 66988
rect 123484 63028 123536 63034
rect 123484 62970 123536 62976
rect 75920 62960 75972 62966
rect 75920 62902 75972 62908
rect 71044 62892 71096 62898
rect 71044 62834 71096 62840
rect 65524 62824 65576 62830
rect 65524 62766 65576 62772
rect 57610 61704 57666 61713
rect 57610 61639 57666 61648
rect 140056 61470 140084 73102
rect 144932 61538 144960 77250
rect 144920 61532 144972 61538
rect 144920 61474 144972 61480
rect 140044 61464 140096 61470
rect 140044 61406 140096 61412
rect 102782 60752 102838 60761
rect 102782 60687 102838 60696
rect 102138 58032 102194 58041
rect 102138 57967 102140 57976
rect 102192 57967 102194 57976
rect 102140 57938 102192 57944
rect 102598 56672 102654 56681
rect 102598 56607 102654 56616
rect 57520 56568 57572 56574
rect 57520 56510 57572 56516
rect 57532 56409 57560 56510
rect 57518 56400 57574 56409
rect 57518 56335 57574 56344
rect 102138 54360 102194 54369
rect 102138 54295 102194 54304
rect 102152 53854 102180 54295
rect 102140 53848 102192 53854
rect 102140 53790 102192 53796
rect 102138 53544 102194 53553
rect 102138 53479 102194 53488
rect 102152 52698 102180 53479
rect 102140 52692 102192 52698
rect 102140 52634 102192 52640
rect 102138 52592 102194 52601
rect 102138 52527 102194 52536
rect 102152 52494 102180 52527
rect 102140 52488 102192 52494
rect 102140 52430 102192 52436
rect 57060 52420 57112 52426
rect 57060 52362 57112 52368
rect 57072 51785 57100 52362
rect 57058 51776 57114 51785
rect 57058 51711 57114 51720
rect 102138 50144 102194 50153
rect 102138 50079 102194 50088
rect 102152 49842 102180 50079
rect 102140 49836 102192 49842
rect 102140 49778 102192 49784
rect 102612 49706 102640 56607
rect 102796 52426 102824 60687
rect 102874 59664 102930 59673
rect 102874 59599 102930 59608
rect 102784 52420 102836 52426
rect 102784 52362 102836 52368
rect 102888 52358 102916 59599
rect 151832 58750 151860 77302
rect 157996 74497 158024 77302
rect 163654 77058 163682 77316
rect 169464 77302 169708 77330
rect 163654 77030 163728 77058
rect 163700 75954 163728 77030
rect 163688 75948 163740 75954
rect 163688 75890 163740 75896
rect 157982 74488 158038 74497
rect 157982 74423 158038 74432
rect 157996 58818 158024 74423
rect 163700 69834 163728 75890
rect 169680 72622 169708 77302
rect 175200 77302 175260 77330
rect 180996 77302 181056 77330
rect 186516 77302 186852 77330
rect 191852 77302 192648 77330
rect 197372 77302 198444 77330
rect 204180 77302 204240 77330
rect 210036 77302 210372 77330
rect 215832 77302 216168 77330
rect 221628 77302 221964 77330
rect 175200 73982 175228 77302
rect 180996 75886 181024 77302
rect 183468 76560 183520 76566
rect 183468 76502 183520 76508
rect 183480 75886 183508 76502
rect 186516 75886 186544 77302
rect 180984 75880 181036 75886
rect 180984 75822 181036 75828
rect 181444 75880 181496 75886
rect 181444 75822 181496 75828
rect 183468 75880 183520 75886
rect 183468 75822 183520 75828
rect 186504 75880 186556 75886
rect 186504 75822 186556 75828
rect 186964 75880 187016 75886
rect 186964 75822 187016 75828
rect 175188 73976 175240 73982
rect 175188 73918 175240 73924
rect 169668 72616 169720 72622
rect 169668 72558 169720 72564
rect 163688 69828 163740 69834
rect 163688 69770 163740 69776
rect 181456 60178 181484 75822
rect 186976 61606 187004 75822
rect 186964 61600 187016 61606
rect 186964 61542 187016 61548
rect 191852 60246 191880 77302
rect 197372 67114 197400 77302
rect 204180 75342 204208 77302
rect 204168 75336 204220 75342
rect 204168 75278 204220 75284
rect 210344 75274 210372 77302
rect 210332 75268 210384 75274
rect 210332 75210 210384 75216
rect 216140 75206 216168 77302
rect 221936 75410 221964 77302
rect 226352 77302 227424 77330
rect 232792 77302 233220 77330
rect 221924 75404 221976 75410
rect 221924 75346 221976 75352
rect 221464 75336 221516 75342
rect 221464 75278 221516 75284
rect 216128 75200 216180 75206
rect 216128 75142 216180 75148
rect 199384 70440 199436 70446
rect 199384 70382 199436 70388
rect 197360 67108 197412 67114
rect 197360 67050 197412 67056
rect 191840 60240 191892 60246
rect 191840 60182 191892 60188
rect 181444 60172 181496 60178
rect 181444 60114 181496 60120
rect 157984 58812 158036 58818
rect 157984 58754 158036 58760
rect 151820 58744 151872 58750
rect 151820 58686 151872 58692
rect 102966 58576 103022 58585
rect 102966 58511 103022 58520
rect 102876 52352 102928 52358
rect 102876 52294 102928 52300
rect 102980 51066 103008 58511
rect 104164 57996 104216 58002
rect 104164 57938 104216 57944
rect 103058 55584 103114 55593
rect 103058 55519 103114 55528
rect 102968 51060 103020 51066
rect 102968 51002 103020 51008
rect 102600 49700 102652 49706
rect 102600 49642 102652 49648
rect 102138 49192 102194 49201
rect 102138 49127 102194 49136
rect 102152 48890 102180 49127
rect 102140 48884 102192 48890
rect 102140 48826 102192 48832
rect 103072 48278 103100 55519
rect 103888 52692 103940 52698
rect 103888 52634 103940 52640
rect 103242 51096 103298 51105
rect 103242 51031 103298 51040
rect 103060 48272 103112 48278
rect 103060 48214 103112 48220
rect 102966 47696 103022 47705
rect 102966 47631 103022 47640
rect 102598 47016 102654 47025
rect 102598 46951 102654 46960
rect 57520 46912 57572 46918
rect 57518 46880 57520 46889
rect 57572 46880 57574 46889
rect 57518 46815 57574 46824
rect 60004 44192 60056 44198
rect 60004 44134 60056 44140
rect 57152 42764 57204 42770
rect 57152 42706 57204 42712
rect 57164 42129 57192 42706
rect 57150 42120 57206 42129
rect 57150 42055 57206 42064
rect 57060 37256 57112 37262
rect 57060 37198 57112 37204
rect 57072 36961 57100 37198
rect 57058 36952 57114 36961
rect 57058 36887 57114 36896
rect 57612 31748 57664 31754
rect 57612 31690 57664 31696
rect 57624 31657 57652 31690
rect 57610 31648 57666 31657
rect 57610 31583 57666 31592
rect 57244 27600 57296 27606
rect 57244 27542 57296 27548
rect 57256 27169 57284 27542
rect 57242 27160 57298 27169
rect 57242 27095 57298 27104
rect 60016 22302 60044 44134
rect 102322 43344 102378 43353
rect 102322 43279 102378 43288
rect 102138 42936 102194 42945
rect 102138 42871 102194 42880
rect 102152 40730 102180 42871
rect 102230 41440 102286 41449
rect 102230 41375 102286 41384
rect 102140 40724 102192 40730
rect 102140 40666 102192 40672
rect 102138 40080 102194 40089
rect 102138 40015 102194 40024
rect 102152 37262 102180 40015
rect 102244 38622 102272 41375
rect 102336 40050 102364 43279
rect 102612 42702 102640 46951
rect 102874 45792 102930 45801
rect 102874 45727 102930 45736
rect 102600 42696 102652 42702
rect 102600 42638 102652 42644
rect 102888 41410 102916 45727
rect 102980 42770 103008 47631
rect 103256 45558 103284 51031
rect 103900 46918 103928 52634
rect 104176 49638 104204 57938
rect 109040 53848 109092 53854
rect 109040 53790 109092 53796
rect 104440 49836 104492 49842
rect 104440 49778 104492 49784
rect 104164 49632 104216 49638
rect 104164 49574 104216 49580
rect 104348 48884 104400 48890
rect 104348 48826 104400 48832
rect 103888 46912 103940 46918
rect 103888 46854 103940 46860
rect 103244 45552 103296 45558
rect 103244 45494 103296 45500
rect 103426 44432 103482 44441
rect 103482 44390 103560 44418
rect 103426 44367 103482 44376
rect 102968 42764 103020 42770
rect 102968 42706 103020 42712
rect 102876 41404 102928 41410
rect 102876 41346 102928 41352
rect 102324 40044 102376 40050
rect 102324 39986 102376 39992
rect 103532 39982 103560 44390
rect 104360 44130 104388 48826
rect 104452 44878 104480 49778
rect 109052 48210 109080 53790
rect 196164 52488 196216 52494
rect 196164 52430 196216 52436
rect 195980 52420 196032 52426
rect 195980 52362 196032 52368
rect 195992 52329 196020 52362
rect 196072 52352 196124 52358
rect 195978 52320 196034 52329
rect 196072 52294 196124 52300
rect 195978 52255 196034 52264
rect 196084 51785 196112 52294
rect 196070 51776 196126 51785
rect 196070 51711 196126 51720
rect 195980 51060 196032 51066
rect 195980 51002 196032 51008
rect 195992 50969 196020 51002
rect 195978 50960 196034 50969
rect 195978 50895 196034 50904
rect 196072 49700 196124 49706
rect 196072 49642 196124 49648
rect 195980 49632 196032 49638
rect 195978 49600 195980 49609
rect 196032 49600 196034 49609
rect 195978 49535 196034 49544
rect 196084 49473 196112 49642
rect 196070 49464 196126 49473
rect 196070 49399 196126 49408
rect 195980 48272 196032 48278
rect 195978 48240 195980 48249
rect 196032 48240 196034 48249
rect 109040 48204 109092 48210
rect 195978 48175 196034 48184
rect 196072 48204 196124 48210
rect 109040 48146 109092 48152
rect 196072 48146 196124 48152
rect 196084 47705 196112 48146
rect 196070 47696 196126 47705
rect 196070 47631 196126 47640
rect 195980 46912 196032 46918
rect 195978 46880 195980 46889
rect 196032 46880 196034 46889
rect 195978 46815 196034 46824
rect 196176 46209 196204 52430
rect 196162 46200 196218 46209
rect 196162 46135 196218 46144
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 195992 45257 196020 45494
rect 195978 45248 196034 45257
rect 195978 45183 196034 45192
rect 104440 44872 104492 44878
rect 104440 44814 104492 44820
rect 196072 44872 196124 44878
rect 196072 44814 196124 44820
rect 196084 44169 196112 44814
rect 196070 44160 196126 44169
rect 104348 44124 104400 44130
rect 104348 44066 104400 44072
rect 195980 44124 196032 44130
rect 196070 44095 196126 44104
rect 195980 44066 196032 44072
rect 195992 43761 196020 44066
rect 195978 43752 196034 43761
rect 195978 43687 196034 43696
rect 195980 42764 196032 42770
rect 195980 42706 196032 42712
rect 195992 42537 196020 42706
rect 196072 42696 196124 42702
rect 196072 42638 196124 42644
rect 195978 42528 196034 42537
rect 195978 42463 196034 42472
rect 196084 42129 196112 42638
rect 196070 42120 196126 42129
rect 196070 42055 196126 42064
rect 195980 41404 196032 41410
rect 195980 41346 196032 41352
rect 195992 41177 196020 41346
rect 195978 41168 196034 41177
rect 195978 41103 196034 41112
rect 196164 40724 196216 40730
rect 196164 40666 196216 40672
rect 196072 40044 196124 40050
rect 196072 39986 196124 39992
rect 103520 39976 103572 39982
rect 195980 39976 196032 39982
rect 103520 39918 103572 39924
rect 195978 39944 195980 39953
rect 196032 39944 196034 39953
rect 195978 39879 196034 39888
rect 196084 39545 196112 39986
rect 196070 39536 196126 39545
rect 196070 39471 196126 39480
rect 102782 38992 102838 39001
rect 102782 38927 102838 38936
rect 102232 38616 102284 38622
rect 102232 38558 102284 38564
rect 102690 37904 102746 37913
rect 102690 37839 102746 37848
rect 102140 37256 102192 37262
rect 102140 37198 102192 37204
rect 102598 36136 102654 36145
rect 102598 36071 102654 36080
rect 102138 34640 102194 34649
rect 102138 34575 102194 34584
rect 102152 33114 102180 34575
rect 102612 34406 102640 36071
rect 102704 35834 102732 37839
rect 102796 35902 102824 38927
rect 195980 38616 196032 38622
rect 196176 38593 196204 40666
rect 195980 38558 196032 38564
rect 196162 38584 196218 38593
rect 195992 38049 196020 38558
rect 196162 38519 196218 38528
rect 195978 38040 196034 38049
rect 195978 37975 196034 37984
rect 102874 37360 102930 37369
rect 102874 37295 102930 37304
rect 102784 35896 102836 35902
rect 102784 35838 102836 35844
rect 102692 35828 102744 35834
rect 102692 35770 102744 35776
rect 102888 34474 102916 37295
rect 195980 37256 196032 37262
rect 195980 37198 196032 37204
rect 195992 37097 196020 37198
rect 195978 37088 196034 37097
rect 195978 37023 196034 37032
rect 195980 35896 196032 35902
rect 195978 35864 195980 35873
rect 196032 35864 196034 35873
rect 195978 35799 196034 35808
rect 196072 35828 196124 35834
rect 196072 35770 196124 35776
rect 196084 35465 196112 35770
rect 196070 35456 196126 35465
rect 196070 35391 196126 35400
rect 102876 34468 102928 34474
rect 102876 34410 102928 34416
rect 195980 34468 196032 34474
rect 195980 34410 196032 34416
rect 102600 34400 102652 34406
rect 195992 34377 196020 34410
rect 196072 34400 196124 34406
rect 102600 34342 102652 34348
rect 195978 34368 196034 34377
rect 196072 34342 196124 34348
rect 195978 34303 196034 34312
rect 196084 33833 196112 34342
rect 196070 33824 196126 33833
rect 196070 33759 196126 33768
rect 102322 33552 102378 33561
rect 102322 33487 102378 33496
rect 102140 33108 102192 33114
rect 102140 33050 102192 33056
rect 102138 32464 102194 32473
rect 102138 32399 102194 32408
rect 102152 31686 102180 32399
rect 102230 31784 102286 31793
rect 102336 31754 102364 33487
rect 195980 33108 196032 33114
rect 195980 33050 196032 33056
rect 195992 33017 196020 33050
rect 195978 33008 196034 33017
rect 195978 32943 196034 32952
rect 102230 31719 102286 31728
rect 102324 31748 102376 31754
rect 102140 31680 102192 31686
rect 102140 31622 102192 31628
rect 102138 30560 102194 30569
rect 102138 30495 102194 30504
rect 102152 30258 102180 30495
rect 102244 30326 102272 31719
rect 102324 31690 102376 31696
rect 195980 31748 196032 31754
rect 195980 31690 196032 31696
rect 195992 31657 196020 31690
rect 196072 31680 196124 31686
rect 195978 31648 196034 31657
rect 196072 31622 196124 31628
rect 195978 31583 196034 31592
rect 196084 31249 196112 31622
rect 196070 31240 196126 31249
rect 196070 31175 196126 31184
rect 102232 30320 102284 30326
rect 195980 30320 196032 30326
rect 102232 30262 102284 30268
rect 195978 30288 195980 30297
rect 196032 30288 196034 30297
rect 102140 30252 102192 30258
rect 195978 30223 196034 30232
rect 196072 30252 196124 30258
rect 102140 30194 102192 30200
rect 196072 30194 196124 30200
rect 196084 29753 196112 30194
rect 196070 29744 196126 29753
rect 196070 29679 196126 29688
rect 102138 29336 102194 29345
rect 102138 29271 102194 29280
rect 102152 28966 102180 29271
rect 102140 28960 102192 28966
rect 195980 28960 196032 28966
rect 102140 28902 102192 28908
rect 195978 28928 195980 28937
rect 196032 28928 196034 28937
rect 195978 28863 196034 28872
rect 102138 28520 102194 28529
rect 102138 28455 102194 28464
rect 102152 28286 102180 28455
rect 102140 28280 102192 28286
rect 102140 28222 102192 28228
rect 195980 28280 196032 28286
rect 195980 28222 196032 28228
rect 195992 28121 196020 28222
rect 195978 28112 196034 28121
rect 195978 28047 196034 28056
rect 102138 27704 102194 27713
rect 102138 27639 102194 27648
rect 102152 27606 102180 27639
rect 102140 27600 102192 27606
rect 102140 27542 102192 27548
rect 195980 27600 196032 27606
rect 195980 27542 196032 27548
rect 195992 27305 196020 27542
rect 195978 27296 196034 27305
rect 195978 27231 196034 27240
rect 102782 26344 102838 26353
rect 102782 26279 102838 26288
rect 102796 26246 102824 26279
rect 102784 26240 102836 26246
rect 195980 26240 196032 26246
rect 102784 26182 102836 26188
rect 195978 26208 195980 26217
rect 196032 26208 196034 26217
rect 195978 26143 196034 26152
rect 60004 22296 60056 22302
rect 60004 22238 60056 22244
rect 62316 22098 62344 24140
rect 66272 24126 66746 24154
rect 62304 22092 62356 22098
rect 62304 22034 62356 22040
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 3424 10328 3476 10334
rect 3424 10270 3476 10276
rect 3436 6497 3464 10270
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 66272 3466 66300 24126
rect 71148 17270 71176 24140
rect 74552 24126 75578 24154
rect 78692 24126 79994 24154
rect 84212 24126 84410 24154
rect 88352 24126 88826 24154
rect 92492 24126 93242 24154
rect 96632 24126 97658 24154
rect 71136 17264 71188 17270
rect 71136 17206 71188 17212
rect 74552 15910 74580 24126
rect 74540 15904 74592 15910
rect 74540 15846 74592 15852
rect 78692 6186 78720 24126
rect 84212 8974 84240 24126
rect 85488 23520 85540 23526
rect 85488 23462 85540 23468
rect 85500 22098 85528 23462
rect 85488 22092 85540 22098
rect 85488 22034 85540 22040
rect 84200 8968 84252 8974
rect 84200 8910 84252 8916
rect 88352 7614 88380 24126
rect 88340 7608 88392 7614
rect 88340 7550 88392 7556
rect 92492 6254 92520 24126
rect 92480 6248 92532 6254
rect 92480 6190 92532 6196
rect 78680 6180 78732 6186
rect 78680 6122 78732 6128
rect 96632 4826 96660 24126
rect 199396 22098 199424 70382
rect 220912 66904 220964 66910
rect 220912 66846 220964 66852
rect 215944 65680 215996 65686
rect 215944 65622 215996 65628
rect 202880 65544 202932 65550
rect 202880 65486 202932 65492
rect 202892 54754 202920 65486
rect 209320 64388 209372 64394
rect 209320 64330 209372 64336
rect 206008 60036 206060 60042
rect 206008 59978 206060 59984
rect 204720 57248 204772 57254
rect 204720 57190 204772 57196
rect 202892 54726 203090 54754
rect 204732 54740 204760 57190
rect 206020 54754 206048 59978
rect 208032 57316 208084 57322
rect 208032 57258 208084 57264
rect 206020 54726 206402 54754
rect 208044 54740 208072 57258
rect 209332 54754 209360 64330
rect 212632 64252 212684 64258
rect 212632 64194 212684 64200
rect 211344 57384 211396 57390
rect 211344 57326 211396 57332
rect 209332 54726 209714 54754
rect 211356 54740 211384 57326
rect 212644 54754 212672 64194
rect 214288 58676 214340 58682
rect 214288 58618 214340 58624
rect 214300 54754 214328 58618
rect 215956 54754 215984 65622
rect 219440 65612 219492 65618
rect 219440 65554 219492 65560
rect 217600 64184 217652 64190
rect 217600 64126 217652 64132
rect 217612 54754 217640 64126
rect 218058 61432 218114 61441
rect 218058 61367 218114 61376
rect 218072 57322 218100 61367
rect 218060 57316 218112 57322
rect 218060 57258 218112 57264
rect 219452 54754 219480 65554
rect 220728 58880 220780 58886
rect 220728 58822 220780 58828
rect 220740 57254 220768 58822
rect 220728 57248 220780 57254
rect 220728 57190 220780 57196
rect 220924 54754 220952 66846
rect 221476 60110 221504 75278
rect 221556 67108 221608 67114
rect 221556 67050 221608 67056
rect 221464 60104 221516 60110
rect 221464 60046 221516 60052
rect 221568 57254 221596 67050
rect 226352 62082 226380 77302
rect 231860 73976 231912 73982
rect 231860 73918 231912 73924
rect 231308 72616 231360 72622
rect 231308 72558 231360 72564
rect 231320 71738 231348 72558
rect 230848 71732 230900 71738
rect 230848 71674 230900 71680
rect 231308 71732 231360 71738
rect 231308 71674 231360 71680
rect 229192 69828 229244 69834
rect 229192 69770 229244 69776
rect 226340 62076 226392 62082
rect 226340 62018 226392 62024
rect 221740 61532 221792 61538
rect 221740 61474 221792 61480
rect 221752 57934 221780 61474
rect 222568 61464 222620 61470
rect 222568 61406 222620 61412
rect 222108 61396 222160 61402
rect 222108 61338 222160 61344
rect 221740 57928 221792 57934
rect 221740 57870 221792 57876
rect 222120 57390 222148 61338
rect 222108 57384 222160 57390
rect 222108 57326 222160 57332
rect 221556 57248 221608 57254
rect 221556 57190 221608 57196
rect 222580 54754 222608 61406
rect 227720 58812 227772 58818
rect 227720 58754 227772 58760
rect 225880 58744 225932 58750
rect 225880 58686 225932 58692
rect 224592 57928 224644 57934
rect 224592 57870 224644 57876
rect 212644 54726 213026 54754
rect 214300 54726 214682 54754
rect 215956 54726 216338 54754
rect 217612 54726 217994 54754
rect 219452 54726 219650 54754
rect 220924 54726 221306 54754
rect 222580 54726 222962 54754
rect 224604 54740 224632 57870
rect 225892 54754 225920 58686
rect 227732 54754 227760 58754
rect 229204 54754 229232 69770
rect 230860 54754 230888 71674
rect 231872 55214 231900 73918
rect 232792 64874 232820 77302
rect 235276 73982 235304 77823
rect 239016 77302 239352 77330
rect 244812 77302 245056 77330
rect 235264 73976 235316 73982
rect 235264 73918 235316 73924
rect 239324 70378 239352 77302
rect 245028 73166 245056 77302
rect 247052 74534 247080 77959
rect 250608 77302 250852 77330
rect 256404 77302 256648 77330
rect 247052 74506 247448 74534
rect 250824 74526 250852 77302
rect 252560 76560 252612 76566
rect 252560 76502 252612 76508
rect 245016 73160 245068 73166
rect 245016 73102 245068 73108
rect 239312 70372 239364 70378
rect 239312 70314 239364 70320
rect 231964 64846 232820 64874
rect 231964 58750 231992 64846
rect 236000 61600 236052 61606
rect 236000 61542 236052 61548
rect 234160 60172 234212 60178
rect 234160 60114 234212 60120
rect 231952 58744 232004 58750
rect 231952 58686 232004 58692
rect 231872 55186 232544 55214
rect 232516 54754 232544 55186
rect 234172 54754 234200 60114
rect 236012 54754 236040 61542
rect 237380 60240 237432 60246
rect 237380 60182 237432 60188
rect 244278 60208 244334 60217
rect 237392 59362 237420 60182
rect 242440 60172 242492 60178
rect 244278 60143 244334 60152
rect 242440 60114 242492 60120
rect 240782 60072 240838 60081
rect 240782 60007 240838 60016
rect 237380 59356 237432 59362
rect 237380 59298 237432 59304
rect 237392 55214 237420 59298
rect 239496 57248 239548 57254
rect 239496 57190 239548 57196
rect 237392 55186 237512 55214
rect 237484 54754 237512 55186
rect 225892 54726 226274 54754
rect 227732 54726 227930 54754
rect 229204 54726 229586 54754
rect 230860 54726 231242 54754
rect 232516 54726 232898 54754
rect 234172 54726 234554 54754
rect 236012 54726 236210 54754
rect 237484 54726 237866 54754
rect 239508 54740 239536 57190
rect 240796 54754 240824 60007
rect 242452 54754 242480 60114
rect 244292 54754 244320 60143
rect 245750 59936 245806 59945
rect 245750 59871 245806 59880
rect 245764 54754 245792 59871
rect 247420 54754 247448 74506
rect 250812 74520 250864 74526
rect 250812 74462 250864 74468
rect 251088 57520 251140 57526
rect 251088 57462 251140 57468
rect 249430 57216 249486 57225
rect 249430 57151 249486 57160
rect 240796 54726 241178 54754
rect 242452 54726 242834 54754
rect 244292 54726 244490 54754
rect 245764 54726 246146 54754
rect 247420 54726 247802 54754
rect 249444 54740 249472 57151
rect 251100 54740 251128 57462
rect 252572 54754 252600 76502
rect 256620 69018 256648 77302
rect 261772 77302 262200 77330
rect 256608 69012 256660 69018
rect 256608 68954 256660 68960
rect 255688 67040 255740 67046
rect 255688 66982 255740 66988
rect 254400 57248 254452 57254
rect 254400 57190 254452 57196
rect 252572 54726 252770 54754
rect 254412 54740 254440 57190
rect 255700 54754 255728 66982
rect 261772 64874 261800 77302
rect 263598 76528 263654 76537
rect 263598 76463 263654 76472
rect 263612 74534 263640 76463
rect 264992 74534 265020 77998
rect 269120 77988 269172 77994
rect 269120 77930 269172 77936
rect 267752 77302 267996 77330
rect 266360 76628 266412 76634
rect 266360 76570 266412 76576
rect 266372 74534 266400 76570
rect 263612 74506 264008 74534
rect 264992 74506 265664 74534
rect 266372 74506 267320 74534
rect 260852 64846 261800 64874
rect 260852 59294 260880 64846
rect 260840 59288 260892 59294
rect 260840 59230 260892 59236
rect 261576 58744 261628 58750
rect 261576 58686 261628 58692
rect 261588 57662 261616 58686
rect 261576 57656 261628 57662
rect 261576 57598 261628 57604
rect 259368 57588 259420 57594
rect 259368 57530 259420 57536
rect 257712 57452 257764 57458
rect 257712 57394 257764 57400
rect 255700 54726 256082 54754
rect 257724 54740 257752 57394
rect 259380 54740 259408 57530
rect 262678 57488 262734 57497
rect 262678 57423 262734 57432
rect 261022 57352 261078 57361
rect 261022 57287 261078 57296
rect 261036 54740 261064 57287
rect 262692 54740 262720 57423
rect 263980 54754 264008 74506
rect 265636 54754 265664 74506
rect 267292 54754 267320 74506
rect 267752 67590 267780 77302
rect 267740 67584 267792 67590
rect 267740 67526 267792 67532
rect 269132 54754 269160 77930
rect 273364 77302 273792 77330
rect 273260 75336 273312 75342
rect 273260 75278 273312 75284
rect 270592 71256 270644 71262
rect 270592 71198 270644 71204
rect 270604 54754 270632 71198
rect 272524 64320 272576 64326
rect 272524 64262 272576 64268
rect 272536 57254 272564 64262
rect 272616 57384 272668 57390
rect 272616 57326 272668 57332
rect 272524 57248 272576 57254
rect 272524 57190 272576 57196
rect 263980 54726 264362 54754
rect 265636 54726 266018 54754
rect 267292 54726 267674 54754
rect 269132 54726 269330 54754
rect 270604 54726 270986 54754
rect 272628 54740 272656 57326
rect 273272 55214 273300 75278
rect 273364 60246 273392 77302
rect 274548 75268 274600 75274
rect 274548 75210 274600 75216
rect 277400 75268 277452 75274
rect 277400 75210 277452 75216
rect 274560 73982 274588 75210
rect 274548 73976 274600 73982
rect 274548 73918 274600 73924
rect 273352 60240 273404 60246
rect 273352 60182 273404 60188
rect 275928 57316 275980 57322
rect 275928 57258 275980 57264
rect 273272 55186 273944 55214
rect 273916 54754 273944 55186
rect 273916 54726 274298 54754
rect 275940 54740 275968 57258
rect 277412 54754 277440 75210
rect 278792 58886 278820 78066
rect 284956 77302 285384 77330
rect 284208 75404 284260 75410
rect 284208 75346 284260 75352
rect 278872 75200 278924 75206
rect 278872 75142 278924 75148
rect 280160 75200 280212 75206
rect 280160 75142 280212 75148
rect 278884 74050 278912 75142
rect 280172 74534 280200 75142
rect 280172 74506 280568 74534
rect 278872 74044 278924 74050
rect 278872 73986 278924 73992
rect 278780 58880 278832 58886
rect 278780 58822 278832 58828
rect 279240 57248 279292 57254
rect 279240 57190 279292 57196
rect 277412 54726 277610 54754
rect 279252 54740 279280 57190
rect 280540 54754 280568 74506
rect 284220 74118 284248 75346
rect 284208 74112 284260 74118
rect 284208 74054 284260 74060
rect 283840 73976 283892 73982
rect 283840 73918 283892 73924
rect 282184 60104 282236 60110
rect 282184 60046 282236 60052
rect 282196 54754 282224 60046
rect 283852 54754 283880 73918
rect 284956 64874 284984 77302
rect 287152 74112 287204 74118
rect 287152 74054 287204 74060
rect 285680 74044 285732 74050
rect 285680 73986 285732 73992
rect 284312 64846 284984 64874
rect 284312 61470 284340 64846
rect 284300 61464 284352 61470
rect 284300 61406 284352 61412
rect 285692 54754 285720 73986
rect 287164 54754 287192 74054
rect 287716 71738 287744 79319
rect 287704 71732 287756 71738
rect 287704 71674 287756 71680
rect 288452 57594 288480 331842
rect 288544 315858 288572 460935
rect 288636 458046 288664 585754
rect 289084 458856 289136 458862
rect 289084 458798 289136 458804
rect 288624 458040 288676 458046
rect 288624 457982 288676 457988
rect 288532 315852 288584 315858
rect 288532 315794 288584 315800
rect 288544 204202 288572 315794
rect 288532 204196 288584 204202
rect 288532 204138 288584 204144
rect 288544 62082 288572 204138
rect 289096 78062 289124 458798
rect 289832 457910 289860 585890
rect 289820 457904 289872 457910
rect 289820 457846 289872 457852
rect 289176 457496 289228 457502
rect 289176 457438 289228 457444
rect 289188 332450 289216 457438
rect 289832 332518 289860 457846
rect 289924 457502 289952 585958
rect 290016 459202 290044 586026
rect 291292 583432 291344 583438
rect 291292 583374 291344 583380
rect 291200 583296 291252 583302
rect 291200 583238 291252 583244
rect 290096 572144 290148 572150
rect 290096 572086 290148 572092
rect 290004 459196 290056 459202
rect 290004 459138 290056 459144
rect 289912 457496 289964 457502
rect 289912 457438 289964 457444
rect 289820 332512 289872 332518
rect 289820 332454 289872 332460
rect 289176 332444 289228 332450
rect 289176 332386 289228 332392
rect 289832 332110 289860 332454
rect 290016 332382 290044 459138
rect 290108 458114 290136 572086
rect 290188 572076 290240 572082
rect 290188 572018 290240 572024
rect 290200 480254 290228 572018
rect 290200 480226 290320 480254
rect 290292 459542 290320 480226
rect 290280 459536 290332 459542
rect 290280 459478 290332 459484
rect 290096 458108 290148 458114
rect 290096 458050 290148 458056
rect 290004 332376 290056 332382
rect 290004 332318 290056 332324
rect 289820 332104 289872 332110
rect 289820 332046 289872 332052
rect 289820 331968 289872 331974
rect 289820 331910 289872 331916
rect 289728 330540 289780 330546
rect 289728 330482 289780 330488
rect 289740 313342 289768 330482
rect 289728 313336 289780 313342
rect 289728 313278 289780 313284
rect 289176 204944 289228 204950
rect 289176 204886 289228 204892
rect 289188 188902 289216 204886
rect 289176 188896 289228 188902
rect 289176 188838 289228 188844
rect 289084 78056 289136 78062
rect 289084 77998 289136 78004
rect 288532 62076 288584 62082
rect 288532 62018 288584 62024
rect 288808 62076 288860 62082
rect 288808 62018 288860 62024
rect 288440 57588 288492 57594
rect 288440 57530 288492 57536
rect 288820 54754 288848 62018
rect 289832 60178 289860 331910
rect 289912 313336 289964 313342
rect 289912 313278 289964 313284
rect 289924 204474 289952 313278
rect 290016 205018 290044 332318
rect 290108 315722 290136 458050
rect 290188 456340 290240 456346
rect 290188 456282 290240 456288
rect 290200 333305 290228 456282
rect 290186 333296 290242 333305
rect 290292 333266 290320 459478
rect 291212 459406 291240 583238
rect 291304 461378 291332 583374
rect 292764 583364 292816 583370
rect 292764 583306 292816 583312
rect 292580 583228 292632 583234
rect 292580 583170 292632 583176
rect 291384 583160 291436 583166
rect 291384 583102 291436 583108
rect 291292 461372 291344 461378
rect 291292 461314 291344 461320
rect 291396 459474 291424 583102
rect 291844 583024 291896 583030
rect 291844 582966 291896 582972
rect 291856 462602 291884 582966
rect 291844 462596 291896 462602
rect 291844 462538 291896 462544
rect 291476 462324 291528 462330
rect 291476 462266 291528 462272
rect 291488 461038 291516 462266
rect 291568 461372 291620 461378
rect 291568 461314 291620 461320
rect 291476 461032 291528 461038
rect 291476 460974 291528 460980
rect 291384 459468 291436 459474
rect 291384 459410 291436 459416
rect 291200 459400 291252 459406
rect 291200 459342 291252 459348
rect 291212 458318 291240 459342
rect 291200 458312 291252 458318
rect 291200 458254 291252 458260
rect 291396 458250 291424 459410
rect 291384 458244 291436 458250
rect 291384 458186 291436 458192
rect 291384 458040 291436 458046
rect 291384 457982 291436 457988
rect 291396 335354 291424 457982
rect 291304 335326 291424 335354
rect 290186 333231 290242 333240
rect 290280 333260 290332 333266
rect 290280 333202 290332 333208
rect 291304 332994 291332 335326
rect 291488 333334 291516 460974
rect 291476 333328 291528 333334
rect 291476 333270 291528 333276
rect 291292 332988 291344 332994
rect 291292 332930 291344 332936
rect 290556 332036 290608 332042
rect 290556 331978 290608 331984
rect 290464 331968 290516 331974
rect 290464 331910 290516 331916
rect 290096 315716 290148 315722
rect 290096 315658 290148 315664
rect 290108 314702 290136 315658
rect 290096 314696 290148 314702
rect 290096 314638 290148 314644
rect 290004 205012 290056 205018
rect 290004 204954 290056 204960
rect 289912 204468 289964 204474
rect 289912 204410 289964 204416
rect 289912 203584 289964 203590
rect 289912 203526 289964 203532
rect 289820 60172 289872 60178
rect 289820 60114 289872 60120
rect 289924 57458 289952 203526
rect 290002 202872 290058 202881
rect 290002 202807 290058 202816
rect 290016 69018 290044 202807
rect 290476 76634 290504 331910
rect 290568 78062 290596 331978
rect 291200 314696 291252 314702
rect 291200 314638 291252 314644
rect 291212 204610 291240 314638
rect 291304 209774 291332 332930
rect 291474 331800 291530 331809
rect 291474 331735 291530 331744
rect 291304 209746 291424 209774
rect 291200 204604 291252 204610
rect 291200 204546 291252 204552
rect 291200 204264 291252 204270
rect 291200 204206 291252 204212
rect 291396 204218 291424 209746
rect 291488 204338 291516 331735
rect 291580 315790 291608 461314
rect 291856 461106 291884 462538
rect 292592 462482 292620 583170
rect 292500 462454 292620 462482
rect 291844 461100 291896 461106
rect 291844 461042 291896 461048
rect 292500 460970 292528 462454
rect 292580 462392 292632 462398
rect 292580 462334 292632 462340
rect 292592 461174 292620 462334
rect 292580 461168 292632 461174
rect 292580 461110 292632 461116
rect 292488 460964 292540 460970
rect 292488 460906 292540 460912
rect 292500 334014 292528 460906
rect 292776 459338 292804 583306
rect 293960 583092 294012 583098
rect 293960 583034 294012 583040
rect 293224 580440 293276 580446
rect 293224 580382 293276 580388
rect 292948 462596 293000 462602
rect 292948 462538 293000 462544
rect 292764 459332 292816 459338
rect 292764 459274 292816 459280
rect 292672 458244 292724 458250
rect 292672 458186 292724 458192
rect 292488 334008 292540 334014
rect 292488 333950 292540 333956
rect 291752 333328 291804 333334
rect 291752 333270 291804 333276
rect 291764 332790 291792 333270
rect 291752 332784 291804 332790
rect 291752 332726 291804 332732
rect 291568 315784 291620 315790
rect 291568 315726 291620 315732
rect 291580 314702 291608 315726
rect 291568 314696 291620 314702
rect 291568 314638 291620 314644
rect 291660 204604 291712 204610
rect 291660 204546 291712 204552
rect 291476 204332 291528 204338
rect 291476 204274 291528 204280
rect 291212 203658 291240 204206
rect 291396 204190 291516 204218
rect 291384 204128 291436 204134
rect 291384 204070 291436 204076
rect 291396 203998 291424 204070
rect 291384 203992 291436 203998
rect 291384 203934 291436 203940
rect 291200 203652 291252 203658
rect 291200 203594 291252 203600
rect 290556 78056 290608 78062
rect 290556 77998 290608 78004
rect 290464 76628 290516 76634
rect 290464 76570 290516 76576
rect 290004 69012 290056 69018
rect 290004 68954 290056 68960
rect 291108 69012 291160 69018
rect 291108 68954 291160 68960
rect 291120 68610 291148 68954
rect 291108 68604 291160 68610
rect 291108 68546 291160 68552
rect 291212 57974 291240 203594
rect 291396 74050 291424 203934
rect 291488 202842 291516 204190
rect 291476 202836 291528 202842
rect 291476 202778 291528 202784
rect 291488 74526 291516 202778
rect 291568 185904 291620 185910
rect 291568 185846 291620 185852
rect 291580 79393 291608 185846
rect 291566 79384 291622 79393
rect 291566 79319 291622 79328
rect 291476 74520 291528 74526
rect 291476 74462 291528 74468
rect 291488 74050 291516 74462
rect 291384 74044 291436 74050
rect 291384 73986 291436 73992
rect 291476 74044 291528 74050
rect 291476 73986 291528 73992
rect 291672 73166 291700 204546
rect 291764 204134 291792 332726
rect 292500 332722 292528 333950
rect 292488 332716 292540 332722
rect 292488 332658 292540 332664
rect 292580 332648 292632 332654
rect 292580 332590 292632 332596
rect 291752 204128 291804 204134
rect 291752 204070 291804 204076
rect 292592 201482 292620 332590
rect 292684 330546 292712 458186
rect 292776 331158 292804 459274
rect 292856 458312 292908 458318
rect 292856 458254 292908 458260
rect 292868 333334 292896 458254
rect 292856 333328 292908 333334
rect 292856 333270 292908 333276
rect 292960 331809 292988 462538
rect 293236 462398 293264 580382
rect 293316 572008 293368 572014
rect 293316 571950 293368 571956
rect 293224 462392 293276 462398
rect 293224 462334 293276 462340
rect 293328 458250 293356 571950
rect 293972 460902 294000 583034
rect 294052 580304 294104 580310
rect 294052 580246 294104 580252
rect 294064 462330 294092 580246
rect 294604 572212 294656 572218
rect 294604 572154 294656 572160
rect 294052 462324 294104 462330
rect 294052 462266 294104 462272
rect 293960 460896 294012 460902
rect 293960 460838 294012 460844
rect 293972 459610 294000 460838
rect 293960 459604 294012 459610
rect 293960 459546 294012 459552
rect 293316 458244 293368 458250
rect 293316 458186 293368 458192
rect 293960 458244 294012 458250
rect 293960 458186 294012 458192
rect 293972 345014 294000 458186
rect 293972 344986 294092 345014
rect 294064 332858 294092 344986
rect 294052 332852 294104 332858
rect 294052 332794 294104 332800
rect 293040 332444 293092 332450
rect 293040 332386 293092 332392
rect 292946 331800 293002 331809
rect 292946 331735 293002 331744
rect 292764 331152 292816 331158
rect 292764 331094 292816 331100
rect 292672 330540 292724 330546
rect 292672 330482 292724 330488
rect 292776 204814 292804 331094
rect 292948 315376 293000 315382
rect 292948 315318 293000 315324
rect 292856 314696 292908 314702
rect 292856 314638 292908 314644
rect 292764 204808 292816 204814
rect 292764 204750 292816 204756
rect 292776 204542 292804 204750
rect 292764 204536 292816 204542
rect 292764 204478 292816 204484
rect 292868 204270 292896 314638
rect 292856 204264 292908 204270
rect 292670 204232 292726 204241
rect 292856 204206 292908 204212
rect 292670 204167 292726 204176
rect 292684 203833 292712 204167
rect 292960 204082 292988 315318
rect 293052 204241 293080 332386
rect 293960 332104 294012 332110
rect 293960 332046 294012 332052
rect 293132 205012 293184 205018
rect 293132 204954 293184 204960
rect 293038 204232 293094 204241
rect 293038 204167 293094 204176
rect 292776 204066 292988 204082
rect 292764 204060 292988 204066
rect 292816 204054 292988 204060
rect 292764 204002 292816 204008
rect 292670 203824 292726 203833
rect 292670 203759 292726 203768
rect 292580 201476 292632 201482
rect 292580 201418 292632 201424
rect 292684 74534 292712 203759
rect 292592 74506 292712 74534
rect 291660 73160 291712 73166
rect 291660 73102 291712 73108
rect 291672 72758 291700 73102
rect 291660 72752 291712 72758
rect 291660 72694 291712 72700
rect 292120 69828 292172 69834
rect 292120 69770 292172 69776
rect 291120 57946 291240 57974
rect 291120 57662 291148 57946
rect 291108 57656 291160 57662
rect 291108 57598 291160 57604
rect 289912 57452 289964 57458
rect 289912 57394 289964 57400
rect 291120 54754 291148 57598
rect 280540 54726 280922 54754
rect 282196 54726 282578 54754
rect 283852 54726 284234 54754
rect 285692 54726 285890 54754
rect 287164 54726 287546 54754
rect 288820 54726 289202 54754
rect 290858 54726 291148 54754
rect 292132 54754 292160 69770
rect 292592 67590 292620 74506
rect 292776 70378 292804 204002
rect 292948 202836 293000 202842
rect 292948 202778 293000 202784
rect 292960 202162 292988 202778
rect 292948 202156 293000 202162
rect 292948 202098 293000 202104
rect 292856 186924 292908 186930
rect 292856 186866 292908 186872
rect 292764 70372 292816 70378
rect 292764 70314 292816 70320
rect 292580 67584 292632 67590
rect 292580 67526 292632 67532
rect 292592 67114 292620 67526
rect 292580 67108 292632 67114
rect 292580 67050 292632 67056
rect 292868 60110 292896 186866
rect 292856 60104 292908 60110
rect 292856 60046 292908 60052
rect 292960 59294 292988 202098
rect 293144 78130 293172 204954
rect 293972 202842 294000 332046
rect 294064 204921 294092 332794
rect 294050 204912 294106 204921
rect 294050 204847 294106 204856
rect 294142 204232 294198 204241
rect 294142 204167 294198 204176
rect 294156 203697 294184 204167
rect 294142 203688 294198 203697
rect 294142 203623 294198 203632
rect 293960 202836 294012 202842
rect 293960 202778 294012 202784
rect 294052 186380 294104 186386
rect 294052 186322 294104 186328
rect 293132 78124 293184 78130
rect 293132 78066 293184 78072
rect 293960 72616 294012 72622
rect 293960 72558 294012 72564
rect 293500 70372 293552 70378
rect 293500 70314 293552 70320
rect 293512 69970 293540 70314
rect 293500 69964 293552 69970
rect 293500 69906 293552 69912
rect 292580 59288 292632 59294
rect 292580 59230 292632 59236
rect 292948 59288 293000 59294
rect 292948 59230 293000 59236
rect 292592 57594 292620 59230
rect 292580 57588 292632 57594
rect 292580 57530 292632 57536
rect 293972 54754 294000 72558
rect 294064 59362 294092 186322
rect 294156 73982 294184 203623
rect 294144 73976 294196 73982
rect 294144 73918 294196 73924
rect 294616 60110 294644 572154
rect 294696 458924 294748 458930
rect 294696 458866 294748 458872
rect 294604 60104 294656 60110
rect 294604 60046 294656 60052
rect 294052 59356 294104 59362
rect 294052 59298 294104 59304
rect 294708 57458 294736 458866
rect 295260 76906 295288 700470
rect 413664 700466 413692 703520
rect 462332 701010 462360 703520
rect 462320 701004 462372 701010
rect 462320 700946 462372 700952
rect 300584 700460 300636 700466
rect 300584 700402 300636 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 300596 588674 300624 700402
rect 478524 700398 478552 703520
rect 300676 700392 300728 700398
rect 300676 700334 300728 700340
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 300584 588668 300636 588674
rect 300584 588610 300636 588616
rect 300688 586566 300716 700334
rect 300768 700324 300820 700330
rect 300768 700266 300820 700272
rect 300676 586560 300728 586566
rect 300676 586502 300728 586508
rect 300492 586152 300544 586158
rect 300492 586094 300544 586100
rect 297824 585880 297876 585886
rect 297824 585822 297876 585828
rect 297732 583296 297784 583302
rect 297732 583238 297784 583244
rect 296628 583024 296680 583030
rect 296628 582966 296680 582972
rect 296536 580576 296588 580582
rect 296536 580518 296588 580524
rect 296444 580440 296496 580446
rect 296444 580382 296496 580388
rect 296456 461145 296484 580382
rect 296442 461136 296498 461145
rect 296442 461071 296498 461080
rect 295432 459604 295484 459610
rect 295432 459546 295484 459552
rect 295444 331226 295472 459546
rect 295616 334008 295668 334014
rect 295616 333950 295668 333956
rect 295432 331220 295484 331226
rect 295432 331162 295484 331168
rect 295340 204808 295392 204814
rect 295340 204750 295392 204756
rect 295248 76900 295300 76906
rect 295248 76842 295300 76848
rect 295352 74118 295380 204750
rect 295444 204406 295472 331162
rect 295524 316056 295576 316062
rect 295524 315998 295576 316004
rect 295536 204950 295564 315998
rect 295524 204944 295576 204950
rect 295524 204886 295576 204892
rect 295432 204400 295484 204406
rect 295432 204342 295484 204348
rect 295628 204241 295656 333950
rect 296260 332716 296312 332722
rect 296260 332658 296312 332664
rect 295614 204232 295670 204241
rect 295614 204167 295670 204176
rect 295984 203788 296036 203794
rect 295984 203730 296036 203736
rect 295996 76702 296024 203730
rect 296272 188426 296300 332658
rect 296456 317529 296484 461071
rect 296548 460902 296576 580518
rect 296640 462466 296668 582966
rect 296628 462460 296680 462466
rect 296628 462402 296680 462408
rect 296536 460896 296588 460902
rect 296536 460838 296588 460844
rect 296442 317520 296498 317529
rect 296442 317455 296498 317464
rect 296548 316034 296576 460838
rect 296640 333266 296668 462402
rect 296720 462392 296772 462398
rect 296720 462334 296772 462340
rect 296628 333260 296680 333266
rect 296628 333202 296680 333208
rect 296732 332654 296760 462334
rect 297744 462262 297772 583238
rect 297836 462330 297864 585822
rect 299388 585812 299440 585818
rect 299388 585754 299440 585760
rect 298836 583228 298888 583234
rect 298836 583170 298888 583176
rect 297916 583092 297968 583098
rect 297916 583034 297968 583040
rect 297824 462324 297876 462330
rect 297824 462266 297876 462272
rect 297732 462256 297784 462262
rect 297732 462198 297784 462204
rect 297928 460934 297956 583034
rect 298008 580372 298060 580378
rect 298008 580314 298060 580320
rect 297836 460906 297956 460934
rect 297836 459474 297864 460906
rect 297824 459468 297876 459474
rect 297824 459410 297876 459416
rect 297730 458280 297786 458289
rect 297730 458215 297786 458224
rect 297364 443692 297416 443698
rect 297364 443634 297416 443640
rect 296720 332648 296772 332654
rect 296720 332590 296772 332596
rect 296364 316006 296576 316034
rect 296364 315858 296392 316006
rect 296352 315852 296404 315858
rect 296352 315794 296404 315800
rect 296364 189009 296392 315794
rect 296720 313948 296772 313954
rect 296720 313890 296772 313896
rect 296536 204944 296588 204950
rect 296536 204886 296588 204892
rect 296350 189000 296406 189009
rect 296350 188935 296406 188944
rect 296444 188964 296496 188970
rect 296444 188906 296496 188912
rect 296260 188420 296312 188426
rect 296260 188362 296312 188368
rect 295984 76696 296036 76702
rect 295984 76638 296036 76644
rect 295340 74112 295392 74118
rect 295340 74054 295392 74060
rect 295432 73976 295484 73982
rect 295432 73918 295484 73924
rect 294696 57452 294748 57458
rect 294696 57394 294748 57400
rect 295444 54754 295472 73918
rect 296456 60178 296484 188906
rect 296548 73166 296576 204886
rect 296732 189038 296760 313890
rect 296720 189032 296772 189038
rect 296720 188974 296772 188980
rect 296628 187060 296680 187066
rect 296628 187002 296680 187008
rect 296536 73160 296588 73166
rect 296536 73102 296588 73108
rect 296444 60172 296496 60178
rect 296444 60114 296496 60120
rect 296640 59362 296668 187002
rect 297088 67040 297140 67046
rect 297088 66982 297140 66988
rect 296628 59356 296680 59362
rect 296628 59298 296680 59304
rect 297100 54754 297128 66982
rect 297376 57361 297404 443634
rect 297456 331900 297508 331906
rect 297456 331842 297508 331848
rect 297468 57526 297496 331842
rect 297744 316034 297772 458215
rect 297836 332722 297864 459410
rect 298020 456550 298048 580314
rect 298744 462256 298796 462262
rect 298744 462198 298796 462204
rect 298756 460970 298784 462198
rect 298744 460964 298796 460970
rect 298744 460906 298796 460912
rect 298008 456544 298060 456550
rect 298008 456486 298060 456492
rect 297916 455388 297968 455394
rect 297916 455330 297968 455336
rect 297824 332716 297876 332722
rect 297824 332658 297876 332664
rect 297928 317422 297956 455330
rect 298756 451274 298784 460906
rect 298848 458726 298876 583170
rect 299204 583160 299256 583166
rect 299204 583102 299256 583108
rect 299112 580304 299164 580310
rect 299112 580246 299164 580252
rect 299124 463593 299152 580246
rect 299110 463584 299166 463593
rect 299110 463519 299166 463528
rect 299216 460934 299244 583102
rect 299296 461168 299348 461174
rect 299296 461110 299348 461116
rect 299032 460906 299244 460934
rect 299032 459406 299060 460906
rect 299020 459400 299072 459406
rect 299020 459342 299072 459348
rect 298836 458720 298888 458726
rect 298836 458662 298888 458668
rect 298756 451246 298968 451274
rect 298836 332648 298888 332654
rect 298836 332590 298888 332596
rect 298742 317520 298798 317529
rect 298742 317455 298744 317464
rect 298796 317455 298798 317464
rect 298744 317426 298796 317432
rect 297916 317416 297968 317422
rect 297916 317358 297968 317364
rect 297744 316006 298140 316034
rect 298008 315376 298060 315382
rect 298008 315318 298060 315324
rect 297548 315308 297600 315314
rect 297548 315250 297600 315256
rect 297560 57526 297588 315250
rect 298020 205766 298048 315318
rect 298112 315314 298140 316006
rect 298100 315308 298152 315314
rect 298100 315250 298152 315256
rect 298008 205760 298060 205766
rect 298008 205702 298060 205708
rect 297640 203584 297692 203590
rect 297640 203526 297692 203532
rect 297652 76566 297680 203526
rect 298112 188970 298140 315250
rect 298848 204950 298876 332590
rect 298940 315654 298968 451246
rect 299032 332858 299060 459342
rect 299202 459232 299258 459241
rect 299202 459167 299204 459176
rect 299256 459167 299258 459176
rect 299204 459138 299256 459144
rect 299112 458244 299164 458250
rect 299112 458186 299164 458192
rect 299124 332926 299152 458186
rect 299204 456544 299256 456550
rect 299204 456486 299256 456492
rect 299112 332920 299164 332926
rect 299112 332862 299164 332868
rect 299020 332852 299072 332858
rect 299020 332794 299072 332800
rect 299032 332654 299060 332794
rect 299020 332648 299072 332654
rect 299020 332590 299072 332596
rect 299020 331288 299072 331294
rect 299020 331230 299072 331236
rect 298928 315648 298980 315654
rect 298928 315590 298980 315596
rect 298940 314702 298968 315590
rect 298928 314696 298980 314702
rect 298928 314638 298980 314644
rect 298836 204944 298888 204950
rect 298836 204886 298888 204892
rect 299032 204134 299060 331230
rect 299124 325694 299152 332862
rect 299216 330546 299244 456486
rect 299308 332450 299336 461110
rect 299400 459338 299428 585754
rect 300400 580508 300452 580514
rect 300400 580450 300452 580456
rect 300412 470594 300440 580450
rect 300136 470566 300440 470594
rect 300136 462398 300164 470566
rect 300124 462392 300176 462398
rect 300124 462334 300176 462340
rect 299388 459332 299440 459338
rect 299388 459274 299440 459280
rect 299400 458250 299428 459274
rect 299388 458244 299440 458250
rect 299388 458186 299440 458192
rect 299296 332444 299348 332450
rect 299296 332386 299348 332392
rect 299308 331294 299336 332386
rect 299296 331288 299348 331294
rect 299296 331230 299348 331236
rect 299204 330540 299256 330546
rect 299204 330482 299256 330488
rect 299124 325666 299428 325694
rect 299296 314696 299348 314702
rect 299296 314638 299348 314644
rect 299204 204264 299256 204270
rect 299204 204206 299256 204212
rect 299020 204128 299072 204134
rect 299020 204070 299072 204076
rect 299032 200114 299060 204070
rect 299032 200086 299152 200114
rect 298560 189032 298612 189038
rect 298558 189000 298560 189009
rect 298612 189000 298614 189009
rect 298100 188964 298152 188970
rect 298558 188935 298614 188944
rect 298100 188906 298152 188912
rect 298744 188420 298796 188426
rect 298744 188362 298796 188368
rect 298008 186992 298060 186998
rect 298008 186934 298060 186940
rect 297640 76560 297692 76566
rect 297640 76502 297692 76508
rect 298020 58818 298048 186934
rect 298756 69902 298784 188362
rect 299124 78266 299152 200086
rect 299112 78260 299164 78266
rect 299112 78202 299164 78208
rect 299216 76566 299244 204206
rect 299308 187610 299336 314638
rect 299400 204474 299428 325666
rect 300136 315926 300164 462334
rect 300216 462324 300268 462330
rect 300216 462266 300268 462272
rect 300228 461242 300256 462266
rect 300308 461916 300360 461922
rect 300308 461858 300360 461864
rect 300216 461236 300268 461242
rect 300216 461178 300268 461184
rect 300228 333198 300256 461178
rect 300320 461106 300348 461858
rect 300308 461100 300360 461106
rect 300308 461042 300360 461048
rect 300216 333192 300268 333198
rect 300216 333134 300268 333140
rect 300320 332518 300348 461042
rect 300504 459241 300532 586094
rect 300676 586084 300728 586090
rect 300676 586026 300728 586032
rect 300584 585948 300636 585954
rect 300584 585890 300636 585896
rect 300596 461922 300624 585890
rect 300688 462262 300716 586026
rect 300780 462330 300808 700266
rect 527192 697610 527220 703520
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 527180 697604 527232 697610
rect 527180 697546 527232 697552
rect 574100 697604 574152 697610
rect 574100 697546 574152 697552
rect 574112 696998 574140 697546
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 574100 696992 574152 696998
rect 574100 696934 574152 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 304184 588674 304566 588690
rect 304172 588668 304566 588674
rect 304224 588662 304566 588668
rect 304172 588610 304224 588616
rect 310348 586566 310376 587316
rect 310336 586560 310388 586566
rect 310336 586502 310388 586508
rect 316144 586158 316172 587316
rect 316132 586152 316184 586158
rect 316132 586094 316184 586100
rect 321940 586090 321968 587316
rect 321928 586084 321980 586090
rect 321928 586026 321980 586032
rect 327736 586022 327764 587316
rect 302148 586016 302200 586022
rect 302148 585958 302200 585964
rect 327724 586016 327776 586022
rect 327724 585958 327776 585964
rect 302160 470594 302188 585958
rect 333532 585954 333560 587316
rect 333520 585948 333572 585954
rect 333520 585890 333572 585896
rect 339328 585886 339356 587316
rect 339316 585880 339368 585886
rect 339316 585822 339368 585828
rect 345124 585818 345152 587316
rect 350920 585993 350948 587316
rect 350906 585984 350962 585993
rect 350906 585919 350962 585928
rect 345112 585812 345164 585818
rect 345112 585754 345164 585760
rect 356716 583302 356744 587316
rect 356704 583296 356756 583302
rect 356704 583238 356756 583244
rect 362512 583137 362540 587316
rect 368308 583234 368336 587316
rect 368296 583228 368348 583234
rect 368296 583170 368348 583176
rect 374104 583166 374132 587316
rect 374092 583160 374144 583166
rect 362498 583128 362554 583137
rect 374092 583102 374144 583108
rect 379900 583098 379928 587316
rect 362498 583063 362554 583072
rect 379888 583092 379940 583098
rect 379888 583034 379940 583040
rect 385696 583001 385724 587316
rect 391492 583030 391520 587316
rect 391480 583024 391532 583030
rect 385682 582992 385738 583001
rect 391480 582966 391532 582972
rect 385682 582927 385738 582936
rect 397288 580582 397316 587316
rect 397276 580576 397328 580582
rect 397276 580518 397328 580524
rect 403084 580514 403112 587316
rect 408880 586498 408908 587316
rect 414676 586498 414704 587316
rect 408868 586492 408920 586498
rect 408868 586434 408920 586440
rect 414664 586492 414716 586498
rect 414664 586434 414716 586440
rect 408880 585857 408908 586434
rect 408866 585848 408922 585857
rect 408866 585783 408922 585792
rect 403072 580508 403124 580514
rect 403072 580450 403124 580456
rect 420472 580446 420500 587316
rect 420460 580440 420512 580446
rect 420460 580382 420512 580388
rect 426268 580378 426296 587316
rect 426256 580372 426308 580378
rect 426256 580314 426308 580320
rect 432064 580310 432092 587316
rect 432052 580304 432104 580310
rect 437860 580281 437888 587316
rect 443012 587302 443670 587330
rect 432052 580246 432104 580252
rect 437846 580272 437902 580281
rect 437846 580207 437902 580216
rect 443012 572014 443040 587302
rect 449452 580310 449480 587316
rect 455248 583030 455276 587316
rect 460952 587302 461058 587330
rect 466472 587302 466854 587330
rect 455236 583024 455288 583030
rect 455236 582966 455288 582972
rect 449440 580304 449492 580310
rect 449440 580246 449492 580252
rect 460952 572082 460980 587302
rect 460940 572076 460992 572082
rect 460940 572018 460992 572024
rect 443000 572008 443052 572014
rect 466472 571985 466500 587302
rect 472636 583098 472664 587316
rect 478432 585721 478460 587316
rect 478418 585712 478474 585721
rect 478418 585647 478474 585656
rect 484228 583166 484256 587316
rect 490024 583234 490052 587316
rect 495452 587302 495834 587330
rect 490012 583228 490064 583234
rect 490012 583170 490064 583176
rect 484216 583160 484268 583166
rect 484216 583102 484268 583108
rect 472624 583092 472676 583098
rect 472624 583034 472676 583040
rect 495452 572150 495480 587302
rect 501616 583302 501644 587316
rect 507412 585818 507440 587316
rect 507400 585812 507452 585818
rect 507400 585754 507452 585760
rect 513208 583370 513236 587316
rect 519004 585721 519032 587316
rect 524800 585886 524828 587316
rect 529952 587302 530610 587330
rect 524788 585880 524840 585886
rect 524788 585822 524840 585828
rect 518990 585712 519046 585721
rect 518990 585647 519046 585656
rect 513196 583364 513248 583370
rect 513196 583306 513248 583312
rect 501604 583296 501656 583302
rect 501604 583238 501656 583244
rect 529952 572218 529980 587302
rect 536392 585954 536420 587316
rect 542188 586022 542216 587316
rect 547984 586090 548012 587316
rect 553780 586158 553808 587316
rect 559576 586226 559604 587316
rect 559564 586220 559616 586226
rect 559564 586162 559616 586168
rect 553768 586152 553820 586158
rect 553768 586094 553820 586100
rect 547972 586084 548024 586090
rect 547972 586026 548024 586032
rect 542176 586016 542228 586022
rect 542176 585958 542228 585964
rect 536380 585948 536432 585954
rect 536380 585890 536432 585896
rect 565372 585857 565400 587316
rect 569960 586220 570012 586226
rect 569960 586162 570012 586168
rect 568580 585948 568632 585954
rect 568580 585890 568632 585896
rect 565358 585848 565414 585857
rect 565358 585783 565414 585792
rect 529940 572212 529992 572218
rect 529940 572154 529992 572160
rect 495440 572144 495492 572150
rect 495440 572086 495492 572092
rect 443000 571950 443052 571956
rect 466458 571976 466514 571985
rect 466458 571911 466514 571920
rect 302068 470566 302188 470594
rect 300768 462324 300820 462330
rect 300768 462266 300820 462272
rect 300676 462256 300728 462262
rect 300676 462198 300728 462204
rect 300584 461916 300636 461922
rect 300584 461858 300636 461864
rect 302068 461174 302096 470566
rect 302238 463584 302294 463593
rect 302238 463519 302294 463528
rect 302148 462256 302200 462262
rect 302148 462198 302200 462204
rect 302056 461168 302108 461174
rect 302056 461110 302108 461116
rect 300490 459232 300546 459241
rect 300490 459167 300546 459176
rect 300400 458924 300452 458930
rect 300400 458866 300452 458872
rect 300412 458726 300440 458866
rect 300400 458720 300452 458726
rect 300400 458662 300452 458668
rect 300412 332625 300440 458662
rect 300504 345014 300532 459167
rect 302160 458833 302188 462198
rect 302146 458824 302202 458833
rect 302146 458759 302202 458768
rect 300504 344986 300624 345014
rect 300398 332616 300454 332625
rect 300398 332551 300454 332560
rect 300308 332512 300360 332518
rect 300308 332454 300360 332460
rect 300124 315920 300176 315926
rect 300124 315862 300176 315868
rect 300136 315110 300164 315862
rect 300124 315104 300176 315110
rect 300124 315046 300176 315052
rect 299388 204468 299440 204474
rect 299388 204410 299440 204416
rect 299296 187604 299348 187610
rect 299296 187546 299348 187552
rect 299204 76560 299256 76566
rect 299204 76502 299256 76508
rect 299308 72690 299336 187546
rect 299296 72684 299348 72690
rect 299296 72626 299348 72632
rect 298744 69896 298796 69902
rect 298744 69838 298796 69844
rect 298744 68536 298796 68542
rect 298744 68478 298796 68484
rect 298008 58812 298060 58818
rect 298008 58754 298060 58760
rect 297456 57520 297508 57526
rect 297456 57462 297508 57468
rect 297548 57520 297600 57526
rect 297548 57462 297600 57468
rect 297362 57352 297418 57361
rect 297362 57287 297418 57296
rect 298756 54754 298784 68478
rect 299400 57934 299428 204410
rect 300320 204202 300348 332454
rect 300596 332314 300624 344986
rect 300768 333192 300820 333198
rect 300768 333134 300820 333140
rect 300780 332994 300808 333134
rect 300768 332988 300820 332994
rect 300768 332930 300820 332936
rect 300584 332308 300636 332314
rect 300584 332250 300636 332256
rect 300400 315104 300452 315110
rect 300400 315046 300452 315052
rect 300412 206650 300440 315046
rect 300400 206644 300452 206650
rect 300400 206586 300452 206592
rect 300308 204196 300360 204202
rect 300308 204138 300360 204144
rect 300216 203720 300268 203726
rect 300216 203662 300268 203668
rect 300124 203652 300176 203658
rect 300124 203594 300176 203600
rect 300136 77994 300164 203594
rect 300228 78130 300256 203662
rect 300320 200114 300348 204138
rect 300596 203998 300624 332250
rect 300674 314800 300730 314809
rect 300674 314735 300730 314744
rect 300584 203992 300636 203998
rect 300584 203934 300636 203940
rect 300320 200086 300532 200114
rect 300504 78198 300532 200086
rect 300596 78334 300624 203934
rect 300688 190454 300716 314735
rect 300780 204270 300808 332930
rect 302056 332784 302108 332790
rect 302056 332726 302108 332732
rect 302068 332625 302096 332726
rect 302054 332616 302110 332625
rect 302054 332551 302110 332560
rect 302160 332382 302188 458759
rect 302252 455394 302280 463519
rect 391216 462466 391506 462482
rect 391204 462460 391506 462466
rect 391256 462454 391506 462460
rect 437874 462466 438256 462482
rect 437874 462460 438268 462466
rect 437874 462454 438216 462460
rect 391204 462402 391256 462408
rect 438216 462402 438268 462408
rect 402888 462392 402940 462398
rect 443736 462392 443788 462398
rect 402940 462340 403098 462346
rect 402888 462334 403098 462340
rect 304172 462324 304224 462330
rect 402900 462318 403098 462334
rect 443670 462340 443736 462346
rect 443670 462334 443788 462340
rect 443670 462318 443776 462334
rect 304172 462266 304224 462272
rect 304184 462210 304212 462266
rect 304184 462182 304566 462210
rect 455262 461378 455368 461394
rect 455262 461372 455380 461378
rect 455262 461366 455328 461372
rect 455328 461314 455380 461320
rect 567108 461372 567160 461378
rect 567108 461314 567160 461320
rect 513288 461304 513340 461310
rect 306378 461136 306434 461145
rect 306378 461071 306434 461080
rect 303528 461032 303580 461038
rect 303526 461000 303528 461009
rect 303580 461000 303582 461009
rect 303526 460935 303582 460944
rect 305000 459264 305052 459270
rect 304998 459232 305000 459241
rect 305052 459232 305054 459241
rect 304998 459167 305054 459176
rect 305000 457496 305052 457502
rect 305000 457438 305052 457444
rect 305012 456550 305040 457438
rect 306392 456754 306420 461071
rect 310348 459513 310376 461244
rect 310334 459504 310390 459513
rect 310334 459439 310390 459448
rect 316144 459270 316172 461244
rect 321940 459542 321968 461244
rect 327368 461230 327750 461258
rect 327368 461174 327396 461230
rect 327356 461168 327408 461174
rect 327356 461110 327408 461116
rect 333532 461106 333560 461244
rect 336740 461236 336792 461242
rect 336740 461178 336792 461184
rect 333520 461100 333572 461106
rect 333520 461042 333572 461048
rect 336752 459542 336780 461178
rect 339328 459542 339356 461244
rect 318800 459536 318852 459542
rect 318800 459478 318852 459484
rect 321928 459536 321980 459542
rect 321928 459478 321980 459484
rect 336740 459536 336792 459542
rect 336740 459478 336792 459484
rect 339316 459536 339368 459542
rect 339316 459478 339368 459484
rect 316132 459264 316184 459270
rect 316132 459206 316184 459212
rect 318812 458833 318840 459478
rect 345124 459338 345152 461244
rect 350920 461038 350948 461244
rect 350908 461032 350960 461038
rect 350908 460974 350960 460980
rect 356716 460970 356744 461244
rect 362512 461009 362540 461244
rect 362498 461000 362554 461009
rect 356704 460964 356756 460970
rect 362498 460935 362554 460944
rect 356704 460906 356756 460912
rect 345112 459332 345164 459338
rect 345112 459274 345164 459280
rect 368308 458930 368336 461244
rect 374104 459406 374132 461244
rect 379900 459474 379928 461244
rect 379888 459468 379940 459474
rect 379888 459410 379940 459416
rect 374092 459400 374144 459406
rect 374092 459342 374144 459348
rect 385696 459202 385724 461244
rect 397288 460902 397316 461244
rect 397276 460896 397328 460902
rect 397276 460838 397328 460844
rect 408880 459542 408908 461244
rect 414676 459542 414704 461244
rect 408868 459536 408920 459542
rect 408868 459478 408920 459484
rect 414664 459536 414716 459542
rect 414664 459478 414716 459484
rect 385684 459196 385736 459202
rect 385684 459138 385736 459144
rect 368296 458924 368348 458930
rect 368296 458866 368348 458872
rect 408880 458862 408908 459478
rect 408868 458856 408920 458862
rect 318798 458824 318854 458833
rect 408868 458798 408920 458804
rect 318798 458759 318854 458768
rect 420472 456754 420500 461244
rect 426282 461230 426388 461258
rect 426360 458266 426388 461230
rect 426360 458238 426480 458266
rect 426452 457502 426480 458238
rect 426440 457496 426492 457502
rect 426440 457438 426492 457444
rect 306380 456748 306432 456754
rect 306380 456690 306432 456696
rect 420460 456748 420512 456754
rect 420460 456690 420512 456696
rect 305000 456544 305052 456550
rect 305000 456486 305052 456492
rect 432064 456074 432092 461244
rect 449452 460970 449480 461244
rect 449440 460964 449492 460970
rect 449440 460906 449492 460912
rect 461044 460902 461072 461244
rect 461032 460896 461084 460902
rect 461032 460838 461084 460844
rect 466840 459542 466868 461244
rect 471992 461230 472650 461258
rect 477512 461230 478446 461258
rect 466828 459536 466880 459542
rect 466828 459478 466880 459484
rect 307668 456068 307720 456074
rect 307668 456010 307720 456016
rect 432052 456068 432104 456074
rect 432052 456010 432104 456016
rect 307680 455394 307708 456010
rect 302240 455388 302292 455394
rect 302240 455330 302292 455336
rect 307668 455388 307720 455394
rect 307668 455330 307720 455336
rect 471992 444378 472020 461230
rect 477512 444961 477540 461230
rect 484228 461106 484256 461244
rect 484216 461100 484268 461106
rect 484216 461042 484268 461048
rect 490024 459202 490052 461244
rect 490012 459196 490064 459202
rect 490012 459138 490064 459144
rect 495820 458862 495848 461244
rect 501630 461230 501920 461258
rect 507426 461242 507808 461258
rect 513222 461252 513288 461258
rect 513222 461246 513340 461252
rect 507426 461236 507820 461242
rect 507426 461230 507768 461236
rect 501892 461174 501920 461230
rect 513222 461230 513328 461246
rect 507768 461178 507820 461184
rect 501880 461168 501932 461174
rect 501880 461110 501932 461116
rect 495808 458856 495860 458862
rect 495808 458798 495860 458804
rect 519004 458182 519032 461244
rect 524800 459406 524828 461244
rect 524788 459400 524840 459406
rect 524788 459342 524840 459348
rect 530596 459338 530624 461244
rect 530584 459332 530636 459338
rect 530584 459274 530636 459280
rect 518992 458176 519044 458182
rect 518992 458118 519044 458124
rect 536392 458114 536420 461244
rect 536380 458108 536432 458114
rect 536380 458050 536432 458056
rect 542188 458046 542216 461244
rect 547984 459270 548012 461244
rect 547972 459264 548024 459270
rect 547972 459206 548024 459212
rect 553780 458833 553808 461244
rect 559576 459474 559604 461244
rect 561588 461032 561640 461038
rect 561588 460974 561640 460980
rect 559564 459468 559616 459474
rect 559564 459410 559616 459416
rect 561600 459202 561628 460974
rect 561588 459196 561640 459202
rect 561588 459138 561640 459144
rect 553766 458824 553822 458833
rect 553766 458759 553822 458768
rect 565372 458250 565400 461244
rect 565360 458244 565412 458250
rect 565360 458186 565412 458192
rect 565820 458176 565872 458182
rect 565818 458144 565820 458153
rect 565872 458144 565874 458153
rect 565818 458079 565874 458088
rect 542176 458040 542228 458046
rect 542176 457982 542228 457988
rect 477498 444952 477554 444961
rect 477498 444887 477554 444896
rect 471980 444372 472032 444378
rect 471980 444314 472032 444320
rect 567120 443698 567148 461314
rect 567752 461236 567804 461242
rect 567752 461178 567804 461184
rect 567764 461145 567792 461178
rect 567750 461136 567806 461145
rect 567750 461071 567806 461080
rect 568592 460934 568620 585890
rect 569316 585880 569368 585886
rect 569316 585822 569368 585828
rect 568672 585812 568724 585818
rect 568672 585754 568724 585760
rect 568684 461242 568712 585754
rect 569224 485104 569276 485110
rect 569224 485046 569276 485052
rect 568762 463584 568818 463593
rect 568762 463519 568818 463528
rect 568776 462466 568804 463519
rect 568764 462460 568816 462466
rect 568764 462402 568816 462408
rect 568672 461236 568724 461242
rect 568672 461178 568724 461184
rect 568592 460906 568712 460934
rect 567936 459536 567988 459542
rect 567936 459478 567988 459484
rect 568488 459536 568540 459542
rect 568488 459478 568540 459484
rect 567948 459377 567976 459478
rect 567934 459368 567990 459377
rect 567934 459303 567990 459312
rect 568500 458561 568528 459478
rect 568486 458552 568542 458561
rect 568486 458487 568542 458496
rect 568684 458114 568712 460906
rect 568948 458244 569000 458250
rect 568948 458186 569000 458192
rect 568672 458108 568724 458114
rect 568672 458050 568724 458056
rect 567108 443692 567160 443698
rect 567108 443634 567160 443640
rect 304552 332654 304580 333268
rect 306380 333260 306432 333266
rect 306380 333202 306432 333208
rect 304540 332648 304592 332654
rect 304540 332590 304592 332596
rect 302148 332376 302200 332382
rect 302148 332318 302200 332324
rect 302054 315752 302110 315761
rect 302054 315687 302056 315696
rect 302108 315687 302110 315696
rect 302056 315658 302108 315664
rect 302054 204776 302110 204785
rect 302054 204711 302110 204720
rect 302068 204406 302096 204711
rect 302056 204400 302108 204406
rect 302056 204342 302108 204348
rect 300768 204264 300820 204270
rect 300768 204206 300820 204212
rect 302160 204066 302188 332318
rect 303528 332240 303580 332246
rect 303526 332208 303528 332217
rect 303580 332208 303582 332217
rect 303526 332143 303582 332152
rect 305000 317484 305052 317490
rect 305000 317426 305052 317432
rect 305012 315994 305040 317426
rect 305000 315988 305052 315994
rect 305000 315930 305052 315936
rect 306392 315382 306420 333202
rect 310348 332489 310376 333268
rect 310334 332480 310390 332489
rect 310334 332415 310390 332424
rect 316144 332314 316172 333268
rect 321940 332382 321968 333268
rect 327736 332450 327764 333268
rect 333532 332518 333560 333268
rect 338960 333254 339342 333282
rect 338960 332994 338988 333254
rect 338948 332988 339000 332994
rect 338948 332930 339000 332936
rect 342260 332920 342312 332926
rect 342260 332862 342312 332868
rect 342272 332586 342300 332862
rect 345124 332586 345152 333268
rect 342260 332580 342312 332586
rect 342260 332522 342312 332528
rect 345112 332580 345164 332586
rect 345112 332522 345164 332528
rect 333520 332512 333572 332518
rect 333520 332454 333572 332460
rect 327724 332444 327776 332450
rect 327724 332386 327776 332392
rect 321928 332376 321980 332382
rect 321928 332318 321980 332324
rect 316132 332308 316184 332314
rect 316132 332250 316184 332256
rect 350920 332246 350948 333268
rect 356072 333254 356730 333282
rect 361592 333254 362526 333282
rect 350908 332240 350960 332246
rect 350908 332182 350960 332188
rect 307668 330540 307720 330546
rect 307668 330482 307720 330488
rect 307680 329798 307708 330482
rect 307668 329792 307720 329798
rect 307668 329734 307720 329740
rect 307668 318096 307720 318102
rect 307668 318038 307720 318044
rect 307680 317422 307708 318038
rect 307668 317416 307720 317422
rect 307668 317358 307720 317364
rect 307668 315784 307720 315790
rect 307668 315726 307720 315732
rect 307680 315382 307708 315726
rect 356072 315654 356100 333254
rect 361592 315722 361620 333254
rect 368308 332790 368336 333268
rect 373920 333254 374118 333282
rect 373920 332858 373948 333254
rect 373908 332852 373960 332858
rect 373908 332794 373960 332800
rect 368296 332784 368348 332790
rect 368296 332726 368348 332732
rect 379900 332722 379928 333268
rect 385052 333254 385710 333282
rect 390572 333254 391506 333282
rect 396092 333254 397302 333282
rect 402992 333254 403098 333282
rect 379888 332716 379940 332722
rect 379888 332658 379940 332664
rect 361580 315716 361632 315722
rect 361580 315658 361632 315664
rect 356060 315648 356112 315654
rect 356060 315590 356112 315596
rect 306380 315376 306432 315382
rect 306380 315318 306432 315324
rect 307668 315376 307720 315382
rect 307668 315318 307720 315324
rect 385052 315314 385080 333254
rect 390572 315790 390600 333254
rect 396092 315858 396120 333254
rect 402992 315926 403020 333254
rect 408880 332586 408908 333268
rect 414676 332586 414704 333268
rect 419552 333254 420486 333282
rect 408868 332580 408920 332586
rect 408868 332522 408920 332528
rect 414664 332580 414716 332586
rect 414664 332522 414716 332528
rect 408880 331974 408908 332522
rect 408868 331968 408920 331974
rect 408868 331910 408920 331916
rect 419552 315994 419580 333254
rect 426268 329798 426296 333268
rect 431972 333254 432078 333282
rect 437492 333254 437874 333282
rect 425704 329792 425756 329798
rect 425704 329734 425756 329740
rect 426256 329792 426308 329798
rect 426256 329734 426308 329740
rect 425716 316742 425744 329734
rect 431972 318102 432000 333254
rect 437492 318170 437520 333254
rect 443656 331974 443684 333268
rect 448532 333254 449466 333282
rect 443644 331968 443696 331974
rect 443644 331910 443696 331916
rect 437480 318164 437532 318170
rect 437480 318106 437532 318112
rect 431960 318096 432012 318102
rect 431960 318038 432012 318044
rect 425704 316736 425756 316742
rect 425704 316678 425756 316684
rect 448532 315994 448560 333254
rect 455248 331294 455276 333268
rect 453948 331288 454000 331294
rect 453948 331230 454000 331236
rect 455236 331288 455288 331294
rect 455236 331230 455288 331236
rect 419540 315988 419592 315994
rect 419540 315930 419592 315936
rect 448520 315988 448572 315994
rect 448520 315930 448572 315936
rect 402980 315920 403032 315926
rect 402980 315862 403032 315868
rect 396080 315852 396132 315858
rect 396080 315794 396132 315800
rect 390560 315784 390612 315790
rect 390560 315726 390612 315732
rect 385040 315308 385092 315314
rect 385040 315250 385092 315256
rect 453960 314634 453988 331230
rect 461044 329798 461072 333268
rect 466472 333254 466854 333282
rect 461032 329792 461084 329798
rect 461032 329734 461084 329740
rect 466472 315314 466500 333254
rect 472636 332722 472664 333268
rect 472624 332716 472676 332722
rect 472624 332658 472676 332664
rect 478432 331906 478460 333268
rect 478420 331900 478472 331906
rect 478420 331842 478472 331848
rect 484228 331294 484256 333268
rect 482928 331288 482980 331294
rect 482928 331230 482980 331236
rect 484216 331288 484268 331294
rect 484216 331230 484268 331236
rect 482940 315926 482968 331230
rect 490024 329730 490052 333268
rect 495452 333254 495834 333282
rect 500972 333254 501630 333282
rect 506492 333254 507426 333282
rect 490012 329724 490064 329730
rect 490012 329666 490064 329672
rect 482928 315920 482980 315926
rect 482928 315862 482980 315868
rect 495452 315858 495480 333254
rect 500972 331242 501000 333254
rect 500880 331214 501000 331242
rect 495440 315852 495492 315858
rect 495440 315794 495492 315800
rect 500880 315790 500908 331214
rect 500868 315784 500920 315790
rect 500868 315726 500920 315732
rect 506492 315722 506520 333254
rect 513208 332790 513236 333268
rect 513196 332784 513248 332790
rect 513196 332726 513248 332732
rect 519004 332518 519032 333268
rect 524800 332586 524828 333268
rect 529952 333254 530610 333282
rect 524788 332580 524840 332586
rect 524788 332522 524840 332528
rect 518992 332512 519044 332518
rect 518992 332454 519044 332460
rect 506480 315716 506532 315722
rect 506480 315658 506532 315664
rect 529952 315654 529980 333254
rect 536392 332450 536420 333268
rect 536380 332444 536432 332450
rect 536380 332386 536432 332392
rect 542188 332382 542216 333268
rect 542176 332376 542228 332382
rect 542176 332318 542228 332324
rect 547984 332314 548012 333268
rect 547972 332308 548024 332314
rect 547972 332250 548024 332256
rect 553780 331809 553808 333268
rect 559576 332246 559604 333268
rect 559564 332240 559616 332246
rect 559564 332182 559616 332188
rect 561588 331968 561640 331974
rect 561588 331910 561640 331916
rect 553766 331800 553822 331809
rect 553766 331735 553822 331744
rect 561600 331226 561628 331910
rect 565372 331906 565400 333268
rect 567108 333260 567160 333266
rect 567108 333202 567160 333208
rect 565820 332512 565872 332518
rect 565820 332454 565872 332460
rect 565832 332353 565860 332454
rect 565818 332344 565874 332353
rect 565818 332279 565874 332288
rect 565360 331900 565412 331906
rect 565360 331842 565412 331848
rect 561588 331220 561640 331226
rect 561588 331162 561640 331168
rect 562324 318164 562376 318170
rect 562324 318106 562376 318112
rect 562336 317422 562364 318106
rect 562324 317416 562376 317422
rect 562324 317358 562376 317364
rect 565820 316736 565872 316742
rect 565820 316678 565872 316684
rect 529940 315648 529992 315654
rect 529940 315590 529992 315596
rect 466460 315308 466512 315314
rect 466460 315250 466512 315256
rect 453948 314628 454000 314634
rect 453948 314570 454000 314576
rect 565832 313954 565860 316678
rect 567120 315926 567148 333202
rect 568684 332450 568712 458050
rect 568672 332444 568724 332450
rect 568672 332386 568724 332392
rect 567108 315920 567160 315926
rect 567108 315862 567160 315868
rect 567120 314702 567148 315862
rect 567474 315752 567530 315761
rect 567474 315687 567476 315696
rect 567528 315687 567530 315696
rect 567476 315658 567528 315664
rect 567108 314696 567160 314702
rect 567108 314638 567160 314644
rect 568486 314664 568542 314673
rect 568486 314599 568488 314608
rect 568540 314599 568542 314608
rect 568488 314570 568540 314576
rect 565820 313948 565872 313954
rect 565820 313890 565872 313896
rect 307024 206644 307076 206650
rect 307024 206586 307076 206592
rect 305000 205760 305052 205766
rect 305000 205702 305052 205708
rect 302884 205692 302936 205698
rect 302884 205634 302936 205640
rect 302148 204060 302200 204066
rect 302148 204002 302200 204008
rect 300688 190426 300808 190454
rect 300780 187678 300808 190426
rect 300768 187672 300820 187678
rect 300768 187614 300820 187620
rect 300584 78328 300636 78334
rect 300584 78270 300636 78276
rect 300492 78192 300544 78198
rect 300492 78134 300544 78140
rect 300216 78124 300268 78130
rect 300216 78066 300268 78072
rect 300124 77988 300176 77994
rect 300124 77930 300176 77936
rect 300400 71188 300452 71194
rect 300400 71130 300452 71136
rect 299388 57928 299440 57934
rect 299388 57870 299440 57876
rect 300412 54754 300440 71130
rect 300780 61538 300808 187614
rect 302160 78402 302188 204002
rect 302896 186425 302924 205634
rect 304264 204332 304316 204338
rect 304264 204274 304316 204280
rect 303712 202156 303764 202162
rect 303712 202098 303764 202104
rect 303528 201476 303580 201482
rect 303528 201418 303580 201424
rect 303540 201385 303568 201418
rect 303526 201376 303582 201385
rect 303526 201311 303582 201320
rect 302882 186416 302938 186425
rect 302882 186351 302938 186360
rect 303724 185609 303752 202098
rect 304276 187066 304304 204274
rect 304552 204241 304580 205292
rect 305012 204338 305040 205702
rect 305000 204332 305052 204338
rect 305000 204274 305052 204280
rect 304538 204232 304594 204241
rect 304538 204167 304594 204176
rect 307036 188358 307064 206586
rect 560208 206372 560260 206378
rect 560208 206314 560260 206320
rect 495440 206304 495492 206310
rect 495440 206246 495492 206252
rect 310428 205692 310480 205698
rect 310428 205634 310480 205640
rect 310348 204105 310376 205292
rect 310334 204096 310390 204105
rect 310334 204031 310390 204040
rect 310440 202842 310468 205634
rect 316144 203998 316172 205292
rect 321940 204066 321968 205292
rect 327736 204134 327764 205292
rect 333532 204202 333560 205292
rect 339328 204270 339356 205292
rect 340880 204468 340932 204474
rect 340880 204410 340932 204416
rect 340892 204270 340920 204410
rect 345124 204270 345152 205292
rect 339316 204264 339368 204270
rect 339316 204206 339368 204212
rect 340880 204264 340932 204270
rect 340880 204206 340932 204212
rect 345112 204264 345164 204270
rect 345112 204206 345164 204212
rect 333520 204196 333572 204202
rect 333520 204138 333572 204144
rect 327724 204128 327776 204134
rect 327724 204070 327776 204076
rect 321928 204060 321980 204066
rect 321928 204002 321980 204008
rect 316132 203992 316184 203998
rect 316132 203934 316184 203940
rect 310428 202836 310480 202842
rect 310428 202778 310480 202784
rect 350920 201482 350948 205292
rect 356072 205278 356730 205306
rect 361592 205278 362526 205306
rect 350908 201476 350960 201482
rect 350908 201418 350960 201424
rect 307024 188352 307076 188358
rect 307024 188294 307076 188300
rect 308036 188352 308088 188358
rect 308036 188294 308088 188300
rect 304264 187060 304316 187066
rect 304264 187002 304316 187008
rect 308048 186998 308076 188294
rect 356072 187610 356100 205278
rect 361592 187678 361620 205278
rect 366272 204400 366324 204406
rect 366272 204342 366324 204348
rect 366284 204270 366312 204342
rect 368308 204270 368336 205292
rect 374012 205278 374118 205306
rect 379532 205278 379914 205306
rect 385052 205278 385710 205306
rect 374012 204950 374040 205278
rect 374000 204944 374052 204950
rect 374000 204886 374052 204892
rect 366272 204264 366324 204270
rect 366272 204206 366324 204212
rect 368296 204264 368348 204270
rect 368296 204206 368348 204212
rect 379532 188426 379560 205278
rect 385052 188970 385080 205278
rect 391492 204338 391520 205292
rect 396092 205278 397302 205306
rect 402992 205278 403098 205306
rect 391480 204332 391532 204338
rect 391480 204274 391532 204280
rect 396092 189038 396120 205278
rect 396080 189032 396132 189038
rect 396080 188974 396132 188980
rect 385040 188964 385092 188970
rect 385040 188906 385092 188912
rect 379520 188420 379572 188426
rect 379520 188362 379572 188368
rect 402992 188358 403020 205278
rect 408880 204270 408908 205292
rect 414676 204270 414704 205292
rect 419552 205278 420486 205306
rect 408868 204264 408920 204270
rect 408868 204206 408920 204212
rect 414664 204264 414716 204270
rect 414664 204206 414716 204212
rect 408880 203658 408908 204206
rect 408868 203652 408920 203658
rect 408868 203594 408920 203600
rect 419552 189009 419580 205278
rect 426268 204202 426296 205292
rect 426256 204196 426308 204202
rect 426256 204138 426308 204144
rect 426268 202842 426296 204138
rect 432064 204066 432092 205292
rect 437492 205278 437874 205306
rect 443012 205278 443670 205306
rect 448532 205278 449466 205306
rect 454052 205278 455262 205306
rect 460952 205278 461058 205306
rect 466854 205278 467144 205306
rect 432052 204060 432104 204066
rect 432052 204002 432104 204008
rect 426256 202836 426308 202842
rect 426256 202778 426308 202784
rect 432064 202162 432092 204002
rect 432052 202156 432104 202162
rect 432052 202098 432104 202104
rect 437492 189038 437520 205278
rect 443012 202994 443040 205278
rect 442920 202966 443040 202994
rect 437480 189032 437532 189038
rect 419538 189000 419594 189009
rect 437480 188974 437532 188980
rect 442920 188970 442948 202966
rect 419538 188935 419594 188944
rect 442908 188964 442960 188970
rect 402980 188352 403032 188358
rect 402980 188294 403032 188300
rect 361580 187672 361632 187678
rect 361580 187614 361632 187620
rect 356060 187604 356112 187610
rect 356060 187546 356112 187552
rect 419552 186998 419580 188935
rect 442908 188906 442960 188912
rect 448532 188358 448560 205278
rect 454052 188834 454080 205278
rect 460952 188902 460980 205278
rect 467116 204950 467144 205278
rect 467104 204944 467156 204950
rect 467104 204886 467156 204892
rect 472636 202910 472664 205292
rect 478432 203590 478460 205292
rect 483032 205278 484242 205306
rect 478420 203584 478472 203590
rect 478420 203526 478472 203532
rect 471888 202904 471940 202910
rect 471888 202846 471940 202852
rect 472624 202904 472676 202910
rect 472624 202846 472676 202852
rect 460940 188896 460992 188902
rect 460940 188838 460992 188844
rect 454040 188828 454092 188834
rect 454040 188770 454092 188776
rect 471900 188766 471928 202846
rect 471888 188760 471940 188766
rect 471888 188702 471940 188708
rect 483032 188698 483060 205278
rect 490024 200802 490052 205292
rect 495452 204202 495480 206246
rect 495820 204270 495848 205292
rect 495808 204264 495860 204270
rect 495808 204206 495860 204212
rect 495440 204196 495492 204202
rect 495440 204138 495492 204144
rect 501616 201482 501644 205292
rect 507412 204338 507440 205292
rect 513208 204406 513236 205292
rect 518912 205278 519018 205306
rect 513196 204400 513248 204406
rect 513196 204342 513248 204348
rect 507400 204332 507452 204338
rect 507400 204274 507452 204280
rect 518912 202874 518940 205278
rect 524800 204202 524828 205292
rect 530610 205278 530992 205306
rect 530964 204542 530992 205278
rect 530952 204536 531004 204542
rect 530952 204478 531004 204484
rect 524788 204196 524840 204202
rect 524788 204138 524840 204144
rect 536392 204134 536420 205292
rect 540888 205012 540940 205018
rect 540888 204954 540940 204960
rect 536380 204128 536432 204134
rect 536380 204070 536432 204076
rect 540900 204066 540928 204954
rect 542188 204270 542216 205292
rect 542176 204264 542228 204270
rect 542176 204206 542228 204212
rect 547984 204066 548012 205292
rect 540888 204060 540940 204066
rect 540888 204002 540940 204008
rect 547972 204060 548024 204066
rect 547972 204002 548024 204008
rect 553780 203590 553808 205292
rect 559576 203998 559604 205292
rect 559564 203992 559616 203998
rect 559564 203934 559616 203940
rect 553768 203584 553820 203590
rect 553768 203526 553820 203532
rect 518820 202846 518940 202874
rect 501604 201476 501656 201482
rect 501604 201418 501656 201424
rect 490012 200796 490064 200802
rect 490012 200738 490064 200744
rect 483020 188692 483072 188698
rect 483020 188634 483072 188640
rect 448520 188352 448572 188358
rect 448520 188294 448572 188300
rect 518820 187649 518848 202846
rect 560220 188834 560248 206314
rect 565372 203658 565400 205292
rect 567290 204368 567346 204377
rect 567290 204303 567292 204312
rect 567344 204303 567346 204312
rect 567292 204274 567344 204280
rect 568684 204134 568712 332386
rect 568856 314696 568908 314702
rect 568856 314638 568908 314644
rect 568764 204400 568816 204406
rect 568764 204342 568816 204348
rect 568672 204128 568724 204134
rect 568672 204070 568724 204076
rect 565360 203652 565412 203658
rect 565360 203594 565412 203600
rect 560208 188828 560260 188834
rect 560208 188770 560260 188776
rect 560220 188426 560248 188770
rect 560208 188420 560260 188426
rect 560208 188362 560260 188368
rect 518806 187640 518862 187649
rect 518806 187575 518862 187584
rect 308036 186992 308088 186998
rect 308036 186934 308088 186940
rect 419540 186992 419592 186998
rect 419540 186934 419592 186940
rect 303710 185600 303766 185609
rect 303710 185535 303766 185544
rect 302330 79928 302386 79937
rect 302330 79863 302386 79872
rect 302148 78396 302200 78402
rect 302148 78338 302200 78344
rect 302240 69964 302292 69970
rect 302240 69906 302292 69912
rect 300768 61532 300820 61538
rect 300768 61474 300820 61480
rect 302252 54754 302280 69906
rect 302344 64870 302372 79863
rect 313280 78396 313332 78402
rect 313280 78338 313332 78344
rect 310362 77994 310468 78010
rect 310362 77988 310480 77994
rect 310362 77982 310428 77988
rect 310428 77930 310480 77936
rect 304552 75993 304580 77316
rect 304538 75984 304594 75993
rect 304538 75919 304594 75928
rect 313292 75886 313320 78338
rect 315948 78328 316000 78334
rect 316000 78276 316080 78282
rect 315948 78270 316080 78276
rect 315960 78254 316080 78270
rect 472650 78266 473032 78282
rect 316052 77330 316080 78254
rect 324320 78260 324372 78266
rect 324320 78202 324372 78208
rect 471980 78260 472032 78266
rect 472650 78260 473044 78266
rect 472650 78254 472992 78260
rect 471980 78202 472032 78208
rect 472992 78202 473044 78208
rect 316052 77302 316158 77330
rect 313280 75880 313332 75886
rect 313280 75822 313332 75828
rect 313292 74534 313320 75822
rect 313292 74506 313688 74534
rect 305368 74044 305420 74050
rect 305368 73986 305420 73992
rect 303712 72752 303764 72758
rect 303712 72694 303764 72700
rect 302332 64864 302384 64870
rect 302332 64806 302384 64812
rect 302344 64394 302372 64806
rect 302332 64388 302384 64394
rect 302332 64330 302384 64336
rect 303724 54754 303752 72694
rect 303804 62076 303856 62082
rect 303804 62018 303856 62024
rect 303816 61441 303844 62018
rect 303802 61432 303858 61441
rect 303802 61367 303858 61376
rect 305380 54754 305408 73986
rect 307024 68604 307076 68610
rect 307024 68546 307076 68552
rect 307036 54754 307064 68546
rect 310520 67108 310572 67114
rect 310520 67050 310572 67056
rect 309048 57588 309100 57594
rect 309048 57530 309100 57536
rect 292132 54726 292514 54754
rect 293972 54726 294170 54754
rect 295444 54726 295826 54754
rect 297100 54726 297482 54754
rect 298756 54726 299138 54754
rect 300412 54726 300794 54754
rect 302252 54726 302450 54754
rect 303724 54726 304106 54754
rect 305380 54726 305762 54754
rect 307036 54726 307418 54754
rect 309060 54740 309088 57530
rect 310532 54754 310560 67050
rect 312360 56636 312412 56642
rect 312360 56578 312412 56584
rect 310532 54726 310730 54754
rect 312372 54740 312400 56578
rect 313660 54754 313688 74506
rect 315304 61600 315356 61606
rect 315304 61542 315356 61548
rect 315316 54754 315344 61542
rect 316052 56642 316080 77302
rect 321940 75886 321968 77316
rect 324332 75886 324360 78202
rect 328460 78192 328512 78198
rect 328460 78134 328512 78140
rect 333244 78192 333296 78198
rect 454040 78192 454092 78198
rect 333296 78140 333546 78146
rect 333244 78134 333546 78140
rect 455328 78192 455380 78198
rect 454040 78134 454092 78140
rect 455262 78140 455328 78146
rect 455262 78134 455380 78140
rect 327736 75886 327764 77316
rect 321928 75880 321980 75886
rect 321928 75822 321980 75828
rect 323584 75880 323636 75886
rect 323584 75822 323636 75828
rect 324320 75880 324372 75886
rect 324320 75822 324372 75828
rect 327724 75880 327776 75886
rect 327724 75822 327776 75828
rect 322940 72684 322992 72690
rect 322940 72626 322992 72632
rect 318800 60376 318852 60382
rect 318800 60318 318852 60324
rect 316960 58948 317012 58954
rect 316960 58890 317012 58896
rect 316040 56636 316092 56642
rect 316040 56578 316092 56584
rect 316972 54754 317000 58890
rect 318812 54754 318840 60318
rect 321928 60308 321980 60314
rect 321928 60250 321980 60256
rect 320088 60240 320140 60246
rect 320088 60182 320140 60188
rect 320100 57594 320128 60182
rect 321940 59265 321968 60250
rect 321926 59256 321982 59265
rect 321926 59191 321982 59200
rect 320824 58880 320876 58886
rect 320824 58822 320876 58828
rect 320836 57934 320864 58822
rect 320824 57928 320876 57934
rect 320824 57870 320876 57876
rect 320088 57588 320140 57594
rect 320088 57530 320140 57536
rect 320836 54754 320864 57870
rect 313660 54726 314042 54754
rect 315316 54726 315698 54754
rect 316972 54726 317354 54754
rect 318812 54726 319010 54754
rect 320666 54726 320864 54754
rect 321940 54754 321968 59191
rect 322952 55214 322980 72626
rect 323596 61606 323624 75822
rect 328472 75682 328500 78134
rect 333256 78118 333546 78134
rect 365720 78124 365772 78130
rect 365720 78066 365772 78072
rect 449808 78124 449860 78130
rect 449808 78066 449860 78072
rect 333244 76560 333296 76566
rect 333244 76502 333296 76508
rect 333256 75886 333284 76502
rect 339328 75886 339356 77316
rect 333244 75880 333296 75886
rect 333244 75822 333296 75828
rect 339316 75880 339368 75886
rect 339316 75822 339368 75828
rect 327724 75676 327776 75682
rect 327724 75618 327776 75624
rect 328460 75676 328512 75682
rect 328460 75618 328512 75624
rect 323584 61600 323636 61606
rect 323584 61542 323636 61548
rect 325240 61532 325292 61538
rect 325240 61474 325292 61480
rect 322952 55186 323624 55214
rect 323596 54754 323624 55186
rect 325252 54754 325280 61474
rect 327736 58954 327764 75618
rect 329748 74044 329800 74050
rect 329748 73986 329800 73992
rect 329760 73166 329788 73986
rect 328552 73160 328604 73166
rect 328552 73102 328604 73108
rect 329748 73160 329800 73166
rect 329748 73102 329800 73108
rect 327724 58948 327776 58954
rect 327724 58890 327776 58896
rect 328368 58744 328420 58750
rect 328368 58686 328420 58692
rect 328380 58585 328408 58686
rect 327078 58576 327134 58585
rect 327078 58511 327134 58520
rect 328366 58576 328422 58585
rect 328366 58511 328422 58520
rect 327092 54754 327120 58511
rect 328564 54754 328592 73102
rect 330208 69896 330260 69902
rect 330208 69838 330260 69844
rect 330220 54754 330248 69838
rect 333256 60382 333284 75822
rect 345124 74594 345152 77316
rect 350552 77302 350934 77330
rect 338764 74588 338816 74594
rect 338764 74530 338816 74536
rect 345112 74588 345164 74594
rect 345112 74530 345164 74536
rect 338488 73840 338540 73846
rect 338488 73782 338540 73788
rect 336648 67108 336700 67114
rect 336648 67050 336700 67056
rect 336660 66881 336688 67050
rect 335358 66872 335414 66881
rect 335358 66807 335414 66816
rect 336646 66872 336702 66881
rect 336646 66807 336702 66816
rect 333244 60376 333296 60382
rect 333244 60318 333296 60324
rect 331864 60240 331916 60246
rect 331864 60182 331916 60188
rect 331876 54754 331904 60182
rect 332968 60172 333020 60178
rect 332968 60114 333020 60120
rect 332980 59362 333008 60114
rect 332968 59356 333020 59362
rect 332968 59298 333020 59304
rect 333520 59356 333572 59362
rect 333520 59298 333572 59304
rect 333532 54754 333560 59298
rect 335372 54754 335400 66807
rect 336832 58812 336884 58818
rect 336832 58754 336884 58760
rect 336844 54754 336872 58754
rect 338500 54754 338528 73782
rect 338776 58886 338804 74530
rect 340144 72480 340196 72486
rect 340144 72422 340196 72428
rect 338764 58880 338816 58886
rect 338764 58822 338816 58828
rect 340156 54754 340184 72422
rect 341800 69692 341852 69698
rect 341800 69634 341852 69640
rect 341812 54754 341840 69634
rect 343640 68332 343692 68338
rect 343640 68274 343692 68280
rect 343652 54754 343680 68274
rect 345112 63028 345164 63034
rect 345112 62970 345164 62976
rect 345124 54754 345152 62970
rect 350080 62960 350132 62966
rect 350080 62902 350132 62908
rect 348424 62892 348476 62898
rect 348424 62834 348476 62840
rect 346768 62824 346820 62830
rect 346768 62766 346820 62772
rect 346780 54754 346808 62766
rect 348436 54754 348464 62834
rect 350092 54754 350120 62902
rect 350552 60314 350580 77302
rect 356716 72690 356744 77316
rect 362052 77302 362526 77330
rect 362052 74534 362080 77302
rect 361592 74506 362080 74534
rect 365732 74534 365760 78066
rect 385040 78056 385092 78062
rect 385040 77998 385092 78004
rect 420736 78056 420788 78062
rect 420736 77998 420788 78004
rect 367112 77302 368322 77330
rect 365732 74506 366680 74534
rect 356704 72684 356756 72690
rect 356704 72626 356756 72632
rect 355048 72548 355100 72554
rect 355048 72490 355100 72496
rect 353392 71052 353444 71058
rect 353392 70994 353444 71000
rect 351920 68400 351972 68406
rect 351920 68342 351972 68348
rect 350540 60308 350592 60314
rect 350540 60250 350592 60256
rect 351932 54754 351960 68342
rect 353404 54754 353432 70994
rect 355060 54754 355088 72490
rect 360200 71120 360252 71126
rect 360200 71062 360252 71068
rect 356704 69760 356756 69766
rect 356704 69702 356756 69708
rect 356716 54754 356744 69702
rect 358360 68468 358412 68474
rect 358360 68410 358412 68416
rect 358372 54754 358400 68410
rect 360212 54754 360240 71062
rect 361592 61538 361620 74506
rect 363328 73908 363380 73914
rect 363328 73850 363380 73856
rect 361672 66972 361724 66978
rect 361672 66914 361724 66920
rect 361580 61532 361632 61538
rect 361580 61474 361632 61480
rect 361684 54754 361712 66914
rect 363340 54754 363368 73850
rect 365352 57588 365404 57594
rect 365352 57530 365404 57536
rect 321940 54726 322322 54754
rect 323596 54726 323978 54754
rect 325252 54726 325634 54754
rect 327092 54726 327290 54754
rect 328564 54726 328946 54754
rect 330220 54726 330602 54754
rect 331876 54726 332258 54754
rect 333532 54726 333914 54754
rect 335372 54726 335570 54754
rect 336844 54726 337226 54754
rect 338500 54726 338882 54754
rect 340156 54726 340538 54754
rect 341812 54726 342194 54754
rect 343652 54726 343850 54754
rect 345124 54726 345506 54754
rect 346780 54726 347162 54754
rect 348436 54726 348818 54754
rect 350092 54726 350474 54754
rect 351932 54726 352130 54754
rect 353404 54726 353786 54754
rect 355060 54726 355442 54754
rect 356716 54726 357098 54754
rect 358372 54726 358754 54754
rect 360212 54726 360410 54754
rect 361684 54726 362066 54754
rect 363340 54726 363722 54754
rect 365364 54740 365392 57530
rect 366652 54754 366680 74506
rect 367112 58750 367140 77302
rect 372620 76560 372672 76566
rect 372620 76502 372672 76508
rect 372632 74534 372660 76502
rect 372632 74506 373304 74534
rect 371608 60104 371660 60110
rect 371608 60046 371660 60052
rect 367100 58744 367152 58750
rect 367100 58686 367152 58692
rect 368664 57520 368716 57526
rect 368664 57462 368716 57468
rect 366652 54726 367034 54754
rect 368676 54740 368704 57462
rect 370320 57452 370372 57458
rect 370320 57394 370372 57400
rect 370332 54740 370360 57394
rect 371620 54754 371648 60046
rect 373276 54754 373304 74506
rect 374104 74050 374132 77316
rect 376760 76628 376812 76634
rect 376760 76570 376812 76576
rect 374182 76528 374238 76537
rect 374182 76463 374238 76472
rect 374196 74534 374224 76463
rect 374196 74506 374960 74534
rect 374092 74044 374144 74050
rect 374092 73986 374144 73992
rect 374932 54754 374960 74506
rect 376772 54754 376800 76570
rect 378232 73840 378284 73846
rect 378232 73782 378284 73788
rect 378244 54754 378272 73782
rect 379900 69902 379928 77316
rect 382280 76696 382332 76702
rect 382280 76638 382332 76644
rect 382292 74534 382320 76638
rect 382292 74506 383240 74534
rect 379888 69896 379940 69902
rect 379888 69838 379940 69844
rect 379888 62824 379940 62830
rect 379888 62766 379940 62772
rect 379900 54754 379928 62766
rect 381544 61464 381596 61470
rect 381544 61406 381596 61412
rect 381556 54754 381584 61406
rect 383212 54754 383240 74506
rect 385052 54754 385080 77998
rect 420748 77330 420776 77998
rect 449820 77330 449848 78066
rect 385236 77302 385710 77330
rect 390664 77302 391506 77330
rect 396092 77302 397302 77330
rect 402992 77302 403098 77330
rect 385236 64874 385264 77302
rect 390560 76832 390612 76838
rect 390560 76774 390612 76780
rect 389178 76664 389234 76673
rect 389178 76599 389234 76608
rect 389192 74534 389220 76599
rect 389192 74506 389864 74534
rect 385144 64846 385264 64874
rect 385144 60246 385172 64846
rect 385132 60240 385184 60246
rect 385132 60182 385184 60188
rect 386878 57352 386934 57361
rect 386878 57287 386934 57296
rect 371620 54726 372002 54754
rect 373276 54726 373658 54754
rect 374932 54726 375314 54754
rect 376772 54726 376970 54754
rect 378244 54726 378626 54754
rect 379900 54726 380282 54754
rect 381556 54726 381938 54754
rect 383212 54726 383594 54754
rect 385052 54726 385250 54754
rect 386892 54740 386920 57287
rect 388534 57216 388590 57225
rect 388534 57151 388590 57160
rect 388548 54740 388576 57151
rect 389836 54754 389864 74506
rect 390572 55214 390600 76774
rect 390664 60178 390692 77302
rect 393320 76764 393372 76770
rect 393320 76706 393372 76712
rect 390652 60172 390704 60178
rect 390652 60114 390704 60120
rect 390572 55186 391520 55214
rect 391492 54754 391520 55186
rect 393332 54754 393360 76706
rect 394700 76696 394752 76702
rect 394700 76638 394752 76644
rect 394712 74534 394740 76638
rect 394712 74506 394832 74534
rect 394804 54754 394832 74506
rect 396092 67114 396120 77302
rect 398840 76900 398892 76906
rect 398840 76842 398892 76848
rect 396080 67108 396132 67114
rect 396080 67050 396132 67056
rect 396448 58744 396500 58750
rect 396448 58686 396500 58692
rect 396460 54754 396488 58686
rect 389836 54726 390218 54754
rect 391492 54726 391874 54754
rect 393332 54726 393530 54754
rect 394804 54726 395186 54754
rect 396460 54726 396842 54754
rect 356992 24274 357374 24290
rect 356980 24268 357374 24274
rect 357032 24262 357374 24268
rect 356980 24210 357032 24216
rect 398852 24206 398880 76842
rect 402992 58818 403020 77302
rect 408880 75886 408908 77316
rect 414676 75886 414704 77316
rect 420288 77314 420776 77330
rect 419540 77308 419592 77314
rect 419540 77250 419592 77256
rect 420276 77308 420776 77314
rect 420328 77302 420776 77308
rect 425072 77302 426282 77330
rect 431972 77302 432078 77330
rect 437874 77302 438164 77330
rect 420276 77250 420328 77256
rect 408868 75880 408920 75886
rect 408868 75822 408920 75828
rect 414664 75880 414716 75886
rect 414664 75822 414716 75828
rect 408880 71262 408908 75822
rect 408868 71256 408920 71262
rect 408868 71198 408920 71204
rect 419552 60042 419580 77250
rect 425072 62082 425100 77302
rect 431972 64870 432000 77302
rect 438136 71738 438164 77302
rect 438124 71732 438176 71738
rect 438124 71674 438176 71680
rect 431960 64864 432012 64870
rect 431960 64806 432012 64812
rect 425060 62076 425112 62082
rect 425060 62018 425112 62024
rect 438136 61402 438164 71674
rect 443656 71670 443684 77316
rect 449268 77314 449848 77330
rect 448520 77308 448572 77314
rect 448520 77250 448572 77256
rect 449256 77308 449848 77314
rect 449308 77302 449848 77308
rect 449256 77250 449308 77256
rect 443644 71664 443696 71670
rect 443644 71606 443696 71612
rect 443656 64258 443684 71606
rect 443644 64252 443696 64258
rect 443644 64194 443696 64200
rect 438124 61396 438176 61402
rect 438124 61338 438176 61344
rect 419540 60036 419592 60042
rect 419540 59978 419592 59984
rect 402980 58812 403032 58818
rect 402980 58754 403032 58760
rect 448532 58682 448560 77250
rect 454052 65686 454080 78134
rect 455262 78118 455368 78134
rect 461044 73166 461072 77316
rect 466854 77302 467144 77330
rect 467116 75886 467144 77302
rect 467104 75880 467156 75886
rect 467104 75822 467156 75828
rect 461032 73160 461084 73166
rect 461032 73102 461084 73108
rect 461044 72350 461072 73102
rect 461032 72344 461084 72350
rect 461032 72286 461084 72292
rect 461584 72344 461636 72350
rect 461584 72286 461636 72292
rect 454040 65680 454092 65686
rect 454040 65622 454092 65628
rect 461596 64190 461624 72286
rect 467116 65618 467144 75822
rect 471992 66910 472020 78202
rect 477512 77302 478446 77330
rect 483676 77302 484242 77330
rect 471980 66904 472032 66910
rect 471980 66846 472032 66852
rect 467104 65612 467156 65618
rect 467104 65554 467156 65560
rect 477512 64326 477540 77302
rect 483676 75818 483704 77302
rect 483664 75812 483716 75818
rect 483664 75754 483716 75760
rect 477500 64320 477552 64326
rect 477500 64262 477552 64268
rect 461584 64184 461636 64190
rect 461584 64126 461636 64132
rect 448520 58676 448572 58682
rect 448520 58618 448572 58624
rect 483676 57390 483704 75754
rect 490024 75342 490052 77316
rect 495834 77302 496124 77330
rect 491208 75744 491260 75750
rect 491208 75686 491260 75692
rect 491220 75342 491248 75686
rect 496096 75682 496124 77302
rect 496084 75676 496136 75682
rect 496084 75618 496136 75624
rect 490012 75336 490064 75342
rect 490012 75278 490064 75284
rect 491208 75336 491260 75342
rect 491208 75278 491260 75284
rect 483664 57384 483716 57390
rect 483664 57326 483716 57332
rect 496096 57322 496124 75618
rect 501616 75614 501644 77316
rect 507136 77302 507426 77330
rect 501604 75608 501656 75614
rect 501604 75550 501656 75556
rect 501616 75274 501644 75550
rect 501604 75268 501656 75274
rect 501604 75210 501656 75216
rect 507136 74497 507164 77302
rect 513208 75546 513236 77316
rect 519004 75857 519032 77316
rect 518990 75848 519046 75857
rect 518990 75783 519046 75792
rect 513196 75540 513248 75546
rect 513196 75482 513248 75488
rect 513208 75206 513236 75482
rect 513196 75200 513248 75206
rect 513196 75142 513248 75148
rect 507122 74488 507178 74497
rect 507122 74423 507178 74432
rect 496084 57316 496136 57322
rect 496084 57258 496136 57264
rect 507136 57254 507164 74423
rect 519004 69834 519032 75783
rect 524800 74526 524828 77316
rect 524788 74520 524840 74526
rect 524788 74462 524840 74468
rect 524800 72622 524828 74462
rect 530596 74458 530624 77316
rect 536116 77302 536406 77330
rect 530584 74452 530636 74458
rect 530584 74394 530636 74400
rect 530596 73982 530624 74394
rect 536116 74390 536144 77302
rect 536104 74384 536156 74390
rect 536104 74326 536156 74332
rect 530584 73976 530636 73982
rect 530584 73918 530636 73924
rect 524788 72616 524840 72622
rect 524788 72558 524840 72564
rect 518992 69828 519044 69834
rect 518992 69770 519044 69776
rect 536116 67046 536144 74326
rect 542188 74322 542216 77316
rect 547892 77302 547998 77330
rect 553412 77302 553794 77330
rect 542176 74316 542228 74322
rect 542176 74258 542228 74264
rect 542188 68542 542216 74258
rect 547892 74254 547920 77302
rect 547880 74248 547932 74254
rect 547880 74190 547932 74196
rect 547892 71194 547920 74190
rect 547880 71188 547932 71194
rect 547880 71130 547932 71136
rect 542176 68536 542228 68542
rect 542176 68478 542228 68484
rect 536104 67040 536156 67046
rect 536104 66982 536156 66988
rect 553412 62830 553440 77302
rect 559576 74186 559604 77316
rect 565004 77302 565386 77330
rect 559564 74180 559616 74186
rect 559564 74122 559616 74128
rect 559576 65550 559604 74122
rect 559564 65544 559616 65550
rect 559564 65486 559616 65492
rect 565004 64874 565032 77302
rect 568684 74390 568712 204070
rect 568776 75546 568804 204342
rect 568868 188698 568896 314638
rect 568856 188692 568908 188698
rect 568856 188634 568908 188640
rect 568868 187746 568896 188634
rect 568856 187740 568908 187746
rect 568856 187682 568908 187688
rect 568960 76838 568988 458186
rect 568948 76832 569000 76838
rect 568948 76774 569000 76780
rect 568764 75540 568816 75546
rect 568764 75482 568816 75488
rect 568672 74384 568724 74390
rect 568672 74326 568724 74332
rect 564452 64846 565032 64874
rect 553400 62824 553452 62830
rect 553400 62766 553452 62772
rect 564452 58750 564480 64846
rect 564440 58744 564492 58750
rect 564440 58686 564492 58692
rect 507124 57248 507176 57254
rect 507124 57190 507176 57196
rect 400218 54496 400274 54505
rect 400218 54431 400274 54440
rect 364432 24200 364484 24206
rect 382832 24200 382884 24206
rect 364484 24148 364550 24154
rect 364432 24142 364550 24148
rect 364444 24126 364550 24142
rect 375024 24138 375314 24154
rect 375012 24132 375314 24138
rect 375064 24126 375314 24132
rect 382490 24148 382832 24154
rect 398840 24200 398892 24206
rect 382490 24142 382884 24148
rect 382490 24126 382872 24142
rect 393254 24138 393360 24154
rect 398840 24142 398892 24148
rect 393254 24132 393372 24138
rect 393254 24126 393320 24132
rect 375012 24074 375064 24080
rect 393320 24074 393372 24080
rect 266360 23520 266412 23526
rect 266360 23462 266412 23468
rect 267372 23520 267424 23526
rect 267424 23468 267674 23474
rect 267372 23462 267674 23468
rect 202892 23310 203090 23338
rect 205652 23310 206678 23338
rect 209792 23310 210266 23338
rect 212552 23310 213854 23338
rect 216692 23310 217442 23338
rect 220832 23310 221030 23338
rect 223592 23310 224618 23338
rect 199384 22092 199436 22098
rect 199384 22034 199436 22040
rect 175464 21548 175516 21554
rect 175464 21490 175516 21496
rect 152464 21412 152516 21418
rect 152464 21354 152516 21360
rect 138020 19984 138072 19990
rect 138020 19926 138072 19932
rect 131120 17332 131172 17338
rect 131120 17274 131172 17280
rect 131132 16574 131160 17274
rect 138032 16574 138060 19926
rect 150440 18692 150492 18698
rect 150440 18634 150492 18640
rect 142160 18624 142212 18630
rect 142160 18566 142212 18572
rect 131132 16546 131344 16574
rect 138032 16546 138888 16574
rect 125600 11892 125652 11898
rect 125600 11834 125652 11840
rect 96620 4820 96672 4826
rect 96620 4762 96672 4768
rect 66260 3460 66312 3466
rect 66260 3402 66312 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 11834
rect 128176 7676 128228 7682
rect 128176 7618 128228 7624
rect 128188 480 128216 7618
rect 129372 4956 129424 4962
rect 129372 4898 129424 4904
rect 129384 480 129412 4898
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 135260 15972 135312 15978
rect 135260 15914 135312 15920
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 132972 480 133000 3470
rect 135272 480 135300 15914
rect 136456 14612 136508 14618
rect 136456 14554 136508 14560
rect 136468 480 136496 14554
rect 138860 480 138888 16546
rect 139584 13252 139636 13258
rect 139584 13194 139636 13200
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 13194
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 18566
rect 150452 16574 150480 18634
rect 150452 16546 150664 16574
rect 147128 10396 147180 10402
rect 147128 10338 147180 10344
rect 143540 6384 143592 6390
rect 143540 6326 143592 6332
rect 143552 480 143580 6326
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 145944 480 145972 3538
rect 147140 480 147168 10338
rect 149520 3868 149572 3874
rect 149520 3810 149572 3816
rect 149532 480 149560 3810
rect 150636 480 150664 16546
rect 151820 11756 151872 11762
rect 151820 11698 151872 11704
rect 151832 3398 151860 11698
rect 152476 3874 152504 21354
rect 162860 20052 162912 20058
rect 162860 19994 162912 20000
rect 155960 18828 156012 18834
rect 155960 18770 156012 18776
rect 155972 16574 156000 18770
rect 162872 16574 162900 19994
rect 175280 18760 175332 18766
rect 175280 18702 175332 18708
rect 171140 17400 171192 17406
rect 171140 17342 171192 17348
rect 171152 16574 171180 17342
rect 175292 16574 175320 18702
rect 175476 18630 175504 21490
rect 187700 21480 187752 21486
rect 187700 21422 187752 21428
rect 178040 20120 178092 20126
rect 178040 20062 178092 20068
rect 175464 18624 175516 18630
rect 175464 18566 175516 18572
rect 178052 16574 178080 20062
rect 187712 18834 187740 21422
rect 187700 18828 187752 18834
rect 187700 18770 187752 18776
rect 184940 18624 184992 18630
rect 184940 18566 184992 18572
rect 155972 16546 156184 16574
rect 162872 16546 163728 16574
rect 171152 16546 172008 16574
rect 175292 16546 175504 16574
rect 178052 16546 178632 16574
rect 153752 11960 153804 11966
rect 153752 11902 153804 11908
rect 152464 3868 152516 3874
rect 152464 3810 152516 3816
rect 151820 3392 151872 3398
rect 151820 3334 151872 3340
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 11902
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 160100 13184 160152 13190
rect 160100 13126 160152 13132
rect 156604 10464 156656 10470
rect 156604 10406 156656 10412
rect 156616 3534 156644 10406
rect 157800 7744 157852 7750
rect 157800 7686 157852 7692
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157812 480 157840 7686
rect 160112 3534 160140 13126
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 160100 2848 160152 2854
rect 160100 2790 160152 2796
rect 160112 480 160140 2790
rect 161308 480 161336 3470
rect 161400 2854 161428 3470
rect 161388 2848 161440 2854
rect 161388 2790 161440 2796
rect 163700 480 163728 16546
rect 168380 16040 168432 16046
rect 168380 15982 168432 15988
rect 164424 14544 164476 14550
rect 164424 14486 164476 14492
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14486
rect 167184 9036 167236 9042
rect 167184 8978 167236 8984
rect 167196 480 167224 8978
rect 168392 480 168420 15982
rect 170312 14476 170364 14482
rect 170312 14418 170364 14424
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 14418
rect 171980 480 172008 16546
rect 174268 9104 174320 9110
rect 174268 9046 174320 9052
rect 174280 480 174308 9046
rect 175476 480 175504 16546
rect 176660 13116 176712 13122
rect 176660 13058 176712 13064
rect 176672 3398 176700 13058
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 177856 3392 177908 3398
rect 177856 3334 177908 3340
rect 177868 480 177896 3334
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 181444 6316 181496 6322
rect 181444 6258 181496 6264
rect 181456 480 181484 6258
rect 182548 5024 182600 5030
rect 182548 4966 182600 4972
rect 182560 480 182588 4966
rect 184952 480 184980 18566
rect 202892 11898 202920 23310
rect 202880 11892 202932 11898
rect 202880 11834 202932 11840
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 186148 480 186176 11766
rect 205652 4962 205680 23310
rect 209792 10470 209820 23310
rect 212552 14618 212580 23310
rect 212540 14612 212592 14618
rect 212540 14554 212592 14560
rect 216692 13258 216720 23310
rect 216680 13252 216732 13258
rect 216680 13194 216732 13200
rect 209780 10464 209832 10470
rect 209780 10406 209832 10412
rect 220832 6390 220860 23310
rect 223592 10402 223620 23310
rect 228192 18698 228220 23324
rect 230492 23310 231794 23338
rect 234632 23310 235382 23338
rect 238772 23310 238970 23338
rect 241532 23310 242558 23338
rect 245672 23310 246146 23338
rect 228180 18692 228232 18698
rect 228180 18634 228232 18640
rect 230492 11966 230520 23310
rect 230480 11960 230532 11966
rect 230480 11902 230532 11908
rect 223580 10396 223632 10402
rect 223580 10338 223632 10344
rect 234632 7750 234660 23310
rect 238772 13190 238800 23310
rect 241532 14550 241560 23310
rect 242900 17264 242952 17270
rect 242900 17206 242952 17212
rect 241520 14544 241572 14550
rect 241520 14486 241572 14492
rect 238760 13184 238812 13190
rect 238760 13126 238812 13132
rect 241704 8968 241756 8974
rect 241704 8910 241756 8916
rect 234620 7744 234672 7750
rect 234620 7686 234672 7692
rect 235908 7744 235960 7750
rect 235908 7686 235960 7692
rect 220820 6384 220872 6390
rect 220820 6326 220872 6332
rect 205640 4956 205692 4962
rect 205640 4898 205692 4904
rect 188528 4888 188580 4894
rect 188528 4830 188580 4836
rect 188540 480 188568 4830
rect 235920 3602 235948 7686
rect 235908 3596 235960 3602
rect 235908 3538 235960 3544
rect 239312 3460 239364 3466
rect 239312 3402 239364 3408
rect 239324 480 239352 3402
rect 241716 480 241744 8910
rect 242912 480 242940 17206
rect 245672 16046 245700 23310
rect 249720 17406 249748 23324
rect 253308 18766 253336 23324
rect 256896 20126 256924 23324
rect 259472 23310 260498 23338
rect 263612 23310 264086 23338
rect 256884 20120 256936 20126
rect 256884 20062 256936 20068
rect 253296 18760 253348 18766
rect 253296 18702 253348 18708
rect 249708 17400 249760 17406
rect 249708 17342 249760 17348
rect 245660 16040 245712 16046
rect 245660 15982 245712 15988
rect 245936 15904 245988 15910
rect 245936 15846 245988 15852
rect 245200 7608 245252 7614
rect 245200 7550 245252 7556
rect 245212 480 245240 7550
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 15846
rect 248788 6248 248840 6254
rect 248788 6190 248840 6196
rect 248800 480 248828 6190
rect 249984 6180 250036 6186
rect 249984 6122 250036 6128
rect 249996 480 250024 6122
rect 259472 5030 259500 23310
rect 263612 11830 263640 23310
rect 263600 11824 263652 11830
rect 263600 11766 263652 11772
rect 259460 5024 259512 5030
rect 259460 4966 259512 4972
rect 252376 4820 252428 4826
rect 252376 4762 252428 4768
rect 252388 480 252416 4762
rect 266372 3466 266400 23462
rect 267384 23446 267674 23462
rect 270512 23310 271262 23338
rect 270512 7682 270540 23310
rect 274836 17338 274864 23324
rect 277412 23310 278438 23338
rect 274824 17332 274876 17338
rect 274824 17274 274876 17280
rect 277412 15978 277440 23310
rect 282012 19990 282040 23324
rect 285600 21554 285628 23324
rect 288452 23310 289202 23338
rect 285588 21548 285640 21554
rect 285588 21490 285640 21496
rect 282000 19984 282052 19990
rect 282000 19926 282052 19932
rect 277400 15972 277452 15978
rect 277400 15914 277452 15920
rect 288452 7750 288480 23310
rect 292776 21418 292804 23324
rect 295352 23310 296378 23338
rect 292764 21412 292816 21418
rect 292764 21354 292816 21360
rect 295352 11762 295380 23310
rect 299952 21486 299980 23324
rect 302252 23310 303554 23338
rect 299940 21480 299992 21486
rect 299940 21422 299992 21428
rect 295340 11756 295392 11762
rect 295340 11698 295392 11704
rect 288440 7744 288492 7750
rect 288440 7686 288492 7692
rect 270500 7676 270552 7682
rect 270500 7618 270552 7624
rect 302252 3534 302280 23310
rect 307128 20058 307156 23324
rect 310532 23310 310730 23338
rect 313292 23310 314318 23338
rect 317432 23310 317906 23338
rect 320192 23310 321494 23338
rect 324332 23310 325082 23338
rect 307116 20052 307168 20058
rect 307116 19994 307168 20000
rect 310532 9042 310560 23310
rect 313292 14482 313320 23310
rect 313280 14476 313332 14482
rect 313280 14418 313332 14424
rect 317432 9110 317460 23310
rect 320192 13122 320220 23310
rect 320180 13116 320232 13122
rect 320180 13058 320232 13064
rect 317420 9104 317472 9110
rect 317420 9046 317472 9052
rect 310520 9036 310572 9042
rect 310520 8978 310572 8984
rect 324332 6322 324360 23310
rect 328656 18630 328684 23324
rect 331232 23310 332258 23338
rect 328644 18624 328696 18630
rect 328644 18566 328696 18572
rect 324320 6316 324372 6322
rect 324320 6258 324372 6264
rect 331232 4894 331260 23310
rect 335832 22234 335860 23324
rect 338132 23310 339434 23338
rect 335820 22228 335872 22234
rect 335820 22170 335872 22176
rect 338132 10334 338160 23310
rect 343008 21865 343036 23324
rect 346596 22166 346624 23324
rect 346584 22160 346636 22166
rect 346584 22102 346636 22108
rect 350184 22098 350212 23324
rect 353772 22302 353800 23324
rect 353760 22296 353812 22302
rect 353760 22238 353812 22244
rect 350172 22092 350224 22098
rect 350172 22034 350224 22040
rect 360948 21962 360976 23324
rect 368124 22001 368152 23324
rect 371712 22030 371740 23324
rect 371700 22024 371752 22030
rect 368110 21992 368166 22001
rect 360936 21956 360988 21962
rect 371700 21966 371752 21972
rect 378888 21962 378916 23324
rect 386064 22098 386092 23324
rect 389652 22137 389680 23324
rect 389638 22128 389694 22137
rect 386052 22092 386104 22098
rect 389638 22063 389694 22072
rect 386052 22034 386104 22040
rect 396828 22030 396856 23324
rect 396816 22024 396868 22030
rect 396816 21966 396868 21972
rect 400232 21962 400260 54431
rect 569236 24138 569264 485046
rect 569328 459610 569356 585822
rect 569316 459604 569368 459610
rect 569316 459546 569368 459552
rect 569328 459406 569356 459546
rect 569972 459474 570000 586162
rect 572720 586152 572772 586158
rect 572720 586094 572772 586100
rect 570144 586084 570196 586090
rect 570144 586026 570196 586032
rect 570052 586016 570104 586022
rect 570052 585958 570104 585964
rect 569960 459468 570012 459474
rect 569960 459410 570012 459416
rect 569316 459400 569368 459406
rect 569316 459342 569368 459348
rect 569316 458856 569368 458862
rect 569316 458798 569368 458804
rect 569328 315858 569356 458798
rect 569972 458590 570000 459410
rect 569960 458584 570012 458590
rect 569960 458526 570012 458532
rect 569960 458448 570012 458454
rect 569960 458390 570012 458396
rect 569972 332314 570000 458390
rect 570064 458046 570092 585958
rect 570156 459270 570184 586026
rect 571524 583364 571576 583370
rect 571524 583306 571576 583312
rect 571432 583296 571484 583302
rect 571432 583238 571484 583244
rect 571340 583024 571392 583030
rect 571340 582966 571392 582972
rect 570236 572212 570288 572218
rect 570236 572154 570288 572160
rect 570248 459338 570276 572154
rect 570328 462324 570380 462330
rect 570328 462266 570380 462272
rect 570340 461106 570368 462266
rect 571352 461378 571380 582966
rect 571340 461372 571392 461378
rect 571340 461314 571392 461320
rect 571444 461174 571472 583238
rect 571536 461310 571564 583306
rect 571616 583160 571668 583166
rect 571616 583102 571668 583108
rect 571628 462330 571656 583102
rect 571708 572144 571760 572150
rect 571708 572086 571760 572092
rect 571616 462324 571668 462330
rect 571616 462266 571668 462272
rect 571524 461304 571576 461310
rect 571524 461246 571576 461252
rect 571432 461168 571484 461174
rect 571432 461110 571484 461116
rect 570328 461100 570380 461106
rect 570328 461042 570380 461048
rect 570236 459332 570288 459338
rect 570236 459274 570288 459280
rect 570144 459264 570196 459270
rect 570144 459206 570196 459212
rect 570156 458454 570184 459206
rect 570144 458448 570196 458454
rect 570144 458390 570196 458396
rect 570248 458250 570276 459274
rect 570236 458244 570288 458250
rect 570236 458186 570288 458192
rect 570052 458040 570104 458046
rect 570052 457982 570104 457988
rect 570064 451274 570092 457982
rect 570064 451246 570184 451274
rect 570156 335354 570184 451246
rect 570236 443692 570288 443698
rect 570236 443634 570288 443640
rect 570248 336705 570276 443634
rect 570234 336696 570290 336705
rect 570234 336631 570290 336640
rect 570064 335326 570184 335354
rect 570064 332382 570092 335326
rect 570340 333266 570368 461042
rect 571536 460934 571564 461246
rect 571352 460906 571564 460934
rect 570420 458584 570472 458590
rect 570420 458526 570472 458532
rect 570432 458182 570460 458526
rect 570420 458176 570472 458182
rect 570420 458118 570472 458124
rect 570604 378820 570656 378826
rect 570604 378762 570656 378768
rect 570328 333260 570380 333266
rect 570328 333202 570380 333208
rect 570052 332376 570104 332382
rect 570052 332318 570104 332324
rect 569960 332308 570012 332314
rect 569960 332250 570012 332256
rect 569316 315852 569368 315858
rect 569316 315794 569368 315800
rect 569328 314702 569356 315794
rect 569316 314696 569368 314702
rect 569316 314638 569368 314644
rect 569972 204066 570000 332250
rect 570064 204270 570092 332318
rect 570052 204264 570104 204270
rect 570052 204206 570104 204212
rect 569960 204060 570012 204066
rect 569960 204002 570012 204008
rect 569972 74254 570000 204002
rect 570064 74322 570092 204206
rect 570144 187740 570196 187746
rect 570144 187682 570196 187688
rect 570156 75818 570184 187682
rect 570144 75812 570196 75818
rect 570144 75754 570196 75760
rect 570052 74316 570104 74322
rect 570052 74258 570104 74264
rect 569960 74248 570012 74254
rect 569960 74190 570012 74196
rect 569224 24132 569276 24138
rect 569224 24074 569276 24080
rect 570616 22030 570644 378762
rect 571352 332926 571380 460906
rect 571616 459604 571668 459610
rect 571616 459546 571668 459552
rect 571430 458552 571486 458561
rect 571430 458487 571486 458496
rect 571340 332920 571392 332926
rect 571340 332862 571392 332868
rect 571352 332722 571380 332862
rect 571340 332716 571392 332722
rect 571340 332658 571392 332664
rect 571340 331900 571392 331906
rect 571340 331842 571392 331848
rect 571248 313336 571300 313342
rect 571248 313278 571300 313284
rect 571260 204950 571288 313278
rect 571248 204944 571300 204950
rect 571248 204886 571300 204892
rect 571352 76770 571380 331842
rect 571444 315314 571472 458487
rect 571524 458244 571576 458250
rect 571524 458186 571576 458192
rect 571536 325694 571564 458186
rect 571628 332586 571656 459546
rect 571720 458862 571748 572086
rect 571708 458856 571760 458862
rect 571708 458798 571760 458804
rect 571708 458176 571760 458182
rect 571708 458118 571760 458124
rect 571720 345014 571748 458118
rect 571720 344986 571932 345014
rect 571616 332580 571668 332586
rect 571616 332522 571668 332528
rect 571628 331294 571656 332522
rect 571904 332246 571932 344986
rect 571892 332240 571944 332246
rect 571892 332182 571944 332188
rect 571616 331288 571668 331294
rect 571616 331230 571668 331236
rect 571536 325666 571840 325694
rect 571812 315654 571840 325666
rect 571800 315648 571852 315654
rect 571800 315590 571852 315596
rect 571432 315308 571484 315314
rect 571432 315250 571484 315256
rect 571444 313342 571472 315250
rect 571524 314696 571576 314702
rect 571524 314638 571576 314644
rect 571432 313336 571484 313342
rect 571432 313278 571484 313284
rect 571432 204808 571484 204814
rect 571432 204750 571484 204756
rect 571444 204542 571472 204750
rect 571432 204536 571484 204542
rect 571432 204478 571484 204484
rect 571340 76764 571392 76770
rect 571340 76706 571392 76712
rect 571444 74458 571472 204478
rect 571536 204474 571564 314638
rect 571708 314628 571760 314634
rect 571708 314570 571760 314576
rect 571720 206378 571748 314570
rect 571708 206372 571760 206378
rect 571708 206314 571760 206320
rect 571812 204814 571840 315590
rect 571800 204808 571852 204814
rect 571800 204750 571852 204756
rect 571904 204626 571932 332182
rect 571628 204598 571932 204626
rect 571524 204468 571576 204474
rect 571524 204410 571576 204416
rect 571536 75682 571564 204410
rect 571628 203998 571656 204598
rect 571616 203992 571668 203998
rect 571616 203934 571668 203940
rect 571524 75676 571576 75682
rect 571524 75618 571576 75624
rect 571432 74452 571484 74458
rect 571432 74394 571484 74400
rect 571628 74186 571656 203934
rect 571708 203584 571760 203590
rect 571708 203526 571760 203532
rect 571616 74180 571668 74186
rect 571616 74122 571668 74128
rect 571720 73846 571748 203526
rect 572732 76566 572760 586094
rect 572812 583092 572864 583098
rect 572812 583034 572864 583040
rect 572824 444378 572852 583034
rect 572904 580304 572956 580310
rect 572904 580246 572956 580252
rect 572916 460970 572944 580246
rect 572996 572076 573048 572082
rect 572996 572018 573048 572024
rect 572904 460964 572956 460970
rect 572904 460906 572956 460912
rect 572812 444372 572864 444378
rect 572812 444314 572864 444320
rect 572824 332790 572852 444314
rect 572812 332784 572864 332790
rect 572812 332726 572864 332732
rect 572810 331800 572866 331809
rect 572810 331735 572866 331744
rect 572824 76634 572852 331735
rect 572916 315994 572944 460906
rect 573008 460902 573036 572018
rect 572996 460896 573048 460902
rect 572996 460838 573048 460844
rect 573008 459610 573036 460838
rect 572996 459604 573048 459610
rect 572996 459546 573048 459552
rect 572996 332716 573048 332722
rect 572996 332658 573048 332664
rect 572904 315988 572956 315994
rect 572904 315930 572956 315936
rect 572916 314770 572944 315930
rect 572904 314764 572956 314770
rect 572904 314706 572956 314712
rect 573008 204406 573036 332658
rect 573088 331288 573140 331294
rect 573088 331230 573140 331236
rect 572996 204400 573048 204406
rect 572996 204342 573048 204348
rect 573100 204218 573128 331230
rect 572916 204202 573128 204218
rect 572904 204196 573128 204202
rect 572956 204190 573128 204196
rect 572904 204138 572956 204144
rect 572812 76628 572864 76634
rect 572812 76570 572864 76576
rect 572720 76560 572772 76566
rect 572720 76502 572772 76508
rect 572916 74526 572944 204138
rect 572996 203652 573048 203658
rect 572996 203594 573048 203600
rect 573008 76702 573036 203594
rect 572996 76696 573048 76702
rect 572996 76638 573048 76644
rect 572904 74520 572956 74526
rect 572904 74462 572956 74468
rect 571708 73840 571760 73846
rect 571708 73782 571760 73788
rect 574112 22098 574140 696934
rect 580446 683904 580502 683913
rect 580446 683839 580502 683848
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 574192 583228 574244 583234
rect 574192 583170 574244 583176
rect 574204 461038 574232 583170
rect 575572 572008 575624 572014
rect 575572 571950 575624 571956
rect 575480 462460 575532 462466
rect 575480 462402 575532 462408
rect 574652 461168 574704 461174
rect 574652 461110 574704 461116
rect 574192 461032 574244 461038
rect 574192 460974 574244 460980
rect 574204 460934 574232 460974
rect 574204 460906 574508 460934
rect 574284 459604 574336 459610
rect 574284 459546 574336 459552
rect 574296 329798 574324 459546
rect 574480 329798 574508 460906
rect 574560 332784 574612 332790
rect 574560 332726 574612 332732
rect 574284 329792 574336 329798
rect 574284 329734 574336 329740
rect 574468 329792 574520 329798
rect 574468 329734 574520 329740
rect 574296 325694 574324 329734
rect 574296 325666 574416 325694
rect 574192 314696 574244 314702
rect 574192 314638 574244 314644
rect 574204 201482 574232 314638
rect 574192 201476 574244 201482
rect 574192 201418 574244 201424
rect 574284 201408 574336 201414
rect 574284 201350 574336 201356
rect 574296 200802 574324 201350
rect 574284 200796 574336 200802
rect 574284 200738 574336 200744
rect 574296 190454 574324 200738
rect 574204 190426 574324 190454
rect 574204 75750 574232 190426
rect 574388 188902 574416 325666
rect 574468 201476 574520 201482
rect 574468 201418 574520 201424
rect 574376 188896 574428 188902
rect 574376 188838 574428 188844
rect 574284 187944 574336 187950
rect 574284 187886 574336 187892
rect 574296 78266 574324 187886
rect 574388 187746 574416 188838
rect 574376 187740 574428 187746
rect 574376 187682 574428 187688
rect 574284 78260 574336 78266
rect 574284 78202 574336 78208
rect 574192 75744 574244 75750
rect 574192 75686 574244 75692
rect 574480 75614 574508 201418
rect 574572 188766 574600 332726
rect 574664 315790 574692 461110
rect 575492 317422 575520 462402
rect 575584 462398 575612 571950
rect 580262 524512 580318 524521
rect 580262 524447 580318 524456
rect 575572 462392 575624 462398
rect 575572 462334 575624 462340
rect 575584 331226 575612 462334
rect 575572 331220 575624 331226
rect 575572 331162 575624 331168
rect 576216 331220 576268 331226
rect 576216 331162 576268 331168
rect 576228 330410 576256 331162
rect 576216 330404 576268 330410
rect 576216 330346 576268 330352
rect 576860 330404 576912 330410
rect 576860 330346 576912 330352
rect 575664 329792 575716 329798
rect 575664 329734 575716 329740
rect 575480 317416 575532 317422
rect 575480 317358 575532 317364
rect 575492 316034 575520 317358
rect 575492 316006 575612 316034
rect 574652 315784 574704 315790
rect 574652 315726 574704 315732
rect 574664 314702 574692 315726
rect 574652 314696 574704 314702
rect 574652 314638 574704 314644
rect 575480 313948 575532 313954
rect 575480 313890 575532 313896
rect 575492 206310 575520 313890
rect 575480 206304 575532 206310
rect 575480 206246 575532 206252
rect 575480 204944 575532 204950
rect 575480 204886 575532 204892
rect 574560 188760 574612 188766
rect 574560 188702 574612 188708
rect 574572 187950 574600 188702
rect 574560 187944 574612 187950
rect 574560 187886 574612 187892
rect 575492 75886 575520 204886
rect 575584 189038 575612 316006
rect 575676 201414 575704 329734
rect 575664 201408 575716 201414
rect 575664 201350 575716 201356
rect 575572 189032 575624 189038
rect 575572 188974 575624 188980
rect 575584 188630 575612 188974
rect 576872 188970 576900 330346
rect 578240 318096 578292 318102
rect 578240 318038 578292 318044
rect 576952 314764 577004 314770
rect 576952 314706 577004 314712
rect 576860 188964 576912 188970
rect 576860 188906 576912 188912
rect 575572 188624 575624 188630
rect 575572 188566 575624 188572
rect 576860 188624 576912 188630
rect 576860 188566 576912 188572
rect 575664 188352 575716 188358
rect 575664 188294 575716 188300
rect 575676 78130 575704 188294
rect 575756 187740 575808 187746
rect 575756 187682 575808 187688
rect 575664 78124 575716 78130
rect 575664 78066 575716 78072
rect 575480 75880 575532 75886
rect 575480 75822 575532 75828
rect 574468 75608 574520 75614
rect 574468 75550 574520 75556
rect 575768 73166 575796 187682
rect 575756 73160 575808 73166
rect 575756 73102 575808 73108
rect 576872 71738 576900 188566
rect 576964 188358 576992 314706
rect 578252 205018 578280 318038
rect 578240 205012 578292 205018
rect 578240 204954 578292 204960
rect 580276 204241 580304 524447
rect 580368 332654 580396 630799
rect 580460 459513 580488 683839
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580920 591025 580948 643991
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580540 485104 580592 485110
rect 580540 485046 580592 485052
rect 580552 484673 580580 485046
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580538 471472 580594 471481
rect 580538 471407 580594 471416
rect 580446 459504 580502 459513
rect 580446 459439 580502 459448
rect 580448 378820 580500 378826
rect 580448 378762 580500 378768
rect 580460 378457 580488 378762
rect 580446 378448 580502 378457
rect 580446 378383 580502 378392
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580356 332648 580408 332654
rect 580356 332590 580408 332596
rect 580262 204232 580318 204241
rect 580262 204167 580318 204176
rect 577136 188964 577188 188970
rect 577136 188906 577188 188912
rect 577044 188420 577096 188426
rect 577044 188362 577096 188368
rect 576952 188352 577004 188358
rect 576952 188294 577004 188300
rect 577056 78198 577084 188362
rect 577044 78192 577096 78198
rect 577044 78134 577096 78140
rect 576860 71732 576912 71738
rect 576860 71674 576912 71680
rect 577148 71670 577176 188906
rect 578240 186992 578292 186998
rect 578240 186934 578292 186940
rect 578252 78062 578280 186934
rect 578240 78056 578292 78062
rect 578240 77998 578292 78004
rect 580460 77994 580488 365055
rect 580552 204105 580580 471407
rect 580644 332489 580672 577623
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 485110 580948 537775
rect 580908 485104 580960 485110
rect 580908 485046 580960 485052
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 378826 580948 431559
rect 580908 378820 580960 378826
rect 580908 378762 580960 378768
rect 580630 332480 580686 332489
rect 580630 332415 580686 332424
rect 580538 204096 580594 204105
rect 580538 204031 580594 204040
rect 580448 77988 580500 77994
rect 580448 77930 580500 77936
rect 577136 71664 577188 71670
rect 577136 71606 577188 71612
rect 574100 22092 574152 22098
rect 574100 22034 574152 22040
rect 570604 22024 570656 22030
rect 570604 21966 570656 21972
rect 368110 21927 368166 21936
rect 378876 21956 378928 21962
rect 360936 21898 360988 21904
rect 378876 21898 378928 21904
rect 400220 21956 400272 21962
rect 400220 21898 400272 21904
rect 342994 21856 343050 21865
rect 342994 21791 343050 21800
rect 338120 10328 338172 10334
rect 338120 10270 338172 10276
rect 331220 4888 331272 4894
rect 331220 4830 331272 4836
rect 302240 3528 302292 3534
rect 302240 3470 302292 3476
rect 266360 3460 266412 3466
rect 266360 3402 266412 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 671200 3478 671256
rect 2778 658144 2834 658200
rect 2870 619112 2926 619168
rect 2778 607144 2834 607200
rect 3422 607144 3478 607200
rect 3422 606056 3478 606112
rect 2778 462576 2834 462632
rect 2778 449520 2834 449576
rect 2870 410488 2926 410544
rect 2778 397432 2834 397488
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 2778 293120 2834 293176
rect 3146 267144 3202 267200
rect 2778 241032 2834 241088
rect 2962 214920 3018 214976
rect 2778 149776 2834 149832
rect 3330 136740 3386 136776
rect 3330 136720 3332 136740
rect 3332 136720 3384 136740
rect 3384 136720 3386 136740
rect 3054 71576 3110 71632
rect 3330 45464 3386 45520
rect 3514 566888 3570 566944
rect 3698 553832 3754 553888
rect 3606 514800 3662 514856
rect 3698 502424 3754 502480
rect 3698 501744 3754 501800
rect 3514 188808 3570 188864
rect 3606 84632 3662 84688
rect 3514 32408 3570 32464
rect 14738 207712 14794 207768
rect 13726 207576 13782 207632
rect 15106 207576 15162 207632
rect 16394 207712 16450 207768
rect 15014 203496 15070 203552
rect 16394 203496 16450 203552
rect 19246 585928 19302 585984
rect 17866 332424 17922 332480
rect 17590 199960 17646 200016
rect 20350 458904 20406 458960
rect 202786 700304 202842 700360
rect 64878 585928 64934 585984
rect 70582 585792 70638 585848
rect 82174 585656 82230 585712
rect 134338 585656 134394 585712
rect 227626 585792 227682 585848
rect 239310 585928 239366 585984
rect 292578 586336 292634 586392
rect 284298 571920 284354 571976
rect 23386 458768 23442 458824
rect 20350 204176 20406 204232
rect 20258 204040 20314 204096
rect 20258 202816 20314 202872
rect 20534 204176 20590 204232
rect 20626 204040 20682 204096
rect 20534 203632 20590 203688
rect 30930 458904 30986 458960
rect 70582 458088 70638 458144
rect 82174 459448 82230 459504
rect 122838 458768 122894 458824
rect 134338 458768 134394 458824
rect 227396 460944 227452 461000
rect 198646 458904 198702 458960
rect 239310 458088 239366 458144
rect 287610 457816 287666 457872
rect 288530 460944 288586 461000
rect 22006 332852 22062 332888
rect 22006 332832 22008 332852
rect 22008 332832 22060 332852
rect 22060 332832 22062 332852
rect 23386 332172 23442 332208
rect 23386 332152 23388 332172
rect 23388 332152 23440 332172
rect 23440 332152 23442 332172
rect 76378 332424 76434 332480
rect 175186 331744 175242 331800
rect 280802 333240 280858 333296
rect 285586 331336 285642 331392
rect 287794 332424 287850 332480
rect 145930 206352 145986 206408
rect 21822 203768 21878 203824
rect 23386 202836 23442 202872
rect 23386 202816 23388 202836
rect 23388 202816 23440 202836
rect 23440 202816 23442 202836
rect 151910 206216 151966 206272
rect 41602 204176 41658 204232
rect 33138 203632 33194 203688
rect 116950 203496 117006 203552
rect 82174 202816 82230 202872
rect 157522 200640 157578 200696
rect 210330 203632 210386 203688
rect 198646 203496 198702 203552
rect 276662 204856 276718 204912
rect 280066 203768 280122 203824
rect 287334 202816 287390 202872
rect 287886 202816 287942 202872
rect 287702 79328 287758 79384
rect 59266 75792 59322 75848
rect 71042 74296 71098 74352
rect 247038 77968 247094 78024
rect 235262 77832 235318 77888
rect 57610 61648 57666 61704
rect 102782 60696 102838 60752
rect 102138 57996 102194 58032
rect 102138 57976 102140 57996
rect 102140 57976 102192 57996
rect 102192 57976 102194 57996
rect 102598 56616 102654 56672
rect 57518 56344 57574 56400
rect 102138 54304 102194 54360
rect 102138 53488 102194 53544
rect 102138 52536 102194 52592
rect 57058 51720 57114 51776
rect 102138 50088 102194 50144
rect 102874 59608 102930 59664
rect 157982 74432 158038 74488
rect 102966 58520 103022 58576
rect 103058 55528 103114 55584
rect 102138 49136 102194 49192
rect 103242 51040 103298 51096
rect 102966 47640 103022 47696
rect 102598 46960 102654 47016
rect 57518 46860 57520 46880
rect 57520 46860 57572 46880
rect 57572 46860 57574 46880
rect 57518 46824 57574 46860
rect 57150 42064 57206 42120
rect 57058 36896 57114 36952
rect 57610 31592 57666 31648
rect 57242 27104 57298 27160
rect 102322 43288 102378 43344
rect 102138 42880 102194 42936
rect 102230 41384 102286 41440
rect 102138 40024 102194 40080
rect 102874 45736 102930 45792
rect 103426 44376 103482 44432
rect 195978 52264 196034 52320
rect 196070 51720 196126 51776
rect 195978 50904 196034 50960
rect 195978 49580 195980 49600
rect 195980 49580 196032 49600
rect 196032 49580 196034 49600
rect 195978 49544 196034 49580
rect 196070 49408 196126 49464
rect 195978 48220 195980 48240
rect 195980 48220 196032 48240
rect 196032 48220 196034 48240
rect 195978 48184 196034 48220
rect 196070 47640 196126 47696
rect 195978 46860 195980 46880
rect 195980 46860 196032 46880
rect 196032 46860 196034 46880
rect 195978 46824 196034 46860
rect 196162 46144 196218 46200
rect 195978 45192 196034 45248
rect 196070 44104 196126 44160
rect 195978 43696 196034 43752
rect 195978 42472 196034 42528
rect 196070 42064 196126 42120
rect 195978 41112 196034 41168
rect 195978 39924 195980 39944
rect 195980 39924 196032 39944
rect 196032 39924 196034 39944
rect 195978 39888 196034 39924
rect 196070 39480 196126 39536
rect 102782 38936 102838 38992
rect 102690 37848 102746 37904
rect 102598 36080 102654 36136
rect 102138 34584 102194 34640
rect 196162 38528 196218 38584
rect 195978 37984 196034 38040
rect 102874 37304 102930 37360
rect 195978 37032 196034 37088
rect 195978 35844 195980 35864
rect 195980 35844 196032 35864
rect 196032 35844 196034 35864
rect 195978 35808 196034 35844
rect 196070 35400 196126 35456
rect 195978 34312 196034 34368
rect 196070 33768 196126 33824
rect 102322 33496 102378 33552
rect 102138 32408 102194 32464
rect 102230 31728 102286 31784
rect 195978 32952 196034 33008
rect 102138 30504 102194 30560
rect 195978 31592 196034 31648
rect 196070 31184 196126 31240
rect 195978 30268 195980 30288
rect 195980 30268 196032 30288
rect 196032 30268 196034 30288
rect 195978 30232 196034 30268
rect 196070 29688 196126 29744
rect 102138 29280 102194 29336
rect 195978 28908 195980 28928
rect 195980 28908 196032 28928
rect 196032 28908 196034 28928
rect 195978 28872 196034 28908
rect 102138 28464 102194 28520
rect 195978 28056 196034 28112
rect 102138 27648 102194 27704
rect 195978 27240 196034 27296
rect 102782 26288 102838 26344
rect 195978 26188 195980 26208
rect 195980 26188 196032 26208
rect 196032 26188 196034 26208
rect 195978 26152 196034 26188
rect 3422 6432 3478 6488
rect 218058 61376 218114 61432
rect 244278 60152 244334 60208
rect 240782 60016 240838 60072
rect 245750 59880 245806 59936
rect 249430 57160 249486 57216
rect 263598 76472 263654 76528
rect 262678 57432 262734 57488
rect 261022 57296 261078 57352
rect 290186 333240 290242 333296
rect 290002 202816 290058 202872
rect 291474 331744 291530 331800
rect 291566 79328 291622 79384
rect 292946 331744 293002 331800
rect 292670 204176 292726 204232
rect 293038 204176 293094 204232
rect 292670 203768 292726 203824
rect 294050 204856 294106 204912
rect 294142 204176 294198 204232
rect 294142 203632 294198 203688
rect 296442 461080 296498 461136
rect 295614 204176 295670 204232
rect 296442 317464 296498 317520
rect 297730 458224 297786 458280
rect 296350 188944 296406 189000
rect 299110 463528 299166 463584
rect 298742 317484 298798 317520
rect 298742 317464 298744 317484
rect 298744 317464 298796 317484
rect 298796 317464 298798 317484
rect 299202 459196 299258 459232
rect 299202 459176 299204 459196
rect 299204 459176 299256 459196
rect 299256 459176 299258 459196
rect 298558 188980 298560 189000
rect 298560 188980 298612 189000
rect 298612 188980 298614 189000
rect 298558 188944 298614 188980
rect 580170 697176 580226 697232
rect 350906 585928 350962 585984
rect 362498 583072 362554 583128
rect 385682 582936 385738 582992
rect 408866 585792 408922 585848
rect 437846 580216 437902 580272
rect 478418 585656 478474 585712
rect 518990 585656 519046 585712
rect 565358 585792 565414 585848
rect 466458 571920 466514 571976
rect 302238 463528 302294 463584
rect 300490 459176 300546 459232
rect 302146 458768 302202 458824
rect 300398 332560 300454 332616
rect 297362 57296 297418 57352
rect 300674 314744 300730 314800
rect 302054 332560 302110 332616
rect 306378 461080 306434 461136
rect 303526 460980 303528 461000
rect 303528 460980 303580 461000
rect 303580 460980 303582 461000
rect 303526 460944 303582 460980
rect 304998 459212 305000 459232
rect 305000 459212 305052 459232
rect 305052 459212 305054 459232
rect 304998 459176 305054 459212
rect 310334 459448 310390 459504
rect 362498 460944 362554 461000
rect 318798 458768 318854 458824
rect 553766 458768 553822 458824
rect 565818 458124 565820 458144
rect 565820 458124 565872 458144
rect 565872 458124 565874 458144
rect 565818 458088 565874 458124
rect 477498 444896 477554 444952
rect 567750 461080 567806 461136
rect 568762 463528 568818 463584
rect 567934 459312 567990 459368
rect 568486 458496 568542 458552
rect 302054 315716 302110 315752
rect 302054 315696 302056 315716
rect 302056 315696 302108 315716
rect 302108 315696 302110 315716
rect 302054 204720 302110 204776
rect 303526 332188 303528 332208
rect 303528 332188 303580 332208
rect 303580 332188 303582 332208
rect 303526 332152 303582 332188
rect 310334 332424 310390 332480
rect 553766 331744 553822 331800
rect 565818 332288 565874 332344
rect 567474 315716 567530 315752
rect 567474 315696 567476 315716
rect 567476 315696 567528 315716
rect 567528 315696 567530 315716
rect 568486 314628 568542 314664
rect 568486 314608 568488 314628
rect 568488 314608 568540 314628
rect 568540 314608 568542 314628
rect 303526 201320 303582 201376
rect 302882 186360 302938 186416
rect 304538 204176 304594 204232
rect 310334 204040 310390 204096
rect 419538 188944 419594 189000
rect 567290 204332 567346 204368
rect 567290 204312 567292 204332
rect 567292 204312 567344 204332
rect 567344 204312 567346 204332
rect 518806 187584 518862 187640
rect 303710 185544 303766 185600
rect 302330 79872 302386 79928
rect 304538 75928 304594 75984
rect 303802 61376 303858 61432
rect 321926 59200 321982 59256
rect 327078 58520 327134 58576
rect 328366 58520 328422 58576
rect 335358 66816 335414 66872
rect 336646 66816 336702 66872
rect 374182 76472 374238 76528
rect 389178 76608 389234 76664
rect 386878 57296 386934 57352
rect 388534 57160 388590 57216
rect 518990 75792 519046 75848
rect 507122 74432 507178 74488
rect 400218 54440 400274 54496
rect 368110 21936 368166 21992
rect 389638 22072 389694 22128
rect 570234 336640 570290 336696
rect 571430 458496 571486 458552
rect 572810 331744 572866 331800
rect 580446 683848 580502 683904
rect 580354 630808 580410 630864
rect 580262 524456 580318 524512
rect 580906 644000 580962 644056
rect 580906 590960 580962 591016
rect 580630 577632 580686 577688
rect 580538 484608 580594 484664
rect 580538 471416 580594 471472
rect 580446 459448 580502 459504
rect 580446 378392 580502 378448
rect 580446 365064 580502 365120
rect 580262 204176 580318 204232
rect 580906 537784 580962 537840
rect 580906 431568 580962 431624
rect 580630 332424 580686 332480
rect 580538 204040 580594 204096
rect 342994 21800 343050 21856
<< metal3 >>
rect 202781 700362 202847 700365
rect 295926 700362 295932 700364
rect 202781 700360 295932 700362
rect 202781 700304 202786 700360
rect 202842 700304 295932 700360
rect 202781 700302 295932 700304
rect 202781 700299 202847 700302
rect 295926 700300 295932 700302
rect 295996 700300 296002 700364
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580441 683906 580507 683909
rect 583520 683906 584960 683996
rect 580441 683904 584960 683906
rect 580441 683848 580446 683904
rect 580502 683848 584960 683904
rect 580441 683846 584960 683848
rect 580441 683843 580507 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2865 619170 2931 619173
rect -960 619168 2931 619170
rect -960 619112 2870 619168
rect 2926 619112 2931 619168
rect -960 619110 2931 619112
rect -960 619020 480 619110
rect 2865 619107 2931 619110
rect 583520 617388 584960 617628
rect 2773 607202 2839 607205
rect 3417 607202 3483 607205
rect 2773 607200 3483 607202
rect 2773 607144 2778 607200
rect 2834 607144 3422 607200
rect 3478 607144 3483 607200
rect 2773 607142 3483 607144
rect 2773 607139 2839 607142
rect 3417 607139 3483 607142
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 569534 590956 569540 591020
rect 569604 591018 569610 591020
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 569604 591016 584960 591018
rect 569604 590960 580906 591016
rect 580962 590960 584960 591016
rect 569604 590958 584960 590960
rect 569604 590956 569610 590958
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect 292573 586396 292639 586397
rect 292573 586394 292620 586396
rect 292528 586392 292620 586394
rect 292528 586336 292578 586392
rect 292528 586334 292620 586336
rect 292573 586332 292620 586334
rect 292684 586332 292690 586396
rect 292573 586331 292639 586332
rect 19241 585986 19307 585989
rect 64873 585986 64939 585989
rect 19241 585984 64939 585986
rect 19241 585928 19246 585984
rect 19302 585928 64878 585984
rect 64934 585928 64939 585984
rect 19241 585926 64939 585928
rect 19241 585923 19307 585926
rect 64873 585923 64939 585926
rect 239305 585986 239371 585989
rect 285622 585986 285628 585988
rect 239305 585984 285628 585986
rect 239305 585928 239310 585984
rect 239366 585928 285628 585984
rect 239305 585926 285628 585928
rect 239305 585923 239371 585926
rect 285622 585924 285628 585926
rect 285692 585924 285698 585988
rect 303470 585924 303476 585988
rect 303540 585986 303546 585988
rect 350901 585986 350967 585989
rect 303540 585984 350967 585986
rect 303540 585928 350906 585984
rect 350962 585928 350967 585984
rect 303540 585926 350967 585928
rect 303540 585924 303546 585926
rect 350901 585923 350967 585926
rect 23238 585788 23244 585852
rect 23308 585850 23314 585852
rect 70577 585850 70643 585853
rect 23308 585848 70643 585850
rect 23308 585792 70582 585848
rect 70638 585792 70643 585848
rect 23308 585790 70643 585792
rect 23308 585788 23314 585790
rect 70577 585787 70643 585790
rect 227621 585850 227687 585853
rect 287094 585850 287100 585852
rect 227621 585848 287100 585850
rect 227621 585792 227626 585848
rect 227682 585792 287100 585848
rect 227621 585790 287100 585792
rect 227621 585787 227687 585790
rect 287094 585788 287100 585790
rect 287164 585788 287170 585852
rect 299974 585788 299980 585852
rect 300044 585850 300050 585852
rect 408861 585850 408927 585853
rect 300044 585848 408927 585850
rect 300044 585792 408866 585848
rect 408922 585792 408927 585848
rect 300044 585790 408927 585792
rect 300044 585788 300050 585790
rect 408861 585787 408927 585790
rect 565353 585850 565419 585853
rect 570086 585850 570092 585852
rect 565353 585848 570092 585850
rect 565353 585792 565358 585848
rect 565414 585792 570092 585848
rect 565353 585790 570092 585792
rect 565353 585787 565419 585790
rect 570086 585788 570092 585790
rect 570156 585788 570162 585852
rect 21950 585652 21956 585716
rect 22020 585714 22026 585716
rect 82169 585714 82235 585717
rect 22020 585712 82235 585714
rect 22020 585656 82174 585712
rect 82230 585656 82235 585712
rect 22020 585654 82235 585656
rect 22020 585652 22026 585654
rect 82169 585651 82235 585654
rect 134333 585714 134399 585717
rect 288382 585714 288388 585716
rect 134333 585712 288388 585714
rect 134333 585656 134338 585712
rect 134394 585656 288388 585712
rect 134333 585654 288388 585656
rect 134333 585651 134399 585654
rect 288382 585652 288388 585654
rect 288452 585652 288458 585716
rect 291694 585652 291700 585716
rect 291764 585714 291770 585716
rect 478413 585714 478479 585717
rect 291764 585712 478479 585714
rect 291764 585656 478418 585712
rect 478474 585656 478479 585712
rect 291764 585654 478479 585656
rect 291764 585652 291770 585654
rect 478413 585651 478479 585654
rect 518985 585714 519051 585717
rect 565854 585714 565860 585716
rect 518985 585712 565860 585714
rect 518985 585656 518990 585712
rect 519046 585656 565860 585712
rect 518985 585654 565860 585656
rect 518985 585651 519051 585654
rect 565854 585652 565860 585654
rect 565924 585652 565930 585716
rect 301998 583068 302004 583132
rect 302068 583130 302074 583132
rect 362493 583130 362559 583133
rect 302068 583128 362559 583130
rect 302068 583072 362498 583128
rect 362554 583072 362559 583128
rect 302068 583070 362559 583072
rect 302068 583068 302074 583070
rect 362493 583067 362559 583070
rect 298686 582932 298692 582996
rect 298756 582994 298762 582996
rect 385677 582994 385743 582997
rect 298756 582992 385743 582994
rect 298756 582936 385682 582992
rect 385738 582936 385743 582992
rect 298756 582934 385743 582936
rect 298756 582932 298762 582934
rect 385677 582931 385743 582934
rect 437841 580274 437907 580277
rect 568614 580274 568620 580276
rect 437841 580272 568620 580274
rect 437841 580216 437846 580272
rect 437902 580216 568620 580272
rect 437841 580214 568620 580216
rect 437841 580211 437907 580214
rect 568614 580212 568620 580214
rect 568684 580212 568690 580276
rect -960 579852 480 580092
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect 284293 571978 284359 571981
rect 297214 571978 297220 571980
rect 284293 571976 297220 571978
rect 284293 571920 284298 571976
rect 284354 571920 297220 571976
rect 284293 571918 297220 571920
rect 284293 571915 284359 571918
rect 297214 571916 297220 571918
rect 297284 571916 297290 571980
rect 466453 571978 466519 571981
rect 567878 571978 567884 571980
rect 466453 571976 567884 571978
rect 466453 571920 466458 571976
rect 466514 571920 567884 571976
rect 466453 571918 567884 571920
rect 466453 571915 466519 571918
rect 567878 571916 567884 571918
rect 567948 571916 567954 571980
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 580257 524514 580323 524517
rect 583520 524514 584960 524604
rect 580257 524512 584960 524514
rect 580257 524456 580262 524512
rect 580318 524456 584960 524512
rect 580257 524454 584960 524456
rect 580257 524451 580323 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 583520 511172 584960 511412
rect 3693 502482 3759 502485
rect 18454 502482 18460 502484
rect 3693 502480 18460 502482
rect 3693 502424 3698 502480
rect 3754 502424 18460 502480
rect 3693 502422 18460 502424
rect 3693 502419 3759 502422
rect 18454 502420 18460 502422
rect 18524 502420 18530 502484
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 580533 471474 580599 471477
rect 583520 471474 584960 471564
rect 580533 471472 584960 471474
rect 580533 471416 580538 471472
rect 580594 471416 584960 471472
rect 580533 471414 584960 471416
rect 580533 471411 580599 471414
rect 583520 471324 584960 471414
rect 299105 463586 299171 463589
rect 302233 463586 302299 463589
rect 299105 463584 302299 463586
rect 299105 463528 299110 463584
rect 299166 463528 302238 463584
rect 302294 463528 302299 463584
rect 299105 463526 302299 463528
rect 299105 463523 299171 463526
rect 302233 463523 302299 463526
rect 568614 463524 568620 463588
rect 568684 463586 568690 463588
rect 568757 463586 568823 463589
rect 568684 463584 568823 463586
rect 568684 463528 568762 463584
rect 568818 463528 568823 463584
rect 568684 463526 568823 463528
rect 568684 463524 568690 463526
rect 568757 463523 568823 463526
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 301998 461212 302004 461276
rect 302068 461274 302074 461276
rect 302068 461214 316050 461274
rect 302068 461212 302074 461214
rect 296437 461138 296503 461141
rect 306373 461138 306439 461141
rect 296437 461136 306439 461138
rect 296437 461080 296442 461136
rect 296498 461080 306378 461136
rect 306434 461080 306439 461136
rect 296437 461078 306439 461080
rect 296437 461075 296503 461078
rect 306373 461075 306439 461078
rect 227391 461002 227457 461005
rect 287094 461002 287100 461004
rect 227391 461000 287100 461002
rect 227391 460944 227396 461000
rect 227452 460944 287100 461000
rect 227391 460942 287100 460944
rect 227391 460939 227457 460942
rect 287094 460940 287100 460942
rect 287164 461002 287170 461004
rect 288525 461002 288591 461005
rect 303521 461004 303587 461005
rect 287164 461000 288591 461002
rect 287164 460944 288530 461000
rect 288586 460944 288591 461000
rect 287164 460942 288591 460944
rect 287164 460940 287170 460942
rect 288525 460939 288591 460942
rect 303470 460940 303476 461004
rect 303540 461002 303587 461004
rect 315990 461002 316050 461214
rect 567745 461140 567811 461141
rect 567694 461138 567700 461140
rect 567654 461078 567700 461138
rect 567764 461136 567811 461140
rect 567806 461080 567811 461136
rect 567694 461076 567700 461078
rect 567764 461076 567811 461080
rect 567745 461075 567811 461076
rect 362493 461002 362559 461005
rect 303540 461000 303632 461002
rect 303582 460944 303632 461000
rect 303540 460942 303632 460944
rect 315990 461000 362559 461002
rect 315990 460944 362498 461000
rect 362554 460944 362559 461000
rect 315990 460942 362559 460944
rect 303540 460940 303587 460942
rect 303521 460939 303587 460940
rect 362493 460939 362559 460942
rect 21950 459444 21956 459508
rect 22020 459506 22026 459508
rect 82169 459506 82235 459509
rect 22020 459504 82235 459506
rect 22020 459448 82174 459504
rect 82230 459448 82235 459504
rect 22020 459446 82235 459448
rect 22020 459444 22026 459446
rect 82169 459443 82235 459446
rect 310329 459506 310395 459509
rect 580441 459506 580507 459509
rect 310329 459504 580507 459506
rect 310329 459448 310334 459504
rect 310390 459448 580446 459504
rect 580502 459448 580507 459504
rect 310329 459446 580507 459448
rect 310329 459443 310395 459446
rect 580441 459443 580507 459446
rect 567929 459372 567995 459373
rect 567878 459370 567884 459372
rect 567838 459310 567884 459370
rect 567948 459368 567995 459372
rect 567990 459312 567995 459368
rect 567878 459308 567884 459310
rect 567948 459308 567995 459312
rect 567929 459307 567995 459308
rect 298686 459172 298692 459236
rect 298756 459234 298762 459236
rect 299197 459234 299263 459237
rect 298756 459232 299263 459234
rect 298756 459176 299202 459232
rect 299258 459176 299263 459232
rect 298756 459174 299263 459176
rect 298756 459172 298762 459174
rect 299197 459171 299263 459174
rect 300485 459234 300551 459237
rect 304993 459234 305059 459237
rect 300485 459232 305059 459234
rect 300485 459176 300490 459232
rect 300546 459176 304998 459232
rect 305054 459176 305059 459232
rect 300485 459174 305059 459176
rect 300485 459171 300551 459174
rect 304993 459171 305059 459174
rect 20345 458962 20411 458965
rect 30925 458962 30991 458965
rect 20345 458960 30991 458962
rect 20345 458904 20350 458960
rect 20406 458904 30930 458960
rect 30986 458904 30991 458960
rect 20345 458902 30991 458904
rect 20345 458899 20411 458902
rect 30925 458899 30991 458902
rect 198641 458962 198707 458965
rect 291142 458962 291148 458964
rect 198641 458960 291148 458962
rect 198641 458904 198646 458960
rect 198702 458904 291148 458960
rect 198641 458902 291148 458904
rect 198641 458899 198707 458902
rect 291142 458900 291148 458902
rect 291212 458900 291218 458964
rect 23381 458826 23447 458829
rect 122833 458826 122899 458829
rect 23381 458824 122899 458826
rect 23381 458768 23386 458824
rect 23442 458768 122838 458824
rect 122894 458768 122899 458824
rect 23381 458766 122899 458768
rect 23381 458763 23447 458766
rect 122833 458763 122899 458766
rect 134333 458826 134399 458829
rect 289854 458826 289860 458828
rect 134333 458824 289860 458826
rect 134333 458768 134338 458824
rect 134394 458768 289860 458824
rect 134333 458766 289860 458768
rect 134333 458763 134399 458766
rect 289854 458764 289860 458766
rect 289924 458764 289930 458828
rect 302141 458826 302207 458829
rect 318793 458826 318859 458829
rect 302141 458824 318859 458826
rect 302141 458768 302146 458824
rect 302202 458768 318798 458824
rect 318854 458768 318859 458824
rect 302141 458766 318859 458768
rect 302141 458763 302207 458766
rect 318793 458763 318859 458766
rect 553761 458826 553827 458829
rect 571374 458826 571380 458828
rect 553761 458824 571380 458826
rect 553761 458768 553766 458824
rect 553822 458768 571380 458824
rect 553761 458766 571380 458768
rect 553761 458763 553827 458766
rect 571374 458764 571380 458766
rect 571444 458764 571450 458828
rect 568481 458554 568547 458557
rect 571425 458554 571491 458557
rect 568481 458552 571491 458554
rect 568481 458496 568486 458552
rect 568542 458496 571430 458552
rect 571486 458496 571491 458552
rect 568481 458494 571491 458496
rect 568481 458491 568547 458494
rect 571425 458491 571491 458494
rect 297725 458282 297791 458285
rect 298686 458282 298692 458284
rect 297725 458280 298692 458282
rect 297725 458224 297730 458280
rect 297786 458224 298692 458280
rect 297725 458222 298692 458224
rect 297725 458219 297791 458222
rect 298686 458220 298692 458222
rect 298756 458220 298762 458284
rect 23238 458084 23244 458148
rect 23308 458146 23314 458148
rect 70577 458146 70643 458149
rect 23308 458144 70643 458146
rect 23308 458088 70582 458144
rect 70638 458088 70643 458144
rect 23308 458086 70643 458088
rect 23308 458084 23314 458086
rect 70577 458083 70643 458086
rect 239305 458146 239371 458149
rect 285622 458146 285628 458148
rect 239305 458144 285628 458146
rect 239305 458088 239310 458144
rect 239366 458088 285628 458144
rect 239305 458086 285628 458088
rect 239305 458083 239371 458086
rect 285622 458084 285628 458086
rect 285692 458084 285698 458148
rect 565813 458146 565879 458149
rect 566406 458146 566412 458148
rect 565813 458144 566412 458146
rect 565813 458088 565818 458144
rect 565874 458088 566412 458144
rect 565813 458086 566412 458088
rect 565813 458083 565879 458086
rect 566406 458084 566412 458086
rect 566476 458084 566482 458148
rect 583520 457996 584960 458236
rect 287605 457876 287671 457877
rect 287605 457874 287652 457876
rect 287560 457872 287652 457874
rect 287560 457816 287610 457872
rect 287560 457814 287652 457816
rect 287605 457812 287652 457814
rect 287716 457812 287722 457876
rect 287605 457811 287671 457812
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 286174 444892 286180 444956
rect 286244 444954 286250 444956
rect 477493 444954 477559 444957
rect 286244 444952 477559 444954
rect 286244 444896 477498 444952
rect 477554 444896 477559 444952
rect 286244 444894 477559 444896
rect 286244 444892 286250 444894
rect 477493 444891 477559 444894
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 570454 418236 570460 418300
rect 570524 418298 570530 418300
rect 583520 418298 584960 418388
rect 570524 418238 584960 418298
rect 570524 418236 570530 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580441 378450 580507 378453
rect 583520 378450 584960 378540
rect 580441 378448 584960 378450
rect 580441 378392 580446 378448
rect 580502 378392 584960 378448
rect 580441 378390 584960 378392
rect 580441 378387 580507 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect 568430 336636 568436 336700
rect 568500 336698 568506 336700
rect 570229 336698 570295 336701
rect 568500 336696 570295 336698
rect 568500 336640 570234 336696
rect 570290 336640 570295 336696
rect 568500 336638 570295 336640
rect 568500 336636 568506 336638
rect 570229 336635 570295 336638
rect 280797 333298 280863 333301
rect 290181 333298 290247 333301
rect 280797 333296 290247 333298
rect 280797 333240 280802 333296
rect 280858 333240 290186 333296
rect 290242 333240 290247 333296
rect 280797 333238 290247 333240
rect 280797 333235 280863 333238
rect 290181 333235 290247 333238
rect 21214 332828 21220 332892
rect 21284 332890 21290 332892
rect 22001 332890 22067 332893
rect 21284 332888 22067 332890
rect 21284 332832 22006 332888
rect 22062 332832 22067 332888
rect 21284 332830 22067 332832
rect 21284 332828 21290 332830
rect 22001 332827 22067 332830
rect 300393 332618 300459 332621
rect 300894 332618 300900 332620
rect 300393 332616 300900 332618
rect 300393 332560 300398 332616
rect 300454 332560 300900 332616
rect 300393 332558 300900 332560
rect 300393 332555 300459 332558
rect 300894 332556 300900 332558
rect 300964 332618 300970 332620
rect 302049 332618 302115 332621
rect 300964 332616 302115 332618
rect 300964 332560 302054 332616
rect 302110 332560 302115 332616
rect 300964 332558 302115 332560
rect 300964 332556 300970 332558
rect 302049 332555 302115 332558
rect 17861 332482 17927 332485
rect 76373 332482 76439 332485
rect 17861 332480 76439 332482
rect -960 332196 480 332436
rect 17861 332424 17866 332480
rect 17922 332424 76378 332480
rect 76434 332424 76439 332480
rect 17861 332422 76439 332424
rect 17861 332419 17927 332422
rect 76373 332419 76439 332422
rect 287789 332482 287855 332485
rect 288198 332482 288204 332484
rect 287789 332480 288204 332482
rect 287789 332424 287794 332480
rect 287850 332424 288204 332480
rect 287789 332422 288204 332424
rect 287789 332419 287855 332422
rect 288198 332420 288204 332422
rect 288268 332420 288274 332484
rect 310329 332482 310395 332485
rect 580625 332482 580691 332485
rect 310329 332480 580691 332482
rect 310329 332424 310334 332480
rect 310390 332424 580630 332480
rect 580686 332424 580691 332480
rect 310329 332422 580691 332424
rect 310329 332419 310395 332422
rect 580625 332419 580691 332422
rect 565813 332348 565879 332349
rect 565813 332346 565860 332348
rect 565768 332344 565860 332346
rect 565768 332288 565818 332344
rect 565768 332286 565860 332288
rect 565813 332284 565860 332286
rect 565924 332284 565930 332348
rect 565813 332283 565879 332284
rect 22686 332148 22692 332212
rect 22756 332210 22762 332212
rect 23381 332210 23447 332213
rect 22756 332208 23447 332210
rect 22756 332152 23386 332208
rect 23442 332152 23447 332208
rect 22756 332150 23447 332152
rect 22756 332148 22762 332150
rect 23381 332147 23447 332150
rect 302734 332148 302740 332212
rect 302804 332210 302810 332212
rect 303521 332210 303587 332213
rect 302804 332208 303587 332210
rect 302804 332152 303526 332208
rect 303582 332152 303587 332208
rect 302804 332150 303587 332152
rect 302804 332148 302810 332150
rect 303521 332147 303587 332150
rect 175181 331802 175247 331805
rect 291469 331802 291535 331805
rect 292941 331802 293007 331805
rect 175181 331800 293007 331802
rect 175181 331744 175186 331800
rect 175242 331744 291474 331800
rect 291530 331744 292946 331800
rect 293002 331744 293007 331800
rect 175181 331742 293007 331744
rect 175181 331739 175247 331742
rect 291469 331739 291535 331742
rect 292941 331739 293007 331742
rect 553761 331802 553827 331805
rect 572805 331802 572871 331805
rect 553761 331800 572871 331802
rect 553761 331744 553766 331800
rect 553822 331744 572810 331800
rect 572866 331744 572871 331800
rect 553761 331742 572871 331744
rect 553761 331739 553827 331742
rect 572805 331739 572871 331742
rect 285581 331396 285647 331397
rect 285581 331392 285628 331396
rect 285692 331394 285698 331396
rect 285581 331336 285586 331392
rect 285581 331332 285628 331336
rect 285692 331334 285738 331394
rect 285692 331332 285698 331334
rect 285581 331331 285647 331332
rect 583520 325124 584960 325364
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 296437 317522 296503 317525
rect 298737 317524 298803 317525
rect 298686 317522 298692 317524
rect 296437 317520 298692 317522
rect 298756 317520 298803 317524
rect 296437 317464 296442 317520
rect 296498 317464 298692 317520
rect 298798 317464 298803 317520
rect 296437 317462 298692 317464
rect 296437 317459 296503 317462
rect 298686 317460 298692 317462
rect 298756 317460 298803 317464
rect 298737 317459 298803 317460
rect 302049 315756 302115 315757
rect 301998 315692 302004 315756
rect 302068 315754 302115 315756
rect 567469 315754 567535 315757
rect 567694 315754 567700 315756
rect 302068 315752 302160 315754
rect 302110 315696 302160 315752
rect 302068 315694 302160 315696
rect 567469 315752 567700 315754
rect 567469 315696 567474 315752
rect 567530 315696 567700 315752
rect 567469 315694 567700 315696
rect 302068 315692 302115 315694
rect 302049 315691 302115 315692
rect 567469 315691 567535 315694
rect 567694 315692 567700 315694
rect 567764 315692 567770 315756
rect 300669 314802 300735 314805
rect 301998 314802 302004 314804
rect 300669 314800 302004 314802
rect 300669 314744 300674 314800
rect 300730 314744 302004 314800
rect 300669 314742 302004 314744
rect 300669 314739 300735 314742
rect 301998 314740 302004 314742
rect 302068 314740 302074 314804
rect 568481 314668 568547 314669
rect 568430 314666 568436 314668
rect 568390 314606 568436 314666
rect 568500 314664 568547 314668
rect 568542 314608 568547 314664
rect 568430 314604 568436 314606
rect 568500 314604 568547 314608
rect 568481 314603 568547 314604
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214978 480 215068
rect 2957 214978 3023 214981
rect -960 214976 3023 214978
rect -960 214920 2962 214976
rect 3018 214920 3023 214976
rect -960 214918 3023 214920
rect -960 214828 480 214918
rect 2957 214915 3023 214918
rect 14733 207770 14799 207773
rect 16389 207770 16455 207773
rect 21398 207770 21404 207772
rect 14733 207768 21404 207770
rect 14733 207712 14738 207768
rect 14794 207712 16394 207768
rect 16450 207712 21404 207768
rect 14733 207710 21404 207712
rect 14733 207707 14799 207710
rect 16389 207707 16455 207710
rect 21398 207708 21404 207710
rect 21468 207708 21474 207772
rect 13721 207634 13787 207637
rect 15101 207634 15167 207637
rect 22134 207634 22140 207636
rect 13721 207632 22140 207634
rect 13721 207576 13726 207632
rect 13782 207576 15106 207632
rect 15162 207576 22140 207632
rect 13721 207574 22140 207576
rect 13721 207571 13787 207574
rect 15101 207571 15167 207574
rect 22134 207572 22140 207574
rect 22204 207572 22210 207636
rect 22134 206348 22140 206412
rect 22204 206410 22210 206412
rect 145925 206410 145991 206413
rect 22204 206408 145991 206410
rect 22204 206352 145930 206408
rect 145986 206352 145991 206408
rect 22204 206350 145991 206352
rect 22204 206348 22210 206350
rect 145925 206347 145991 206350
rect 21398 206212 21404 206276
rect 21468 206274 21474 206276
rect 151905 206274 151971 206277
rect 21468 206272 151971 206274
rect 21468 206216 151910 206272
rect 151966 206216 151971 206272
rect 21468 206214 151971 206216
rect 21468 206212 21474 206214
rect 151905 206211 151971 206214
rect 583520 205580 584960 205820
rect 276657 204914 276723 204917
rect 294045 204914 294111 204917
rect 276657 204912 294111 204914
rect 276657 204856 276662 204912
rect 276718 204856 294050 204912
rect 294106 204856 294111 204912
rect 276657 204854 294111 204856
rect 276657 204851 276723 204854
rect 294045 204851 294111 204854
rect 302049 204780 302115 204781
rect 300894 204716 300900 204780
rect 300964 204778 300970 204780
rect 301998 204778 302004 204780
rect 300964 204718 302004 204778
rect 302068 204778 302115 204780
rect 302068 204776 302196 204778
rect 302110 204720 302196 204776
rect 300964 204716 300970 204718
rect 301998 204716 302004 204718
rect 302068 204718 302196 204720
rect 302068 204716 302115 204718
rect 302049 204715 302115 204716
rect 567285 204372 567351 204373
rect 567285 204370 567332 204372
rect 567240 204368 567332 204370
rect 567240 204312 567290 204368
rect 567240 204310 567332 204312
rect 567285 204308 567332 204310
rect 567396 204308 567402 204372
rect 567285 204307 567351 204308
rect 20345 204234 20411 204237
rect 20529 204234 20595 204237
rect 41597 204234 41663 204237
rect 20345 204232 20595 204234
rect 20345 204176 20350 204232
rect 20406 204176 20534 204232
rect 20590 204176 20595 204232
rect 20345 204174 20595 204176
rect 20345 204171 20411 204174
rect 20529 204171 20595 204174
rect 26190 204232 41663 204234
rect 26190 204176 41602 204232
rect 41658 204176 41663 204232
rect 26190 204174 41663 204176
rect 20253 204098 20319 204101
rect 20621 204098 20687 204101
rect 26190 204098 26250 204174
rect 41597 204171 41663 204174
rect 292665 204234 292731 204237
rect 293033 204234 293099 204237
rect 292665 204232 293099 204234
rect 292665 204176 292670 204232
rect 292726 204176 293038 204232
rect 293094 204176 293099 204232
rect 292665 204174 293099 204176
rect 292665 204171 292731 204174
rect 293033 204171 293099 204174
rect 294137 204234 294203 204237
rect 295609 204234 295675 204237
rect 294137 204232 295675 204234
rect 294137 204176 294142 204232
rect 294198 204176 295614 204232
rect 295670 204176 295675 204232
rect 294137 204174 295675 204176
rect 294137 204171 294203 204174
rect 295609 204171 295675 204174
rect 304533 204234 304599 204237
rect 580257 204234 580323 204237
rect 304533 204232 580323 204234
rect 304533 204176 304538 204232
rect 304594 204176 580262 204232
rect 580318 204176 580323 204232
rect 304533 204174 580323 204176
rect 304533 204171 304599 204174
rect 580257 204171 580323 204174
rect 20253 204096 26250 204098
rect 20253 204040 20258 204096
rect 20314 204040 20626 204096
rect 20682 204040 26250 204096
rect 20253 204038 26250 204040
rect 310329 204098 310395 204101
rect 580533 204098 580599 204101
rect 310329 204096 580599 204098
rect 310329 204040 310334 204096
rect 310390 204040 580538 204096
rect 580594 204040 580599 204096
rect 310329 204038 580599 204040
rect 20253 204035 20319 204038
rect 20621 204035 20687 204038
rect 310329 204035 310395 204038
rect 580533 204035 580599 204038
rect 21817 203826 21883 203829
rect 21950 203826 21956 203828
rect 21817 203824 21956 203826
rect 21817 203768 21822 203824
rect 21878 203768 21956 203824
rect 21817 203766 21956 203768
rect 21817 203763 21883 203766
rect 21950 203764 21956 203766
rect 22020 203764 22026 203828
rect 280061 203826 280127 203829
rect 292665 203826 292731 203829
rect 280061 203824 292731 203826
rect 280061 203768 280066 203824
rect 280122 203768 292670 203824
rect 292726 203768 292731 203824
rect 280061 203766 292731 203768
rect 280061 203763 280127 203766
rect 292665 203763 292731 203766
rect 20529 203690 20595 203693
rect 33133 203690 33199 203693
rect 20529 203688 33199 203690
rect 20529 203632 20534 203688
rect 20590 203632 33138 203688
rect 33194 203632 33199 203688
rect 20529 203630 33199 203632
rect 20529 203627 20595 203630
rect 33133 203627 33199 203630
rect 210325 203690 210391 203693
rect 294137 203690 294203 203693
rect 210325 203688 294203 203690
rect 210325 203632 210330 203688
rect 210386 203632 294142 203688
rect 294198 203632 294203 203688
rect 210325 203630 294203 203632
rect 210325 203627 210391 203630
rect 294137 203627 294203 203630
rect 15009 203554 15075 203557
rect 16389 203554 16455 203557
rect 116945 203554 117011 203557
rect 15009 203552 117011 203554
rect 15009 203496 15014 203552
rect 15070 203496 16394 203552
rect 16450 203496 116950 203552
rect 117006 203496 117011 203552
rect 15009 203494 117011 203496
rect 15009 203491 15075 203494
rect 16389 203491 16455 203494
rect 116945 203491 117011 203494
rect 198641 203554 198707 203557
rect 287094 203554 287100 203556
rect 198641 203552 287100 203554
rect 198641 203496 198646 203552
rect 198702 203496 287100 203552
rect 198641 203494 287100 203496
rect 198641 203491 198707 203494
rect 287094 203492 287100 203494
rect 287164 203492 287170 203556
rect 20253 202874 20319 202877
rect 21214 202874 21220 202876
rect 20253 202872 21220 202874
rect 20253 202816 20258 202872
rect 20314 202816 21220 202872
rect 20253 202814 21220 202816
rect 20253 202811 20319 202814
rect 21214 202812 21220 202814
rect 21284 202812 21290 202876
rect 22686 202812 22692 202876
rect 22756 202874 22762 202876
rect 23381 202874 23447 202877
rect 82169 202874 82235 202877
rect 287329 202876 287395 202877
rect 287278 202874 287284 202876
rect 22756 202872 23447 202874
rect 22756 202816 23386 202872
rect 23442 202816 23447 202872
rect 22756 202814 23447 202816
rect 22756 202812 22762 202814
rect 21222 202738 21282 202812
rect 23381 202811 23447 202814
rect 26190 202872 82235 202874
rect 26190 202816 82174 202872
rect 82230 202816 82235 202872
rect 26190 202814 82235 202816
rect 287238 202814 287284 202874
rect 287348 202872 287395 202876
rect 287390 202816 287395 202872
rect 26190 202738 26250 202814
rect 82169 202811 82235 202814
rect 287278 202812 287284 202814
rect 287348 202812 287395 202816
rect 287329 202811 287395 202812
rect 287881 202874 287947 202877
rect 288198 202874 288204 202876
rect 287881 202872 288204 202874
rect 287881 202816 287886 202872
rect 287942 202816 288204 202872
rect 287881 202814 288204 202816
rect 287881 202811 287947 202814
rect 288198 202812 288204 202814
rect 288268 202874 288274 202876
rect 289997 202874 290063 202877
rect 288268 202872 290063 202874
rect 288268 202816 290002 202872
rect 290058 202816 290063 202872
rect 288268 202814 290063 202816
rect 288268 202812 288274 202814
rect 289997 202811 290063 202814
rect 21222 202678 26250 202738
rect -960 201772 480 202012
rect 302734 201316 302740 201380
rect 302804 201378 302810 201380
rect 303521 201378 303587 201381
rect 302804 201376 303587 201378
rect 302804 201320 303526 201376
rect 303582 201320 303587 201376
rect 302804 201318 303587 201320
rect 302804 201316 302810 201318
rect 303521 201315 303587 201318
rect 157517 200698 157583 200701
rect 19290 200696 157583 200698
rect 19290 200640 157522 200696
rect 157578 200640 157583 200696
rect 19290 200638 157583 200640
rect 17585 200018 17651 200021
rect 19290 200018 19350 200638
rect 157517 200635 157583 200638
rect 19926 200018 19932 200020
rect 17585 200016 19932 200018
rect 17585 199960 17590 200016
rect 17646 199960 19932 200016
rect 17585 199958 19932 199960
rect 17585 199955 17651 199958
rect 19926 199956 19932 199958
rect 19996 199956 20002 200020
rect 583520 192388 584960 192628
rect 296345 189002 296411 189005
rect 298553 189002 298619 189005
rect 296345 189000 298619 189002
rect -960 188866 480 188956
rect 296345 188944 296350 189000
rect 296406 188944 298558 189000
rect 298614 188944 298619 189000
rect 296345 188942 298619 188944
rect 296345 188939 296411 188942
rect 298510 188939 298619 188942
rect 298686 188940 298692 189004
rect 298756 189002 298762 189004
rect 419533 189002 419599 189005
rect 298756 189000 419599 189002
rect 298756 188944 419538 189000
rect 419594 188944 419599 189000
rect 298756 188942 419599 188944
rect 298756 188940 298762 188942
rect 419533 188939 419599 188942
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect 298510 188866 298570 188939
rect 298870 188866 298876 188868
rect 298510 188806 298876 188866
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 298870 188804 298876 188806
rect 298940 188804 298946 188868
rect 518801 187642 518867 187645
rect 565854 187642 565860 187644
rect 518801 187640 565860 187642
rect 518801 187584 518806 187640
rect 518862 187584 565860 187640
rect 518801 187582 565860 187584
rect 518801 187579 518867 187582
rect 565854 187580 565860 187582
rect 565924 187580 565930 187644
rect 301446 186356 301452 186420
rect 301516 186418 301522 186420
rect 302877 186418 302943 186421
rect 301516 186416 302943 186418
rect 301516 186360 302882 186416
rect 302938 186360 302943 186416
rect 301516 186358 302943 186360
rect 301516 186356 301522 186358
rect 302877 186355 302943 186358
rect 299238 185540 299244 185604
rect 299308 185602 299314 185604
rect 303705 185602 303771 185605
rect 299308 185600 303771 185602
rect 299308 185544 303710 185600
rect 303766 185544 303771 185600
rect 299308 185542 303771 185544
rect 299308 185540 299314 185542
rect 303705 185539 303771 185542
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110666 480 110756
rect -960 110606 6930 110666
rect -960 110516 480 110606
rect 6870 110530 6930 110606
rect 19558 110530 19564 110532
rect 6870 110470 19564 110530
rect 19558 110468 19564 110470
rect 19628 110468 19634 110532
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3601 84690 3667 84693
rect -960 84688 3667 84690
rect -960 84632 3606 84688
rect 3662 84632 3667 84688
rect -960 84630 3667 84632
rect -960 84540 480 84630
rect 3601 84627 3667 84630
rect 19926 80140 19932 80204
rect 19996 80202 20002 80204
rect 23606 80202 23612 80204
rect 19996 80142 23612 80202
rect 19996 80140 20002 80142
rect 23606 80140 23612 80142
rect 23676 80140 23682 80204
rect 300710 80140 300716 80204
rect 300780 80202 300786 80204
rect 303654 80202 303660 80204
rect 300780 80142 303660 80202
rect 300780 80140 300786 80142
rect 303654 80140 303660 80142
rect 303724 80140 303730 80204
rect 299238 79868 299244 79932
rect 299308 79930 299314 79932
rect 302325 79930 302391 79933
rect 299308 79928 302391 79930
rect 299308 79872 302330 79928
rect 302386 79872 302391 79928
rect 299308 79870 302391 79872
rect 299308 79868 299314 79870
rect 302325 79867 302391 79870
rect 287697 79386 287763 79389
rect 291561 79386 291627 79389
rect 287697 79384 291627 79386
rect 287697 79328 287702 79384
rect 287758 79328 291566 79384
rect 291622 79328 291627 79384
rect 287697 79326 291627 79328
rect 287697 79323 287763 79326
rect 291561 79323 291627 79326
rect 247033 78026 247099 78029
rect 291694 78026 291700 78028
rect 247033 78024 291700 78026
rect 247033 77968 247038 78024
rect 247094 77968 291700 78024
rect 247033 77966 291700 77968
rect 247033 77963 247099 77966
rect 291694 77964 291700 77966
rect 291764 77964 291770 78028
rect 235257 77890 235323 77893
rect 287278 77890 287284 77892
rect 235257 77888 287284 77890
rect 235257 77832 235262 77888
rect 235318 77832 287284 77888
rect 235257 77830 287284 77832
rect 235257 77827 235323 77830
rect 287278 77828 287284 77830
rect 287348 77828 287354 77892
rect 389173 76666 389239 76669
rect 570086 76666 570092 76668
rect 389173 76664 570092 76666
rect 389173 76608 389178 76664
rect 389234 76608 570092 76664
rect 389173 76606 570092 76608
rect 389173 76603 389239 76606
rect 570086 76604 570092 76606
rect 570156 76604 570162 76668
rect 263593 76530 263659 76533
rect 299974 76530 299980 76532
rect 263593 76528 299980 76530
rect 263593 76472 263598 76528
rect 263654 76472 299980 76528
rect 263593 76470 299980 76472
rect 263593 76467 263659 76470
rect 299974 76468 299980 76470
rect 300044 76468 300050 76532
rect 374177 76530 374243 76533
rect 571374 76530 571380 76532
rect 374177 76528 571380 76530
rect 374177 76472 374182 76528
rect 374238 76472 571380 76528
rect 374177 76470 571380 76472
rect 374177 76467 374243 76470
rect 571374 76468 571380 76470
rect 571444 76468 571450 76532
rect 304533 75986 304599 75989
rect 570454 75986 570460 75988
rect 304533 75984 570460 75986
rect 304533 75928 304538 75984
rect 304594 75928 570460 75984
rect 304533 75926 570460 75928
rect 304533 75923 304599 75926
rect 570454 75924 570460 75926
rect 570524 75924 570530 75988
rect 21950 75788 21956 75852
rect 22020 75850 22026 75852
rect 59261 75850 59327 75853
rect 22020 75848 59327 75850
rect 22020 75792 59266 75848
rect 59322 75792 59327 75848
rect 22020 75790 59327 75792
rect 22020 75788 22026 75790
rect 59261 75787 59327 75790
rect 518985 75850 519051 75853
rect 565854 75850 565860 75852
rect 518985 75848 565860 75850
rect 518985 75792 518990 75848
rect 519046 75792 565860 75848
rect 518985 75790 565860 75792
rect 518985 75787 519051 75790
rect 565854 75788 565860 75790
rect 565924 75788 565930 75852
rect 23606 74428 23612 74492
rect 23676 74490 23682 74492
rect 157977 74490 158043 74493
rect 23676 74488 158043 74490
rect 23676 74432 157982 74488
rect 158038 74432 158043 74488
rect 23676 74430 158043 74432
rect 23676 74428 23682 74430
rect 157977 74427 158043 74430
rect 507117 74490 507183 74493
rect 566958 74490 566964 74492
rect 507117 74488 566964 74490
rect 507117 74432 507122 74488
rect 507178 74432 566964 74488
rect 507117 74430 566964 74432
rect 507117 74427 507183 74430
rect 566958 74428 566964 74430
rect 567028 74428 567034 74492
rect 23238 74292 23244 74356
rect 23308 74354 23314 74356
rect 71037 74354 71103 74357
rect 23308 74352 71103 74354
rect 23308 74296 71042 74352
rect 71098 74296 71103 74352
rect 23308 74294 71103 74296
rect 23308 74292 23314 74294
rect 71037 74291 71103 74294
rect 583520 72844 584960 73084
rect -960 71634 480 71724
rect 3049 71634 3115 71637
rect -960 71632 3115 71634
rect -960 71576 3054 71632
rect 3110 71576 3115 71632
rect -960 71574 3115 71576
rect -960 71484 480 71574
rect 3049 71571 3115 71574
rect 298870 66812 298876 66876
rect 298940 66874 298946 66876
rect 335353 66874 335419 66877
rect 336641 66874 336707 66877
rect 298940 66872 336707 66874
rect 298940 66816 335358 66872
rect 335414 66816 336646 66872
rect 336702 66816 336707 66872
rect 298940 66814 336707 66816
rect 298940 66812 298946 66814
rect 335353 66811 335419 66814
rect 336641 66811 336707 66814
rect 57605 61706 57671 61709
rect 57605 61704 60106 61706
rect 57605 61648 57610 61704
rect 57666 61648 60106 61704
rect 57605 61646 60106 61648
rect 57605 61643 57671 61646
rect 60046 61064 60106 61646
rect 218053 61434 218119 61437
rect 303654 61434 303660 61436
rect 218053 61432 303660 61434
rect 218053 61376 218058 61432
rect 218114 61376 303660 61432
rect 218053 61374 303660 61376
rect 218053 61371 218119 61374
rect 303654 61372 303660 61374
rect 303724 61434 303730 61436
rect 303797 61434 303863 61437
rect 303724 61432 303863 61434
rect 303724 61376 303802 61432
rect 303858 61376 303863 61432
rect 303724 61374 303863 61376
rect 303724 61372 303730 61374
rect 303797 61371 303863 61374
rect 99790 60754 99850 61336
rect 102777 60754 102843 60757
rect 99790 60752 102843 60754
rect 99790 60696 102782 60752
rect 102838 60696 102843 60752
rect 99790 60694 102843 60696
rect 102777 60691 102843 60694
rect 99790 59666 99850 60248
rect 244273 60210 244339 60213
rect 291142 60210 291148 60212
rect 244273 60208 291148 60210
rect 244273 60152 244278 60208
rect 244334 60152 291148 60208
rect 244273 60150 291148 60152
rect 244273 60147 244339 60150
rect 291142 60148 291148 60150
rect 291212 60148 291218 60212
rect 240777 60074 240843 60077
rect 287094 60074 287100 60076
rect 240777 60072 287100 60074
rect 240777 60016 240782 60072
rect 240838 60016 287100 60072
rect 240777 60014 287100 60016
rect 240777 60011 240843 60014
rect 287094 60012 287100 60014
rect 287164 60012 287170 60076
rect 245745 59938 245811 59941
rect 292614 59938 292620 59940
rect 245745 59936 292620 59938
rect 245745 59880 245750 59936
rect 245806 59880 292620 59936
rect 245745 59878 292620 59880
rect 245745 59875 245811 59878
rect 292614 59876 292620 59878
rect 292684 59876 292690 59940
rect 102869 59666 102935 59669
rect 99790 59664 102935 59666
rect 99790 59608 102874 59664
rect 102930 59608 102935 59664
rect 99790 59606 102935 59608
rect 102869 59603 102935 59606
rect 583520 59516 584960 59756
rect 303470 59196 303476 59260
rect 303540 59258 303546 59260
rect 321921 59258 321987 59261
rect 303540 59256 321987 59258
rect 303540 59200 321926 59256
rect 321982 59200 321987 59256
rect 303540 59198 321987 59200
rect 303540 59196 303546 59198
rect 321921 59195 321987 59198
rect -960 58428 480 58668
rect 99790 58578 99850 59160
rect 102961 58578 103027 58581
rect 99790 58576 103027 58578
rect 99790 58520 102966 58576
rect 103022 58520 103027 58576
rect 99790 58518 103027 58520
rect 102961 58515 103027 58518
rect 301998 58516 302004 58580
rect 302068 58578 302074 58580
rect 327073 58578 327139 58581
rect 328361 58578 328427 58581
rect 302068 58576 328427 58578
rect 302068 58520 327078 58576
rect 327134 58520 328366 58576
rect 328422 58520 328427 58576
rect 302068 58518 328427 58520
rect 302068 58516 302074 58518
rect 327073 58515 327139 58518
rect 328361 58515 328427 58518
rect 99790 58034 99850 58072
rect 102133 58034 102199 58037
rect 99790 58032 102199 58034
rect 99790 57976 102138 58032
rect 102194 57976 102199 58032
rect 99790 57974 102199 57976
rect 102133 57971 102199 57974
rect 262673 57490 262739 57493
rect 288382 57490 288388 57492
rect 262673 57488 288388 57490
rect 262673 57432 262678 57488
rect 262734 57432 288388 57488
rect 262673 57430 288388 57432
rect 262673 57427 262739 57430
rect 288382 57428 288388 57430
rect 288452 57428 288458 57492
rect 261017 57354 261083 57357
rect 289854 57354 289860 57356
rect 261017 57352 289860 57354
rect 261017 57296 261022 57352
rect 261078 57296 289860 57352
rect 261017 57294 289860 57296
rect 261017 57291 261083 57294
rect 289854 57292 289860 57294
rect 289924 57292 289930 57356
rect 297357 57354 297423 57357
rect 386873 57354 386939 57357
rect 297357 57352 386939 57354
rect 297357 57296 297362 57352
rect 297418 57296 386878 57352
rect 386934 57296 386939 57352
rect 297357 57294 386939 57296
rect 297357 57291 297423 57294
rect 386873 57291 386939 57294
rect 249425 57218 249491 57221
rect 286174 57218 286180 57220
rect 249425 57216 286180 57218
rect 249425 57160 249430 57216
rect 249486 57160 286180 57216
rect 249425 57158 286180 57160
rect 249425 57155 249491 57158
rect 286174 57156 286180 57158
rect 286244 57156 286250 57220
rect 297214 57156 297220 57220
rect 297284 57218 297290 57220
rect 388529 57218 388595 57221
rect 297284 57216 388595 57218
rect 297284 57160 388534 57216
rect 388590 57160 388595 57216
rect 297284 57158 388595 57160
rect 297284 57156 297290 57158
rect 388529 57155 388595 57158
rect 99790 56674 99850 56984
rect 102593 56674 102659 56677
rect 99790 56672 102659 56674
rect 99790 56616 102598 56672
rect 102654 56616 102659 56672
rect 99790 56614 102659 56616
rect 102593 56611 102659 56614
rect 57513 56402 57579 56405
rect 57513 56400 60106 56402
rect 57513 56344 57518 56400
rect 57574 56344 60106 56400
rect 57513 56342 60106 56344
rect 57513 56339 57579 56342
rect 60046 56168 60106 56342
rect 99790 55586 99850 55896
rect 103053 55586 103119 55589
rect 99790 55584 103119 55586
rect 99790 55528 103058 55584
rect 103114 55528 103119 55584
rect 99790 55526 103119 55528
rect 103053 55523 103119 55526
rect 99790 54362 99850 54808
rect 295926 54436 295932 54500
rect 295996 54498 296002 54500
rect 400213 54498 400279 54501
rect 295996 54496 400279 54498
rect 295996 54440 400218 54496
rect 400274 54440 400279 54496
rect 295996 54438 400279 54440
rect 295996 54436 296002 54438
rect 400213 54435 400279 54438
rect 102133 54362 102199 54365
rect 99790 54360 102199 54362
rect 99790 54304 102138 54360
rect 102194 54304 102199 54360
rect 99790 54302 102199 54304
rect 102133 54299 102199 54302
rect 99790 53546 99850 53720
rect 102133 53546 102199 53549
rect 99790 53544 102199 53546
rect 99790 53488 102138 53544
rect 102194 53488 102199 53544
rect 99790 53486 102199 53488
rect 102133 53483 102199 53486
rect 99790 52594 99850 52632
rect 102133 52594 102199 52597
rect 99790 52592 102199 52594
rect 99790 52536 102138 52592
rect 102194 52536 102199 52592
rect 99790 52534 102199 52536
rect 102133 52531 102199 52534
rect 195973 52322 196039 52325
rect 195973 52320 199394 52322
rect 195973 52264 195978 52320
rect 196034 52264 199394 52320
rect 195973 52262 199394 52264
rect 195973 52259 196039 52262
rect 199334 52088 199394 52262
rect 57053 51778 57119 51781
rect 196065 51778 196131 51781
rect 57053 51776 60106 51778
rect 57053 51720 57058 51776
rect 57114 51720 60106 51776
rect 57053 51718 60106 51720
rect 57053 51715 57119 51718
rect 60046 51272 60106 51718
rect 196065 51776 199394 51778
rect 196065 51720 196070 51776
rect 196126 51720 199394 51776
rect 196065 51718 199394 51720
rect 196065 51715 196131 51718
rect 99790 51098 99850 51544
rect 199334 51272 199394 51718
rect 103237 51098 103303 51101
rect 99790 51096 103303 51098
rect 99790 51040 103242 51096
rect 103298 51040 103303 51096
rect 99790 51038 103303 51040
rect 103237 51035 103303 51038
rect 195973 50962 196039 50965
rect 195973 50960 199394 50962
rect 195973 50904 195978 50960
rect 196034 50904 199394 50960
rect 195973 50902 199394 50904
rect 195973 50899 196039 50902
rect 199334 50456 199394 50902
rect 99790 50146 99850 50456
rect 102133 50146 102199 50149
rect 99790 50144 102199 50146
rect 99790 50088 102138 50144
rect 102194 50088 102199 50144
rect 99790 50086 102199 50088
rect 102133 50083 102199 50086
rect 195973 49602 196039 49605
rect 199334 49602 199394 49640
rect 195973 49600 199394 49602
rect 195973 49544 195978 49600
rect 196034 49544 199394 49600
rect 195973 49542 199394 49544
rect 195973 49539 196039 49542
rect 196065 49466 196131 49469
rect 196065 49464 199394 49466
rect 196065 49408 196070 49464
rect 196126 49408 199394 49464
rect 196065 49406 199394 49408
rect 196065 49403 196131 49406
rect 99790 49194 99850 49368
rect 102133 49194 102199 49197
rect 99790 49192 102199 49194
rect 99790 49136 102138 49192
rect 102194 49136 102199 49192
rect 99790 49134 102199 49136
rect 102133 49131 102199 49134
rect 199334 48824 199394 49406
rect 99790 47698 99850 48280
rect 195973 48242 196039 48245
rect 195973 48240 199394 48242
rect 195973 48184 195978 48240
rect 196034 48184 199394 48240
rect 195973 48182 199394 48184
rect 195973 48179 196039 48182
rect 199334 48008 199394 48182
rect 102961 47698 103027 47701
rect 99790 47696 103027 47698
rect 99790 47640 102966 47696
rect 103022 47640 103027 47696
rect 99790 47638 103027 47640
rect 102961 47635 103027 47638
rect 196065 47698 196131 47701
rect 196065 47696 199394 47698
rect 196065 47640 196070 47696
rect 196126 47640 199394 47696
rect 196065 47638 199394 47640
rect 196065 47635 196131 47638
rect 199334 47192 199394 47638
rect 99790 47018 99850 47192
rect 102593 47018 102659 47021
rect 99790 47016 102659 47018
rect 99790 46960 102598 47016
rect 102654 46960 102659 47016
rect 99790 46958 102659 46960
rect 102593 46955 102659 46958
rect 57513 46882 57579 46885
rect 195973 46882 196039 46885
rect 57513 46880 60106 46882
rect 57513 46824 57518 46880
rect 57574 46824 60106 46880
rect 57513 46822 60106 46824
rect 57513 46819 57579 46822
rect 60046 46376 60106 46822
rect 195973 46880 199394 46882
rect 195973 46824 195978 46880
rect 196034 46824 199394 46880
rect 195973 46822 199394 46824
rect 195973 46819 196039 46822
rect 199334 46376 199394 46822
rect 196157 46202 196223 46205
rect 196157 46200 199394 46202
rect 196157 46144 196162 46200
rect 196218 46144 199394 46200
rect 583520 46188 584960 46428
rect 196157 46142 199394 46144
rect 196157 46139 196223 46142
rect 99790 45794 99850 46104
rect 102869 45794 102935 45797
rect 99790 45792 102935 45794
rect 99790 45736 102874 45792
rect 102930 45736 102935 45792
rect 99790 45734 102935 45736
rect 102869 45731 102935 45734
rect -960 45522 480 45612
rect 199334 45560 199394 46142
rect 3325 45522 3391 45525
rect -960 45520 3391 45522
rect -960 45464 3330 45520
rect 3386 45464 3391 45520
rect -960 45462 3391 45464
rect -960 45372 480 45462
rect 3325 45459 3391 45462
rect 195973 45250 196039 45253
rect 195973 45248 199394 45250
rect 195973 45192 195978 45248
rect 196034 45192 199394 45248
rect 195973 45190 199394 45192
rect 195973 45187 196039 45190
rect 99790 44434 99850 45016
rect 199334 44744 199394 45190
rect 103421 44434 103487 44437
rect 99790 44432 103487 44434
rect 99790 44376 103426 44432
rect 103482 44376 103487 44432
rect 99790 44374 103487 44376
rect 103421 44371 103487 44374
rect 196065 44162 196131 44165
rect 196065 44160 199394 44162
rect 196065 44104 196070 44160
rect 196126 44104 199394 44160
rect 196065 44102 199394 44104
rect 196065 44099 196131 44102
rect 199334 43928 199394 44102
rect 99790 43346 99850 43928
rect 195973 43754 196039 43757
rect 195973 43752 199394 43754
rect 195973 43696 195978 43752
rect 196034 43696 199394 43752
rect 195973 43694 199394 43696
rect 195973 43691 196039 43694
rect 102317 43346 102383 43349
rect 99790 43344 102383 43346
rect 99790 43288 102322 43344
rect 102378 43288 102383 43344
rect 99790 43286 102383 43288
rect 102317 43283 102383 43286
rect 199334 43112 199394 43694
rect 102133 42938 102199 42941
rect 99790 42936 102199 42938
rect 99790 42880 102138 42936
rect 102194 42880 102199 42936
rect 99790 42878 102199 42880
rect 99790 42840 99850 42878
rect 102133 42875 102199 42878
rect 195973 42530 196039 42533
rect 195973 42528 199394 42530
rect 195973 42472 195978 42528
rect 196034 42472 199394 42528
rect 195973 42470 199394 42472
rect 195973 42467 196039 42470
rect 199334 42296 199394 42470
rect 57145 42122 57211 42125
rect 196065 42122 196131 42125
rect 57145 42120 60106 42122
rect 57145 42064 57150 42120
rect 57206 42064 60106 42120
rect 57145 42062 60106 42064
rect 57145 42059 57211 42062
rect 60046 41480 60106 42062
rect 196065 42120 199394 42122
rect 196065 42064 196070 42120
rect 196126 42064 199394 42120
rect 196065 42062 199394 42064
rect 196065 42059 196131 42062
rect 99790 41442 99850 41752
rect 199334 41480 199394 42062
rect 102225 41442 102291 41445
rect 99790 41440 102291 41442
rect 99790 41384 102230 41440
rect 102286 41384 102291 41440
rect 99790 41382 102291 41384
rect 102225 41379 102291 41382
rect 195973 41170 196039 41173
rect 195973 41168 199394 41170
rect 195973 41112 195978 41168
rect 196034 41112 199394 41168
rect 195973 41110 199394 41112
rect 195973 41107 196039 41110
rect 199334 40664 199394 41110
rect 99790 40082 99850 40664
rect 102133 40082 102199 40085
rect 99790 40080 102199 40082
rect 99790 40024 102138 40080
rect 102194 40024 102199 40080
rect 99790 40022 102199 40024
rect 102133 40019 102199 40022
rect 195973 39946 196039 39949
rect 195973 39944 199394 39946
rect 195973 39888 195978 39944
rect 196034 39888 199394 39944
rect 195973 39886 199394 39888
rect 195973 39883 196039 39886
rect 199334 39848 199394 39886
rect 99790 38994 99850 39576
rect 196065 39538 196131 39541
rect 196065 39536 199394 39538
rect 196065 39480 196070 39536
rect 196126 39480 199394 39536
rect 196065 39478 199394 39480
rect 196065 39475 196131 39478
rect 199334 39032 199394 39478
rect 102777 38994 102843 38997
rect 99790 38992 102843 38994
rect 99790 38936 102782 38992
rect 102838 38936 102843 38992
rect 99790 38934 102843 38936
rect 102777 38931 102843 38934
rect 196157 38586 196223 38589
rect 196157 38584 199394 38586
rect 196157 38528 196162 38584
rect 196218 38528 199394 38584
rect 196157 38526 199394 38528
rect 196157 38523 196223 38526
rect 99790 37906 99850 38488
rect 199334 38216 199394 38526
rect 195973 38042 196039 38045
rect 195973 38040 199394 38042
rect 195973 37984 195978 38040
rect 196034 37984 199394 38040
rect 195973 37982 199394 37984
rect 195973 37979 196039 37982
rect 102685 37906 102751 37909
rect 99790 37904 102751 37906
rect 99790 37848 102690 37904
rect 102746 37848 102751 37904
rect 99790 37846 102751 37848
rect 102685 37843 102751 37846
rect 199334 37400 199394 37982
rect 99790 37362 99850 37400
rect 102869 37362 102935 37365
rect 99790 37360 102935 37362
rect 99790 37304 102874 37360
rect 102930 37304 102935 37360
rect 99790 37302 102935 37304
rect 102869 37299 102935 37302
rect 195973 37090 196039 37093
rect 195973 37088 199394 37090
rect 195973 37032 195978 37088
rect 196034 37032 199394 37088
rect 195973 37030 199394 37032
rect 195973 37027 196039 37030
rect 57053 36954 57119 36957
rect 57053 36952 60106 36954
rect 57053 36896 57058 36952
rect 57114 36896 60106 36952
rect 57053 36894 60106 36896
rect 57053 36891 57119 36894
rect 60046 36584 60106 36894
rect 199334 36584 199394 37030
rect 99790 36138 99850 36312
rect 102593 36138 102659 36141
rect 99790 36136 102659 36138
rect 99790 36080 102598 36136
rect 102654 36080 102659 36136
rect 99790 36078 102659 36080
rect 102593 36075 102659 36078
rect 195973 35866 196039 35869
rect 195973 35864 199394 35866
rect 195973 35808 195978 35864
rect 196034 35808 199394 35864
rect 195973 35806 199394 35808
rect 195973 35803 196039 35806
rect 199334 35768 199394 35806
rect 196065 35458 196131 35461
rect 196065 35456 199394 35458
rect 196065 35400 196070 35456
rect 196126 35400 199394 35456
rect 196065 35398 199394 35400
rect 196065 35395 196131 35398
rect 99790 34642 99850 35224
rect 199334 34952 199394 35398
rect 102133 34642 102199 34645
rect 99790 34640 102199 34642
rect 99790 34584 102138 34640
rect 102194 34584 102199 34640
rect 99790 34582 102199 34584
rect 102133 34579 102199 34582
rect 195973 34370 196039 34373
rect 195973 34368 199394 34370
rect 195973 34312 195978 34368
rect 196034 34312 199394 34368
rect 195973 34310 199394 34312
rect 195973 34307 196039 34310
rect 199334 34136 199394 34310
rect 99790 33554 99850 34136
rect 196065 33826 196131 33829
rect 196065 33824 199394 33826
rect 196065 33768 196070 33824
rect 196126 33768 199394 33824
rect 196065 33766 199394 33768
rect 196065 33763 196131 33766
rect 102317 33554 102383 33557
rect 99790 33552 102383 33554
rect 99790 33496 102322 33552
rect 102378 33496 102383 33552
rect 99790 33494 102383 33496
rect 102317 33491 102383 33494
rect 199334 33320 199394 33766
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect 99790 32466 99850 33048
rect 195973 33010 196039 33013
rect 195973 33008 199394 33010
rect 195973 32952 195978 33008
rect 196034 32952 199394 33008
rect 583520 32996 584960 33236
rect 195973 32950 199394 32952
rect 195973 32947 196039 32950
rect 199334 32504 199394 32950
rect 102133 32466 102199 32469
rect 99790 32464 102199 32466
rect 99790 32408 102138 32464
rect 102194 32408 102199 32464
rect 99790 32406 102199 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 102133 32403 102199 32406
rect 99790 31786 99850 31960
rect 102225 31786 102291 31789
rect 99790 31784 102291 31786
rect 99790 31728 102230 31784
rect 102286 31728 102291 31784
rect 99790 31726 102291 31728
rect 102225 31723 102291 31726
rect 57605 31650 57671 31653
rect 60046 31650 60106 31688
rect 57605 31648 60106 31650
rect 57605 31592 57610 31648
rect 57666 31592 60106 31648
rect 57605 31590 60106 31592
rect 195973 31650 196039 31653
rect 199334 31650 199394 31688
rect 195973 31648 199394 31650
rect 195973 31592 195978 31648
rect 196034 31592 199394 31648
rect 195973 31590 199394 31592
rect 57605 31587 57671 31590
rect 195973 31587 196039 31590
rect 196065 31242 196131 31245
rect 196065 31240 199394 31242
rect 196065 31184 196070 31240
rect 196126 31184 199394 31240
rect 196065 31182 199394 31184
rect 196065 31179 196131 31182
rect 199334 30872 199394 31182
rect 99790 30562 99850 30872
rect 102133 30562 102199 30565
rect 99790 30560 102199 30562
rect 99790 30504 102138 30560
rect 102194 30504 102199 30560
rect 99790 30502 102199 30504
rect 102133 30499 102199 30502
rect 195973 30290 196039 30293
rect 195973 30288 199394 30290
rect 195973 30232 195978 30288
rect 196034 30232 199394 30288
rect 195973 30230 199394 30232
rect 195973 30227 196039 30230
rect 199334 30056 199394 30230
rect 99790 29338 99850 29784
rect 196065 29746 196131 29749
rect 196065 29744 199394 29746
rect 196065 29688 196070 29744
rect 196126 29688 199394 29744
rect 196065 29686 199394 29688
rect 196065 29683 196131 29686
rect 102133 29338 102199 29341
rect 99790 29336 102199 29338
rect 99790 29280 102138 29336
rect 102194 29280 102199 29336
rect 99790 29278 102199 29280
rect 102133 29275 102199 29278
rect 199334 29240 199394 29686
rect 195973 28930 196039 28933
rect 195973 28928 199394 28930
rect 195973 28872 195978 28928
rect 196034 28872 199394 28928
rect 195973 28870 199394 28872
rect 195973 28867 196039 28870
rect 99790 28522 99850 28696
rect 102133 28522 102199 28525
rect 99790 28520 102199 28522
rect 99790 28464 102138 28520
rect 102194 28464 102199 28520
rect 99790 28462 102199 28464
rect 102133 28459 102199 28462
rect 199334 28424 199394 28870
rect 195973 28114 196039 28117
rect 195973 28112 199394 28114
rect 195973 28056 195978 28112
rect 196034 28056 199394 28112
rect 195973 28054 199394 28056
rect 195973 28051 196039 28054
rect 102133 27706 102199 27709
rect 99790 27704 102199 27706
rect 99790 27648 102138 27704
rect 102194 27648 102199 27704
rect 99790 27646 102199 27648
rect 99790 27608 99850 27646
rect 102133 27643 102199 27646
rect 199334 27608 199394 28054
rect 195973 27298 196039 27301
rect 195973 27296 199394 27298
rect 195973 27240 195978 27296
rect 196034 27240 199394 27296
rect 195973 27238 199394 27240
rect 195973 27235 196039 27238
rect 57237 27162 57303 27165
rect 57237 27160 60106 27162
rect 57237 27104 57242 27160
rect 57298 27104 60106 27160
rect 57237 27102 60106 27104
rect 57237 27099 57303 27102
rect 60046 26792 60106 27102
rect 199334 26792 199394 27238
rect 99790 26346 99850 26520
rect 102777 26346 102843 26349
rect 99790 26344 102843 26346
rect 99790 26288 102782 26344
rect 102838 26288 102843 26344
rect 99790 26286 102843 26288
rect 102777 26283 102843 26286
rect 195973 26210 196039 26213
rect 195973 26208 199394 26210
rect 195973 26152 195978 26208
rect 196034 26152 199394 26208
rect 195973 26150 199394 26152
rect 195973 26147 196039 26150
rect 199334 25976 199394 26150
rect 389633 22130 389699 22133
rect 569534 22130 569540 22132
rect 389633 22128 569540 22130
rect 389633 22072 389638 22128
rect 389694 22072 569540 22128
rect 389633 22070 569540 22072
rect 389633 22067 389699 22070
rect 569534 22068 569540 22070
rect 569604 22068 569610 22132
rect 18454 21932 18460 21996
rect 18524 21994 18530 21996
rect 368105 21994 368171 21997
rect 18524 21992 368171 21994
rect 18524 21936 368110 21992
rect 368166 21936 368171 21992
rect 18524 21934 368171 21936
rect 18524 21932 18530 21934
rect 368105 21931 368171 21934
rect 19558 21796 19564 21860
rect 19628 21858 19634 21860
rect 342989 21858 343055 21861
rect 19628 21856 343055 21858
rect 19628 21800 342994 21856
rect 343050 21800 343055 21856
rect 19628 21798 343055 21800
rect 19628 21796 19634 21798
rect 342989 21795 343055 21798
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 295932 700300 295996 700364
rect 569540 590956 569604 591020
rect 292620 586392 292684 586396
rect 292620 586336 292634 586392
rect 292634 586336 292684 586392
rect 292620 586332 292684 586336
rect 285628 585924 285692 585988
rect 303476 585924 303540 585988
rect 23244 585788 23308 585852
rect 287100 585788 287164 585852
rect 299980 585788 300044 585852
rect 570092 585788 570156 585852
rect 21956 585652 22020 585716
rect 288388 585652 288452 585716
rect 291700 585652 291764 585716
rect 565860 585652 565924 585716
rect 302004 583068 302068 583132
rect 298692 582932 298756 582996
rect 568620 580212 568684 580276
rect 297220 571916 297284 571980
rect 567884 571916 567948 571980
rect 18460 502420 18524 502484
rect 568620 463524 568684 463588
rect 302004 461212 302068 461276
rect 287100 460940 287164 461004
rect 303476 461000 303540 461004
rect 567700 461136 567764 461140
rect 567700 461080 567750 461136
rect 567750 461080 567764 461136
rect 567700 461076 567764 461080
rect 303476 460944 303526 461000
rect 303526 460944 303540 461000
rect 303476 460940 303540 460944
rect 21956 459444 22020 459508
rect 567884 459368 567948 459372
rect 567884 459312 567934 459368
rect 567934 459312 567948 459368
rect 567884 459308 567948 459312
rect 298692 459172 298756 459236
rect 291148 458900 291212 458964
rect 289860 458764 289924 458828
rect 571380 458764 571444 458828
rect 298692 458220 298756 458284
rect 23244 458084 23308 458148
rect 285628 458084 285692 458148
rect 566412 458084 566476 458148
rect 287652 457872 287716 457876
rect 287652 457816 287666 457872
rect 287666 457816 287716 457872
rect 287652 457812 287716 457816
rect 286180 444892 286244 444956
rect 570460 418236 570524 418300
rect 568436 336636 568500 336700
rect 21220 332828 21284 332892
rect 300900 332556 300964 332620
rect 288204 332420 288268 332484
rect 565860 332344 565924 332348
rect 565860 332288 565874 332344
rect 565874 332288 565924 332344
rect 565860 332284 565924 332288
rect 22692 332148 22756 332212
rect 302740 332148 302804 332212
rect 285628 331392 285692 331396
rect 285628 331336 285642 331392
rect 285642 331336 285692 331392
rect 285628 331332 285692 331336
rect 298692 317520 298756 317524
rect 298692 317464 298742 317520
rect 298742 317464 298756 317520
rect 298692 317460 298756 317464
rect 302004 315752 302068 315756
rect 302004 315696 302054 315752
rect 302054 315696 302068 315752
rect 302004 315692 302068 315696
rect 567700 315692 567764 315756
rect 302004 314740 302068 314804
rect 568436 314664 568500 314668
rect 568436 314608 568486 314664
rect 568486 314608 568500 314664
rect 568436 314604 568500 314608
rect 21404 207708 21468 207772
rect 22140 207572 22204 207636
rect 22140 206348 22204 206412
rect 21404 206212 21468 206276
rect 300900 204716 300964 204780
rect 302004 204776 302068 204780
rect 302004 204720 302054 204776
rect 302054 204720 302068 204776
rect 302004 204716 302068 204720
rect 567332 204368 567396 204372
rect 567332 204312 567346 204368
rect 567346 204312 567396 204368
rect 567332 204308 567396 204312
rect 21956 203764 22020 203828
rect 287100 203492 287164 203556
rect 21220 202812 21284 202876
rect 22692 202812 22756 202876
rect 287284 202872 287348 202876
rect 287284 202816 287334 202872
rect 287334 202816 287348 202872
rect 287284 202812 287348 202816
rect 288204 202812 288268 202876
rect 302740 201316 302804 201380
rect 19932 199956 19996 200020
rect 298692 188940 298756 189004
rect 298876 188804 298940 188868
rect 565860 187580 565924 187644
rect 301452 186356 301516 186420
rect 299244 185540 299308 185604
rect 19564 110468 19628 110532
rect 19932 80140 19996 80204
rect 23612 80140 23676 80204
rect 300716 80140 300780 80204
rect 303660 80140 303724 80204
rect 299244 79868 299308 79932
rect 291700 77964 291764 78028
rect 287284 77828 287348 77892
rect 570092 76604 570156 76668
rect 299980 76468 300044 76532
rect 571380 76468 571444 76532
rect 570460 75924 570524 75988
rect 21956 75788 22020 75852
rect 565860 75788 565924 75852
rect 23612 74428 23676 74492
rect 566964 74428 567028 74492
rect 23244 74292 23308 74356
rect 298876 66812 298940 66876
rect 303660 61372 303724 61436
rect 291148 60148 291212 60212
rect 287100 60012 287164 60076
rect 292620 59876 292684 59940
rect 303476 59196 303540 59260
rect 302004 58516 302068 58580
rect 288388 57428 288452 57492
rect 289860 57292 289924 57356
rect 286180 57156 286244 57220
rect 297220 57156 297284 57220
rect 295932 54436 295996 54500
rect 569540 22068 569604 22132
rect 18460 21932 18524 21996
rect 19564 21796 19628 21860
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 700000 51914 700398
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 700000 87914 700398
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 700000 123914 700398
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 700000 159914 700398
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 700000 195914 700398
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 700000 231914 700398
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 700000 267914 700398
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 33868 691954 34868 691986
rect 33868 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 34868 691954
rect 33868 691634 34868 691718
rect 33868 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 34868 691634
rect 33868 691366 34868 691398
rect 53868 691954 54868 691986
rect 53868 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 54868 691954
rect 53868 691634 54868 691718
rect 53868 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 54868 691634
rect 53868 691366 54868 691398
rect 73868 691954 74868 691986
rect 73868 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 74868 691954
rect 73868 691634 74868 691718
rect 73868 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 74868 691634
rect 73868 691366 74868 691398
rect 93868 691954 94868 691986
rect 93868 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 94868 691954
rect 93868 691634 94868 691718
rect 93868 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 94868 691634
rect 93868 691366 94868 691398
rect 113868 691954 114868 691986
rect 113868 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 114868 691954
rect 113868 691634 114868 691718
rect 113868 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 114868 691634
rect 113868 691366 114868 691398
rect 133868 691954 134868 691986
rect 133868 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 134868 691954
rect 133868 691634 134868 691718
rect 133868 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 134868 691634
rect 133868 691366 134868 691398
rect 153868 691954 154868 691986
rect 153868 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 154868 691954
rect 153868 691634 154868 691718
rect 153868 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 154868 691634
rect 153868 691366 154868 691398
rect 173868 691954 174868 691986
rect 173868 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 174868 691954
rect 173868 691634 174868 691718
rect 173868 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 174868 691634
rect 173868 691366 174868 691398
rect 193868 691954 194868 691986
rect 193868 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 194868 691954
rect 193868 691634 194868 691718
rect 193868 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 194868 691634
rect 193868 691366 194868 691398
rect 213868 691954 214868 691986
rect 213868 691718 213930 691954
rect 214166 691718 214250 691954
rect 214486 691718 214570 691954
rect 214806 691718 214868 691954
rect 213868 691634 214868 691718
rect 213868 691398 213930 691634
rect 214166 691398 214250 691634
rect 214486 691398 214570 691634
rect 214806 691398 214868 691634
rect 213868 691366 214868 691398
rect 233868 691954 234868 691986
rect 233868 691718 233930 691954
rect 234166 691718 234250 691954
rect 234486 691718 234570 691954
rect 234806 691718 234868 691954
rect 233868 691634 234868 691718
rect 233868 691398 233930 691634
rect 234166 691398 234250 691634
rect 234486 691398 234570 691634
rect 234806 691398 234868 691634
rect 233868 691366 234868 691398
rect 253868 691954 254868 691986
rect 253868 691718 253930 691954
rect 254166 691718 254250 691954
rect 254486 691718 254570 691954
rect 254806 691718 254868 691954
rect 253868 691634 254868 691718
rect 253868 691398 253930 691634
rect 254166 691398 254250 691634
rect 254486 691398 254570 691634
rect 254806 691398 254868 691634
rect 253868 691366 254868 691398
rect 273868 691954 274868 691986
rect 273868 691718 273930 691954
rect 274166 691718 274250 691954
rect 274486 691718 274570 691954
rect 274806 691718 274868 691954
rect 273868 691634 274868 691718
rect 273868 691398 273930 691634
rect 274166 691398 274250 691634
rect 274486 691398 274570 691634
rect 274806 691398 274868 691634
rect 273868 691366 274868 691398
rect 294294 691954 294914 705242
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 295931 700364 295997 700365
rect 295931 700300 295932 700364
rect 295996 700300 295997 700364
rect 295931 700299 295997 700300
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 23868 687454 24868 687486
rect 23868 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 24868 687454
rect 23868 687134 24868 687218
rect 23868 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 24868 687134
rect 23868 686866 24868 686898
rect 43868 687454 44868 687486
rect 43868 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 44868 687454
rect 43868 687134 44868 687218
rect 43868 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 44868 687134
rect 43868 686866 44868 686898
rect 63868 687454 64868 687486
rect 63868 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 64868 687454
rect 63868 687134 64868 687218
rect 63868 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 64868 687134
rect 63868 686866 64868 686898
rect 83868 687454 84868 687486
rect 83868 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 84868 687454
rect 83868 687134 84868 687218
rect 83868 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 84868 687134
rect 83868 686866 84868 686898
rect 103868 687454 104868 687486
rect 103868 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 104868 687454
rect 103868 687134 104868 687218
rect 103868 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 104868 687134
rect 103868 686866 104868 686898
rect 123868 687454 124868 687486
rect 123868 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 124868 687454
rect 123868 687134 124868 687218
rect 123868 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 124868 687134
rect 123868 686866 124868 686898
rect 143868 687454 144868 687486
rect 143868 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 144868 687454
rect 143868 687134 144868 687218
rect 143868 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 144868 687134
rect 143868 686866 144868 686898
rect 163868 687454 164868 687486
rect 163868 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 164868 687454
rect 163868 687134 164868 687218
rect 163868 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 164868 687134
rect 163868 686866 164868 686898
rect 183868 687454 184868 687486
rect 183868 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 184868 687454
rect 183868 687134 184868 687218
rect 183868 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 184868 687134
rect 183868 686866 184868 686898
rect 203868 687454 204868 687486
rect 203868 687218 203930 687454
rect 204166 687218 204250 687454
rect 204486 687218 204570 687454
rect 204806 687218 204868 687454
rect 203868 687134 204868 687218
rect 203868 686898 203930 687134
rect 204166 686898 204250 687134
rect 204486 686898 204570 687134
rect 204806 686898 204868 687134
rect 203868 686866 204868 686898
rect 223868 687454 224868 687486
rect 223868 687218 223930 687454
rect 224166 687218 224250 687454
rect 224486 687218 224570 687454
rect 224806 687218 224868 687454
rect 223868 687134 224868 687218
rect 223868 686898 223930 687134
rect 224166 686898 224250 687134
rect 224486 686898 224570 687134
rect 224806 686898 224868 687134
rect 223868 686866 224868 686898
rect 243868 687454 244868 687486
rect 243868 687218 243930 687454
rect 244166 687218 244250 687454
rect 244486 687218 244570 687454
rect 244806 687218 244868 687454
rect 243868 687134 244868 687218
rect 243868 686898 243930 687134
rect 244166 686898 244250 687134
rect 244486 686898 244570 687134
rect 244806 686898 244868 687134
rect 243868 686866 244868 686898
rect 263868 687454 264868 687486
rect 263868 687218 263930 687454
rect 264166 687218 264250 687454
rect 264486 687218 264570 687454
rect 264806 687218 264868 687454
rect 263868 687134 264868 687218
rect 263868 686898 263930 687134
rect 264166 686898 264250 687134
rect 264486 686898 264570 687134
rect 264806 686898 264868 687134
rect 263868 686866 264868 686898
rect 283868 687454 284868 687486
rect 283868 687218 283930 687454
rect 284166 687218 284250 687454
rect 284486 687218 284570 687454
rect 284806 687218 284868 687454
rect 283868 687134 284868 687218
rect 283868 686898 283930 687134
rect 284166 686898 284250 687134
rect 284486 686898 284570 687134
rect 284806 686898 284868 687134
rect 283868 686866 284868 686898
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 33868 655954 34868 655986
rect 33868 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 34868 655954
rect 33868 655634 34868 655718
rect 33868 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 34868 655634
rect 33868 655366 34868 655398
rect 53868 655954 54868 655986
rect 53868 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 54868 655954
rect 53868 655634 54868 655718
rect 53868 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 54868 655634
rect 53868 655366 54868 655398
rect 73868 655954 74868 655986
rect 73868 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 74868 655954
rect 73868 655634 74868 655718
rect 73868 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 74868 655634
rect 73868 655366 74868 655398
rect 93868 655954 94868 655986
rect 93868 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 94868 655954
rect 93868 655634 94868 655718
rect 93868 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 94868 655634
rect 93868 655366 94868 655398
rect 113868 655954 114868 655986
rect 113868 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 114868 655954
rect 113868 655634 114868 655718
rect 113868 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 114868 655634
rect 113868 655366 114868 655398
rect 133868 655954 134868 655986
rect 133868 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 134868 655954
rect 133868 655634 134868 655718
rect 133868 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 134868 655634
rect 133868 655366 134868 655398
rect 153868 655954 154868 655986
rect 153868 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 154868 655954
rect 153868 655634 154868 655718
rect 153868 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 154868 655634
rect 153868 655366 154868 655398
rect 173868 655954 174868 655986
rect 173868 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 174868 655954
rect 173868 655634 174868 655718
rect 173868 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 174868 655634
rect 173868 655366 174868 655398
rect 193868 655954 194868 655986
rect 193868 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 194868 655954
rect 193868 655634 194868 655718
rect 193868 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 194868 655634
rect 193868 655366 194868 655398
rect 213868 655954 214868 655986
rect 213868 655718 213930 655954
rect 214166 655718 214250 655954
rect 214486 655718 214570 655954
rect 214806 655718 214868 655954
rect 213868 655634 214868 655718
rect 213868 655398 213930 655634
rect 214166 655398 214250 655634
rect 214486 655398 214570 655634
rect 214806 655398 214868 655634
rect 213868 655366 214868 655398
rect 233868 655954 234868 655986
rect 233868 655718 233930 655954
rect 234166 655718 234250 655954
rect 234486 655718 234570 655954
rect 234806 655718 234868 655954
rect 233868 655634 234868 655718
rect 233868 655398 233930 655634
rect 234166 655398 234250 655634
rect 234486 655398 234570 655634
rect 234806 655398 234868 655634
rect 233868 655366 234868 655398
rect 253868 655954 254868 655986
rect 253868 655718 253930 655954
rect 254166 655718 254250 655954
rect 254486 655718 254570 655954
rect 254806 655718 254868 655954
rect 253868 655634 254868 655718
rect 253868 655398 253930 655634
rect 254166 655398 254250 655634
rect 254486 655398 254570 655634
rect 254806 655398 254868 655634
rect 253868 655366 254868 655398
rect 273868 655954 274868 655986
rect 273868 655718 273930 655954
rect 274166 655718 274250 655954
rect 274486 655718 274570 655954
rect 274806 655718 274868 655954
rect 273868 655634 274868 655718
rect 273868 655398 273930 655634
rect 274166 655398 274250 655634
rect 274486 655398 274570 655634
rect 274806 655398 274868 655634
rect 273868 655366 274868 655398
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 23868 651454 24868 651486
rect 23868 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 24868 651454
rect 23868 651134 24868 651218
rect 23868 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 24868 651134
rect 23868 650866 24868 650898
rect 43868 651454 44868 651486
rect 43868 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 44868 651454
rect 43868 651134 44868 651218
rect 43868 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 44868 651134
rect 43868 650866 44868 650898
rect 63868 651454 64868 651486
rect 63868 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 64868 651454
rect 63868 651134 64868 651218
rect 63868 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 64868 651134
rect 63868 650866 64868 650898
rect 83868 651454 84868 651486
rect 83868 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 84868 651454
rect 83868 651134 84868 651218
rect 83868 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 84868 651134
rect 83868 650866 84868 650898
rect 103868 651454 104868 651486
rect 103868 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 104868 651454
rect 103868 651134 104868 651218
rect 103868 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 104868 651134
rect 103868 650866 104868 650898
rect 123868 651454 124868 651486
rect 123868 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 124868 651454
rect 123868 651134 124868 651218
rect 123868 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 124868 651134
rect 123868 650866 124868 650898
rect 143868 651454 144868 651486
rect 143868 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 144868 651454
rect 143868 651134 144868 651218
rect 143868 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 144868 651134
rect 143868 650866 144868 650898
rect 163868 651454 164868 651486
rect 163868 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 164868 651454
rect 163868 651134 164868 651218
rect 163868 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 164868 651134
rect 163868 650866 164868 650898
rect 183868 651454 184868 651486
rect 183868 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 184868 651454
rect 183868 651134 184868 651218
rect 183868 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 184868 651134
rect 183868 650866 184868 650898
rect 203868 651454 204868 651486
rect 203868 651218 203930 651454
rect 204166 651218 204250 651454
rect 204486 651218 204570 651454
rect 204806 651218 204868 651454
rect 203868 651134 204868 651218
rect 203868 650898 203930 651134
rect 204166 650898 204250 651134
rect 204486 650898 204570 651134
rect 204806 650898 204868 651134
rect 203868 650866 204868 650898
rect 223868 651454 224868 651486
rect 223868 651218 223930 651454
rect 224166 651218 224250 651454
rect 224486 651218 224570 651454
rect 224806 651218 224868 651454
rect 223868 651134 224868 651218
rect 223868 650898 223930 651134
rect 224166 650898 224250 651134
rect 224486 650898 224570 651134
rect 224806 650898 224868 651134
rect 223868 650866 224868 650898
rect 243868 651454 244868 651486
rect 243868 651218 243930 651454
rect 244166 651218 244250 651454
rect 244486 651218 244570 651454
rect 244806 651218 244868 651454
rect 243868 651134 244868 651218
rect 243868 650898 243930 651134
rect 244166 650898 244250 651134
rect 244486 650898 244570 651134
rect 244806 650898 244868 651134
rect 243868 650866 244868 650898
rect 263868 651454 264868 651486
rect 263868 651218 263930 651454
rect 264166 651218 264250 651454
rect 264486 651218 264570 651454
rect 264806 651218 264868 651454
rect 263868 651134 264868 651218
rect 263868 650898 263930 651134
rect 264166 650898 264250 651134
rect 264486 650898 264570 651134
rect 264806 650898 264868 651134
rect 263868 650866 264868 650898
rect 283868 651454 284868 651486
rect 283868 651218 283930 651454
rect 284166 651218 284250 651454
rect 284486 651218 284570 651454
rect 284806 651218 284868 651454
rect 283868 651134 284868 651218
rect 283868 650898 283930 651134
rect 284166 650898 284250 651134
rect 284486 650898 284570 651134
rect 284806 650898 284868 651134
rect 283868 650866 284868 650898
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 33868 619954 34868 619986
rect 33868 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 34868 619954
rect 33868 619634 34868 619718
rect 33868 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 34868 619634
rect 33868 619366 34868 619398
rect 53868 619954 54868 619986
rect 53868 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 54868 619954
rect 53868 619634 54868 619718
rect 53868 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 54868 619634
rect 53868 619366 54868 619398
rect 73868 619954 74868 619986
rect 73868 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 74868 619954
rect 73868 619634 74868 619718
rect 73868 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 74868 619634
rect 73868 619366 74868 619398
rect 93868 619954 94868 619986
rect 93868 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 94868 619954
rect 93868 619634 94868 619718
rect 93868 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 94868 619634
rect 93868 619366 94868 619398
rect 113868 619954 114868 619986
rect 113868 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 114868 619954
rect 113868 619634 114868 619718
rect 113868 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 114868 619634
rect 113868 619366 114868 619398
rect 133868 619954 134868 619986
rect 133868 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 134868 619954
rect 133868 619634 134868 619718
rect 133868 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 134868 619634
rect 133868 619366 134868 619398
rect 153868 619954 154868 619986
rect 153868 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 154868 619954
rect 153868 619634 154868 619718
rect 153868 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 154868 619634
rect 153868 619366 154868 619398
rect 173868 619954 174868 619986
rect 173868 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 174868 619954
rect 173868 619634 174868 619718
rect 173868 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 174868 619634
rect 173868 619366 174868 619398
rect 193868 619954 194868 619986
rect 193868 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 194868 619954
rect 193868 619634 194868 619718
rect 193868 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 194868 619634
rect 193868 619366 194868 619398
rect 213868 619954 214868 619986
rect 213868 619718 213930 619954
rect 214166 619718 214250 619954
rect 214486 619718 214570 619954
rect 214806 619718 214868 619954
rect 213868 619634 214868 619718
rect 213868 619398 213930 619634
rect 214166 619398 214250 619634
rect 214486 619398 214570 619634
rect 214806 619398 214868 619634
rect 213868 619366 214868 619398
rect 233868 619954 234868 619986
rect 233868 619718 233930 619954
rect 234166 619718 234250 619954
rect 234486 619718 234570 619954
rect 234806 619718 234868 619954
rect 233868 619634 234868 619718
rect 233868 619398 233930 619634
rect 234166 619398 234250 619634
rect 234486 619398 234570 619634
rect 234806 619398 234868 619634
rect 233868 619366 234868 619398
rect 253868 619954 254868 619986
rect 253868 619718 253930 619954
rect 254166 619718 254250 619954
rect 254486 619718 254570 619954
rect 254806 619718 254868 619954
rect 253868 619634 254868 619718
rect 253868 619398 253930 619634
rect 254166 619398 254250 619634
rect 254486 619398 254570 619634
rect 254806 619398 254868 619634
rect 253868 619366 254868 619398
rect 273868 619954 274868 619986
rect 273868 619718 273930 619954
rect 274166 619718 274250 619954
rect 274486 619718 274570 619954
rect 274806 619718 274868 619954
rect 273868 619634 274868 619718
rect 273868 619398 273930 619634
rect 274166 619398 274250 619634
rect 274486 619398 274570 619634
rect 274806 619398 274868 619634
rect 273868 619366 274868 619398
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 23868 615454 24868 615486
rect 23868 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 24868 615454
rect 23868 615134 24868 615218
rect 23868 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 24868 615134
rect 23868 614866 24868 614898
rect 43868 615454 44868 615486
rect 43868 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 44868 615454
rect 43868 615134 44868 615218
rect 43868 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 44868 615134
rect 43868 614866 44868 614898
rect 63868 615454 64868 615486
rect 63868 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 64868 615454
rect 63868 615134 64868 615218
rect 63868 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 64868 615134
rect 63868 614866 64868 614898
rect 83868 615454 84868 615486
rect 83868 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 84868 615454
rect 83868 615134 84868 615218
rect 83868 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 84868 615134
rect 83868 614866 84868 614898
rect 103868 615454 104868 615486
rect 103868 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 104868 615454
rect 103868 615134 104868 615218
rect 103868 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 104868 615134
rect 103868 614866 104868 614898
rect 123868 615454 124868 615486
rect 123868 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 124868 615454
rect 123868 615134 124868 615218
rect 123868 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 124868 615134
rect 123868 614866 124868 614898
rect 143868 615454 144868 615486
rect 143868 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 144868 615454
rect 143868 615134 144868 615218
rect 143868 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 144868 615134
rect 143868 614866 144868 614898
rect 163868 615454 164868 615486
rect 163868 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 164868 615454
rect 163868 615134 164868 615218
rect 163868 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 164868 615134
rect 163868 614866 164868 614898
rect 183868 615454 184868 615486
rect 183868 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 184868 615454
rect 183868 615134 184868 615218
rect 183868 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 184868 615134
rect 183868 614866 184868 614898
rect 203868 615454 204868 615486
rect 203868 615218 203930 615454
rect 204166 615218 204250 615454
rect 204486 615218 204570 615454
rect 204806 615218 204868 615454
rect 203868 615134 204868 615218
rect 203868 614898 203930 615134
rect 204166 614898 204250 615134
rect 204486 614898 204570 615134
rect 204806 614898 204868 615134
rect 203868 614866 204868 614898
rect 223868 615454 224868 615486
rect 223868 615218 223930 615454
rect 224166 615218 224250 615454
rect 224486 615218 224570 615454
rect 224806 615218 224868 615454
rect 223868 615134 224868 615218
rect 223868 614898 223930 615134
rect 224166 614898 224250 615134
rect 224486 614898 224570 615134
rect 224806 614898 224868 615134
rect 223868 614866 224868 614898
rect 243868 615454 244868 615486
rect 243868 615218 243930 615454
rect 244166 615218 244250 615454
rect 244486 615218 244570 615454
rect 244806 615218 244868 615454
rect 243868 615134 244868 615218
rect 243868 614898 243930 615134
rect 244166 614898 244250 615134
rect 244486 614898 244570 615134
rect 244806 614898 244868 615134
rect 243868 614866 244868 614898
rect 263868 615454 264868 615486
rect 263868 615218 263930 615454
rect 264166 615218 264250 615454
rect 264486 615218 264570 615454
rect 264806 615218 264868 615454
rect 263868 615134 264868 615218
rect 263868 614898 263930 615134
rect 264166 614898 264250 615134
rect 264486 614898 264570 615134
rect 264806 614898 264868 615134
rect 263868 614866 264868 614898
rect 283868 615454 284868 615486
rect 283868 615218 283930 615454
rect 284166 615218 284250 615454
rect 284486 615218 284570 615454
rect 284806 615218 284868 615454
rect 283868 615134 284868 615218
rect 283868 614898 283930 615134
rect 284166 614898 284250 615134
rect 284486 614898 284570 615134
rect 284806 614898 284868 615134
rect 283868 614866 284868 614898
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 292619 586396 292685 586397
rect 292619 586332 292620 586396
rect 292684 586332 292685 586396
rect 292619 586331 292685 586332
rect 285627 585988 285693 585989
rect 285627 585924 285628 585988
rect 285692 585924 285693 585988
rect 285627 585923 285693 585924
rect 23243 585852 23309 585853
rect 23243 585788 23244 585852
rect 23308 585788 23309 585852
rect 23243 585787 23309 585788
rect 21955 585716 22021 585717
rect 21955 585652 21956 585716
rect 22020 585652 22021 585716
rect 21955 585651 22021 585652
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 18459 502484 18525 502485
rect 18459 502420 18460 502484
rect 18524 502420 18525 502484
rect 18459 502419 18525 502420
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 18462 21997 18522 502419
rect 21958 459509 22018 585651
rect 21955 459508 22021 459509
rect 21955 459444 21956 459508
rect 22020 459444 22021 459508
rect 21955 459443 22021 459444
rect 21958 335370 22018 459443
rect 23246 458149 23306 585787
rect 33868 547954 34868 547986
rect 33868 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 34868 547954
rect 33868 547634 34868 547718
rect 33868 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 34868 547634
rect 33868 547366 34868 547398
rect 53868 547954 54868 547986
rect 53868 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 54868 547954
rect 53868 547634 54868 547718
rect 53868 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 54868 547634
rect 53868 547366 54868 547398
rect 73868 547954 74868 547986
rect 73868 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 74868 547954
rect 73868 547634 74868 547718
rect 73868 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 74868 547634
rect 73868 547366 74868 547398
rect 93868 547954 94868 547986
rect 93868 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 94868 547954
rect 93868 547634 94868 547718
rect 93868 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 94868 547634
rect 93868 547366 94868 547398
rect 113868 547954 114868 547986
rect 113868 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 114868 547954
rect 113868 547634 114868 547718
rect 113868 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 114868 547634
rect 113868 547366 114868 547398
rect 133868 547954 134868 547986
rect 133868 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 134868 547954
rect 133868 547634 134868 547718
rect 133868 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 134868 547634
rect 133868 547366 134868 547398
rect 153868 547954 154868 547986
rect 153868 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 154868 547954
rect 153868 547634 154868 547718
rect 153868 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 154868 547634
rect 153868 547366 154868 547398
rect 173868 547954 174868 547986
rect 173868 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 174868 547954
rect 173868 547634 174868 547718
rect 173868 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 174868 547634
rect 173868 547366 174868 547398
rect 193868 547954 194868 547986
rect 193868 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 194868 547954
rect 193868 547634 194868 547718
rect 193868 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 194868 547634
rect 193868 547366 194868 547398
rect 213868 547954 214868 547986
rect 213868 547718 213930 547954
rect 214166 547718 214250 547954
rect 214486 547718 214570 547954
rect 214806 547718 214868 547954
rect 213868 547634 214868 547718
rect 213868 547398 213930 547634
rect 214166 547398 214250 547634
rect 214486 547398 214570 547634
rect 214806 547398 214868 547634
rect 213868 547366 214868 547398
rect 233868 547954 234868 547986
rect 233868 547718 233930 547954
rect 234166 547718 234250 547954
rect 234486 547718 234570 547954
rect 234806 547718 234868 547954
rect 233868 547634 234868 547718
rect 233868 547398 233930 547634
rect 234166 547398 234250 547634
rect 234486 547398 234570 547634
rect 234806 547398 234868 547634
rect 233868 547366 234868 547398
rect 253868 547954 254868 547986
rect 253868 547718 253930 547954
rect 254166 547718 254250 547954
rect 254486 547718 254570 547954
rect 254806 547718 254868 547954
rect 253868 547634 254868 547718
rect 253868 547398 253930 547634
rect 254166 547398 254250 547634
rect 254486 547398 254570 547634
rect 254806 547398 254868 547634
rect 253868 547366 254868 547398
rect 273868 547954 274868 547986
rect 273868 547718 273930 547954
rect 274166 547718 274250 547954
rect 274486 547718 274570 547954
rect 274806 547718 274868 547954
rect 273868 547634 274868 547718
rect 273868 547398 273930 547634
rect 274166 547398 274250 547634
rect 274486 547398 274570 547634
rect 274806 547398 274868 547634
rect 273868 547366 274868 547398
rect 23868 543454 24868 543486
rect 23868 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 24868 543454
rect 23868 543134 24868 543218
rect 23868 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 24868 543134
rect 23868 542866 24868 542898
rect 43868 543454 44868 543486
rect 43868 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 44868 543454
rect 43868 543134 44868 543218
rect 43868 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 44868 543134
rect 43868 542866 44868 542898
rect 63868 543454 64868 543486
rect 63868 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 64868 543454
rect 63868 543134 64868 543218
rect 63868 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 64868 543134
rect 63868 542866 64868 542898
rect 83868 543454 84868 543486
rect 83868 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 84868 543454
rect 83868 543134 84868 543218
rect 83868 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 84868 543134
rect 83868 542866 84868 542898
rect 103868 543454 104868 543486
rect 103868 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 104868 543454
rect 103868 543134 104868 543218
rect 103868 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 104868 543134
rect 103868 542866 104868 542898
rect 123868 543454 124868 543486
rect 123868 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 124868 543454
rect 123868 543134 124868 543218
rect 123868 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 124868 543134
rect 123868 542866 124868 542898
rect 143868 543454 144868 543486
rect 143868 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 144868 543454
rect 143868 543134 144868 543218
rect 143868 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 144868 543134
rect 143868 542866 144868 542898
rect 163868 543454 164868 543486
rect 163868 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 164868 543454
rect 163868 543134 164868 543218
rect 163868 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 164868 543134
rect 163868 542866 164868 542898
rect 183868 543454 184868 543486
rect 183868 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 184868 543454
rect 183868 543134 184868 543218
rect 183868 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 184868 543134
rect 183868 542866 184868 542898
rect 203868 543454 204868 543486
rect 203868 543218 203930 543454
rect 204166 543218 204250 543454
rect 204486 543218 204570 543454
rect 204806 543218 204868 543454
rect 203868 543134 204868 543218
rect 203868 542898 203930 543134
rect 204166 542898 204250 543134
rect 204486 542898 204570 543134
rect 204806 542898 204868 543134
rect 203868 542866 204868 542898
rect 223868 543454 224868 543486
rect 223868 543218 223930 543454
rect 224166 543218 224250 543454
rect 224486 543218 224570 543454
rect 224806 543218 224868 543454
rect 223868 543134 224868 543218
rect 223868 542898 223930 543134
rect 224166 542898 224250 543134
rect 224486 542898 224570 543134
rect 224806 542898 224868 543134
rect 223868 542866 224868 542898
rect 243868 543454 244868 543486
rect 243868 543218 243930 543454
rect 244166 543218 244250 543454
rect 244486 543218 244570 543454
rect 244806 543218 244868 543454
rect 243868 543134 244868 543218
rect 243868 542898 243930 543134
rect 244166 542898 244250 543134
rect 244486 542898 244570 543134
rect 244806 542898 244868 543134
rect 243868 542866 244868 542898
rect 263868 543454 264868 543486
rect 263868 543218 263930 543454
rect 264166 543218 264250 543454
rect 264486 543218 264570 543454
rect 264806 543218 264868 543454
rect 263868 543134 264868 543218
rect 263868 542898 263930 543134
rect 264166 542898 264250 543134
rect 264486 542898 264570 543134
rect 264806 542898 264868 543134
rect 263868 542866 264868 542898
rect 283868 543454 284868 543486
rect 283868 543218 283930 543454
rect 284166 543218 284250 543454
rect 284486 543218 284570 543454
rect 284806 543218 284868 543454
rect 283868 543134 284868 543218
rect 283868 542898 283930 543134
rect 284166 542898 284250 543134
rect 284486 542898 284570 543134
rect 284806 542898 284868 543134
rect 283868 542866 284868 542898
rect 33868 511954 34868 511986
rect 33868 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 34868 511954
rect 33868 511634 34868 511718
rect 33868 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 34868 511634
rect 33868 511366 34868 511398
rect 53868 511954 54868 511986
rect 53868 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 54868 511954
rect 53868 511634 54868 511718
rect 53868 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 54868 511634
rect 53868 511366 54868 511398
rect 73868 511954 74868 511986
rect 73868 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 74868 511954
rect 73868 511634 74868 511718
rect 73868 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 74868 511634
rect 73868 511366 74868 511398
rect 93868 511954 94868 511986
rect 93868 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 94868 511954
rect 93868 511634 94868 511718
rect 93868 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 94868 511634
rect 93868 511366 94868 511398
rect 113868 511954 114868 511986
rect 113868 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 114868 511954
rect 113868 511634 114868 511718
rect 113868 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 114868 511634
rect 113868 511366 114868 511398
rect 133868 511954 134868 511986
rect 133868 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 134868 511954
rect 133868 511634 134868 511718
rect 133868 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 134868 511634
rect 133868 511366 134868 511398
rect 153868 511954 154868 511986
rect 153868 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 154868 511954
rect 153868 511634 154868 511718
rect 153868 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 154868 511634
rect 153868 511366 154868 511398
rect 173868 511954 174868 511986
rect 173868 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 174868 511954
rect 173868 511634 174868 511718
rect 173868 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 174868 511634
rect 173868 511366 174868 511398
rect 193868 511954 194868 511986
rect 193868 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 194868 511954
rect 193868 511634 194868 511718
rect 193868 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 194868 511634
rect 193868 511366 194868 511398
rect 213868 511954 214868 511986
rect 213868 511718 213930 511954
rect 214166 511718 214250 511954
rect 214486 511718 214570 511954
rect 214806 511718 214868 511954
rect 213868 511634 214868 511718
rect 213868 511398 213930 511634
rect 214166 511398 214250 511634
rect 214486 511398 214570 511634
rect 214806 511398 214868 511634
rect 213868 511366 214868 511398
rect 233868 511954 234868 511986
rect 233868 511718 233930 511954
rect 234166 511718 234250 511954
rect 234486 511718 234570 511954
rect 234806 511718 234868 511954
rect 233868 511634 234868 511718
rect 233868 511398 233930 511634
rect 234166 511398 234250 511634
rect 234486 511398 234570 511634
rect 234806 511398 234868 511634
rect 233868 511366 234868 511398
rect 253868 511954 254868 511986
rect 253868 511718 253930 511954
rect 254166 511718 254250 511954
rect 254486 511718 254570 511954
rect 254806 511718 254868 511954
rect 253868 511634 254868 511718
rect 253868 511398 253930 511634
rect 254166 511398 254250 511634
rect 254486 511398 254570 511634
rect 254806 511398 254868 511634
rect 253868 511366 254868 511398
rect 273868 511954 274868 511986
rect 273868 511718 273930 511954
rect 274166 511718 274250 511954
rect 274486 511718 274570 511954
rect 274806 511718 274868 511954
rect 273868 511634 274868 511718
rect 273868 511398 273930 511634
rect 274166 511398 274250 511634
rect 274486 511398 274570 511634
rect 274806 511398 274868 511634
rect 273868 511366 274868 511398
rect 23868 507454 24868 507486
rect 23868 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 24868 507454
rect 23868 507134 24868 507218
rect 23868 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 24868 507134
rect 23868 506866 24868 506898
rect 43868 507454 44868 507486
rect 43868 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 44868 507454
rect 43868 507134 44868 507218
rect 43868 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 44868 507134
rect 43868 506866 44868 506898
rect 63868 507454 64868 507486
rect 63868 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 64868 507454
rect 63868 507134 64868 507218
rect 63868 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 64868 507134
rect 63868 506866 64868 506898
rect 83868 507454 84868 507486
rect 83868 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 84868 507454
rect 83868 507134 84868 507218
rect 83868 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 84868 507134
rect 83868 506866 84868 506898
rect 103868 507454 104868 507486
rect 103868 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 104868 507454
rect 103868 507134 104868 507218
rect 103868 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 104868 507134
rect 103868 506866 104868 506898
rect 123868 507454 124868 507486
rect 123868 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 124868 507454
rect 123868 507134 124868 507218
rect 123868 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 124868 507134
rect 123868 506866 124868 506898
rect 143868 507454 144868 507486
rect 143868 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 144868 507454
rect 143868 507134 144868 507218
rect 143868 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 144868 507134
rect 143868 506866 144868 506898
rect 163868 507454 164868 507486
rect 163868 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 164868 507454
rect 163868 507134 164868 507218
rect 163868 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 164868 507134
rect 163868 506866 164868 506898
rect 183868 507454 184868 507486
rect 183868 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 184868 507454
rect 183868 507134 184868 507218
rect 183868 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 184868 507134
rect 183868 506866 184868 506898
rect 203868 507454 204868 507486
rect 203868 507218 203930 507454
rect 204166 507218 204250 507454
rect 204486 507218 204570 507454
rect 204806 507218 204868 507454
rect 203868 507134 204868 507218
rect 203868 506898 203930 507134
rect 204166 506898 204250 507134
rect 204486 506898 204570 507134
rect 204806 506898 204868 507134
rect 203868 506866 204868 506898
rect 223868 507454 224868 507486
rect 223868 507218 223930 507454
rect 224166 507218 224250 507454
rect 224486 507218 224570 507454
rect 224806 507218 224868 507454
rect 223868 507134 224868 507218
rect 223868 506898 223930 507134
rect 224166 506898 224250 507134
rect 224486 506898 224570 507134
rect 224806 506898 224868 507134
rect 223868 506866 224868 506898
rect 243868 507454 244868 507486
rect 243868 507218 243930 507454
rect 244166 507218 244250 507454
rect 244486 507218 244570 507454
rect 244806 507218 244868 507454
rect 243868 507134 244868 507218
rect 243868 506898 243930 507134
rect 244166 506898 244250 507134
rect 244486 506898 244570 507134
rect 244806 506898 244868 507134
rect 243868 506866 244868 506898
rect 263868 507454 264868 507486
rect 263868 507218 263930 507454
rect 264166 507218 264250 507454
rect 264486 507218 264570 507454
rect 264806 507218 264868 507454
rect 263868 507134 264868 507218
rect 263868 506898 263930 507134
rect 264166 506898 264250 507134
rect 264486 506898 264570 507134
rect 264806 506898 264868 507134
rect 263868 506866 264868 506898
rect 283868 507454 284868 507486
rect 283868 507218 283930 507454
rect 284166 507218 284250 507454
rect 284486 507218 284570 507454
rect 284806 507218 284868 507454
rect 283868 507134 284868 507218
rect 283868 506898 283930 507134
rect 284166 506898 284250 507134
rect 284486 506898 284570 507134
rect 284806 506898 284868 507134
rect 283868 506866 284868 506898
rect 33868 475954 34868 475986
rect 33868 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 34868 475954
rect 33868 475634 34868 475718
rect 33868 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 34868 475634
rect 33868 475366 34868 475398
rect 53868 475954 54868 475986
rect 53868 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 54868 475954
rect 53868 475634 54868 475718
rect 53868 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 54868 475634
rect 53868 475366 54868 475398
rect 73868 475954 74868 475986
rect 73868 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 74868 475954
rect 73868 475634 74868 475718
rect 73868 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 74868 475634
rect 73868 475366 74868 475398
rect 93868 475954 94868 475986
rect 93868 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 94868 475954
rect 93868 475634 94868 475718
rect 93868 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 94868 475634
rect 93868 475366 94868 475398
rect 113868 475954 114868 475986
rect 113868 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 114868 475954
rect 113868 475634 114868 475718
rect 113868 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 114868 475634
rect 113868 475366 114868 475398
rect 133868 475954 134868 475986
rect 133868 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 134868 475954
rect 133868 475634 134868 475718
rect 133868 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 134868 475634
rect 133868 475366 134868 475398
rect 153868 475954 154868 475986
rect 153868 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 154868 475954
rect 153868 475634 154868 475718
rect 153868 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 154868 475634
rect 153868 475366 154868 475398
rect 173868 475954 174868 475986
rect 173868 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 174868 475954
rect 173868 475634 174868 475718
rect 173868 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 174868 475634
rect 173868 475366 174868 475398
rect 193868 475954 194868 475986
rect 193868 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 194868 475954
rect 193868 475634 194868 475718
rect 193868 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 194868 475634
rect 193868 475366 194868 475398
rect 213868 475954 214868 475986
rect 213868 475718 213930 475954
rect 214166 475718 214250 475954
rect 214486 475718 214570 475954
rect 214806 475718 214868 475954
rect 213868 475634 214868 475718
rect 213868 475398 213930 475634
rect 214166 475398 214250 475634
rect 214486 475398 214570 475634
rect 214806 475398 214868 475634
rect 213868 475366 214868 475398
rect 233868 475954 234868 475986
rect 233868 475718 233930 475954
rect 234166 475718 234250 475954
rect 234486 475718 234570 475954
rect 234806 475718 234868 475954
rect 233868 475634 234868 475718
rect 233868 475398 233930 475634
rect 234166 475398 234250 475634
rect 234486 475398 234570 475634
rect 234806 475398 234868 475634
rect 233868 475366 234868 475398
rect 253868 475954 254868 475986
rect 253868 475718 253930 475954
rect 254166 475718 254250 475954
rect 254486 475718 254570 475954
rect 254806 475718 254868 475954
rect 253868 475634 254868 475718
rect 253868 475398 253930 475634
rect 254166 475398 254250 475634
rect 254486 475398 254570 475634
rect 254806 475398 254868 475634
rect 253868 475366 254868 475398
rect 273868 475954 274868 475986
rect 273868 475718 273930 475954
rect 274166 475718 274250 475954
rect 274486 475718 274570 475954
rect 274806 475718 274868 475954
rect 273868 475634 274868 475718
rect 273868 475398 273930 475634
rect 274166 475398 274250 475634
rect 274486 475398 274570 475634
rect 274806 475398 274868 475634
rect 273868 475366 274868 475398
rect 23868 471454 24868 471486
rect 23868 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 24868 471454
rect 23868 471134 24868 471218
rect 23868 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 24868 471134
rect 23868 470866 24868 470898
rect 43868 471454 44868 471486
rect 43868 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 44868 471454
rect 43868 471134 44868 471218
rect 43868 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 44868 471134
rect 43868 470866 44868 470898
rect 63868 471454 64868 471486
rect 63868 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 64868 471454
rect 63868 471134 64868 471218
rect 63868 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 64868 471134
rect 63868 470866 64868 470898
rect 83868 471454 84868 471486
rect 83868 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 84868 471454
rect 83868 471134 84868 471218
rect 83868 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 84868 471134
rect 83868 470866 84868 470898
rect 103868 471454 104868 471486
rect 103868 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 104868 471454
rect 103868 471134 104868 471218
rect 103868 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 104868 471134
rect 103868 470866 104868 470898
rect 123868 471454 124868 471486
rect 123868 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 124868 471454
rect 123868 471134 124868 471218
rect 123868 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 124868 471134
rect 123868 470866 124868 470898
rect 143868 471454 144868 471486
rect 143868 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 144868 471454
rect 143868 471134 144868 471218
rect 143868 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 144868 471134
rect 143868 470866 144868 470898
rect 163868 471454 164868 471486
rect 163868 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 164868 471454
rect 163868 471134 164868 471218
rect 163868 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 164868 471134
rect 163868 470866 164868 470898
rect 183868 471454 184868 471486
rect 183868 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 184868 471454
rect 183868 471134 184868 471218
rect 183868 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 184868 471134
rect 183868 470866 184868 470898
rect 203868 471454 204868 471486
rect 203868 471218 203930 471454
rect 204166 471218 204250 471454
rect 204486 471218 204570 471454
rect 204806 471218 204868 471454
rect 203868 471134 204868 471218
rect 203868 470898 203930 471134
rect 204166 470898 204250 471134
rect 204486 470898 204570 471134
rect 204806 470898 204868 471134
rect 203868 470866 204868 470898
rect 223868 471454 224868 471486
rect 223868 471218 223930 471454
rect 224166 471218 224250 471454
rect 224486 471218 224570 471454
rect 224806 471218 224868 471454
rect 223868 471134 224868 471218
rect 223868 470898 223930 471134
rect 224166 470898 224250 471134
rect 224486 470898 224570 471134
rect 224806 470898 224868 471134
rect 223868 470866 224868 470898
rect 243868 471454 244868 471486
rect 243868 471218 243930 471454
rect 244166 471218 244250 471454
rect 244486 471218 244570 471454
rect 244806 471218 244868 471454
rect 243868 471134 244868 471218
rect 243868 470898 243930 471134
rect 244166 470898 244250 471134
rect 244486 470898 244570 471134
rect 244806 470898 244868 471134
rect 243868 470866 244868 470898
rect 263868 471454 264868 471486
rect 263868 471218 263930 471454
rect 264166 471218 264250 471454
rect 264486 471218 264570 471454
rect 264806 471218 264868 471454
rect 263868 471134 264868 471218
rect 263868 470898 263930 471134
rect 264166 470898 264250 471134
rect 264486 470898 264570 471134
rect 264806 470898 264868 471134
rect 263868 470866 264868 470898
rect 283868 471454 284868 471486
rect 283868 471218 283930 471454
rect 284166 471218 284250 471454
rect 284486 471218 284570 471454
rect 284806 471218 284868 471454
rect 283868 471134 284868 471218
rect 283868 470898 283930 471134
rect 284166 470898 284250 471134
rect 284486 470898 284570 471134
rect 284806 470898 284868 471134
rect 283868 470866 284868 470898
rect 285630 458149 285690 585923
rect 287099 585852 287165 585853
rect 287099 585788 287100 585852
rect 287164 585788 287165 585852
rect 287099 585787 287165 585788
rect 287102 461005 287162 585787
rect 288387 585716 288453 585717
rect 288387 585652 288388 585716
rect 288452 585652 288453 585716
rect 288387 585651 288453 585652
rect 291699 585716 291765 585717
rect 291699 585652 291700 585716
rect 291764 585652 291765 585716
rect 291699 585651 291765 585652
rect 287099 461004 287165 461005
rect 287099 460940 287100 461004
rect 287164 460940 287165 461004
rect 287099 460939 287165 460940
rect 23243 458148 23309 458149
rect 23243 458084 23244 458148
rect 23308 458084 23309 458148
rect 23243 458083 23309 458084
rect 285627 458148 285693 458149
rect 285627 458084 285628 458148
rect 285692 458084 285693 458148
rect 285627 458083 285693 458084
rect 23246 335370 23306 458083
rect 33868 439954 34868 439986
rect 33868 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 34868 439954
rect 33868 439634 34868 439718
rect 33868 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 34868 439634
rect 33868 439366 34868 439398
rect 53868 439954 54868 439986
rect 53868 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 54868 439954
rect 53868 439634 54868 439718
rect 53868 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 54868 439634
rect 53868 439366 54868 439398
rect 73868 439954 74868 439986
rect 73868 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 74868 439954
rect 73868 439634 74868 439718
rect 73868 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 74868 439634
rect 73868 439366 74868 439398
rect 93868 439954 94868 439986
rect 93868 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 94868 439954
rect 93868 439634 94868 439718
rect 93868 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 94868 439634
rect 93868 439366 94868 439398
rect 113868 439954 114868 439986
rect 113868 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 114868 439954
rect 113868 439634 114868 439718
rect 113868 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 114868 439634
rect 113868 439366 114868 439398
rect 133868 439954 134868 439986
rect 133868 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 134868 439954
rect 133868 439634 134868 439718
rect 133868 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 134868 439634
rect 133868 439366 134868 439398
rect 153868 439954 154868 439986
rect 153868 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 154868 439954
rect 153868 439634 154868 439718
rect 153868 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 154868 439634
rect 153868 439366 154868 439398
rect 173868 439954 174868 439986
rect 173868 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 174868 439954
rect 173868 439634 174868 439718
rect 173868 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 174868 439634
rect 173868 439366 174868 439398
rect 193868 439954 194868 439986
rect 193868 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 194868 439954
rect 193868 439634 194868 439718
rect 193868 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 194868 439634
rect 193868 439366 194868 439398
rect 213868 439954 214868 439986
rect 213868 439718 213930 439954
rect 214166 439718 214250 439954
rect 214486 439718 214570 439954
rect 214806 439718 214868 439954
rect 213868 439634 214868 439718
rect 213868 439398 213930 439634
rect 214166 439398 214250 439634
rect 214486 439398 214570 439634
rect 214806 439398 214868 439634
rect 213868 439366 214868 439398
rect 233868 439954 234868 439986
rect 233868 439718 233930 439954
rect 234166 439718 234250 439954
rect 234486 439718 234570 439954
rect 234806 439718 234868 439954
rect 233868 439634 234868 439718
rect 233868 439398 233930 439634
rect 234166 439398 234250 439634
rect 234486 439398 234570 439634
rect 234806 439398 234868 439634
rect 233868 439366 234868 439398
rect 253868 439954 254868 439986
rect 253868 439718 253930 439954
rect 254166 439718 254250 439954
rect 254486 439718 254570 439954
rect 254806 439718 254868 439954
rect 253868 439634 254868 439718
rect 253868 439398 253930 439634
rect 254166 439398 254250 439634
rect 254486 439398 254570 439634
rect 254806 439398 254868 439634
rect 253868 439366 254868 439398
rect 273868 439954 274868 439986
rect 273868 439718 273930 439954
rect 274166 439718 274250 439954
rect 274486 439718 274570 439954
rect 274806 439718 274868 439954
rect 273868 439634 274868 439718
rect 273868 439398 273930 439634
rect 274166 439398 274250 439634
rect 274486 439398 274570 439634
rect 274806 439398 274868 439634
rect 273868 439366 274868 439398
rect 23868 435454 24868 435486
rect 23868 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 24868 435454
rect 23868 435134 24868 435218
rect 23868 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 24868 435134
rect 23868 434866 24868 434898
rect 43868 435454 44868 435486
rect 43868 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 44868 435454
rect 43868 435134 44868 435218
rect 43868 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 44868 435134
rect 43868 434866 44868 434898
rect 63868 435454 64868 435486
rect 63868 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 64868 435454
rect 63868 435134 64868 435218
rect 63868 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 64868 435134
rect 63868 434866 64868 434898
rect 83868 435454 84868 435486
rect 83868 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 84868 435454
rect 83868 435134 84868 435218
rect 83868 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 84868 435134
rect 83868 434866 84868 434898
rect 103868 435454 104868 435486
rect 103868 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 104868 435454
rect 103868 435134 104868 435218
rect 103868 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 104868 435134
rect 103868 434866 104868 434898
rect 123868 435454 124868 435486
rect 123868 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 124868 435454
rect 123868 435134 124868 435218
rect 123868 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 124868 435134
rect 123868 434866 124868 434898
rect 143868 435454 144868 435486
rect 143868 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 144868 435454
rect 143868 435134 144868 435218
rect 143868 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 144868 435134
rect 143868 434866 144868 434898
rect 163868 435454 164868 435486
rect 163868 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 164868 435454
rect 163868 435134 164868 435218
rect 163868 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 164868 435134
rect 163868 434866 164868 434898
rect 183868 435454 184868 435486
rect 183868 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 184868 435454
rect 183868 435134 184868 435218
rect 183868 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 184868 435134
rect 183868 434866 184868 434898
rect 203868 435454 204868 435486
rect 203868 435218 203930 435454
rect 204166 435218 204250 435454
rect 204486 435218 204570 435454
rect 204806 435218 204868 435454
rect 203868 435134 204868 435218
rect 203868 434898 203930 435134
rect 204166 434898 204250 435134
rect 204486 434898 204570 435134
rect 204806 434898 204868 435134
rect 203868 434866 204868 434898
rect 223868 435454 224868 435486
rect 223868 435218 223930 435454
rect 224166 435218 224250 435454
rect 224486 435218 224570 435454
rect 224806 435218 224868 435454
rect 223868 435134 224868 435218
rect 223868 434898 223930 435134
rect 224166 434898 224250 435134
rect 224486 434898 224570 435134
rect 224806 434898 224868 435134
rect 223868 434866 224868 434898
rect 243868 435454 244868 435486
rect 243868 435218 243930 435454
rect 244166 435218 244250 435454
rect 244486 435218 244570 435454
rect 244806 435218 244868 435454
rect 243868 435134 244868 435218
rect 243868 434898 243930 435134
rect 244166 434898 244250 435134
rect 244486 434898 244570 435134
rect 244806 434898 244868 435134
rect 243868 434866 244868 434898
rect 263868 435454 264868 435486
rect 263868 435218 263930 435454
rect 264166 435218 264250 435454
rect 264486 435218 264570 435454
rect 264806 435218 264868 435454
rect 263868 435134 264868 435218
rect 263868 434898 263930 435134
rect 264166 434898 264250 435134
rect 264486 434898 264570 435134
rect 264806 434898 264868 435134
rect 263868 434866 264868 434898
rect 283868 435454 284868 435486
rect 283868 435218 283930 435454
rect 284166 435218 284250 435454
rect 284486 435218 284570 435454
rect 284806 435218 284868 435454
rect 283868 435134 284868 435218
rect 283868 434898 283930 435134
rect 284166 434898 284250 435134
rect 284486 434898 284570 435134
rect 284806 434898 284868 435134
rect 283868 434866 284868 434898
rect 33868 403954 34868 403986
rect 33868 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 34868 403954
rect 33868 403634 34868 403718
rect 33868 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 34868 403634
rect 33868 403366 34868 403398
rect 53868 403954 54868 403986
rect 53868 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 54868 403954
rect 53868 403634 54868 403718
rect 53868 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 54868 403634
rect 53868 403366 54868 403398
rect 73868 403954 74868 403986
rect 73868 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 74868 403954
rect 73868 403634 74868 403718
rect 73868 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 74868 403634
rect 73868 403366 74868 403398
rect 93868 403954 94868 403986
rect 93868 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 94868 403954
rect 93868 403634 94868 403718
rect 93868 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 94868 403634
rect 93868 403366 94868 403398
rect 113868 403954 114868 403986
rect 113868 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 114868 403954
rect 113868 403634 114868 403718
rect 113868 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 114868 403634
rect 113868 403366 114868 403398
rect 133868 403954 134868 403986
rect 133868 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 134868 403954
rect 133868 403634 134868 403718
rect 133868 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 134868 403634
rect 133868 403366 134868 403398
rect 153868 403954 154868 403986
rect 153868 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 154868 403954
rect 153868 403634 154868 403718
rect 153868 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 154868 403634
rect 153868 403366 154868 403398
rect 173868 403954 174868 403986
rect 173868 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 174868 403954
rect 173868 403634 174868 403718
rect 173868 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 174868 403634
rect 173868 403366 174868 403398
rect 193868 403954 194868 403986
rect 193868 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 194868 403954
rect 193868 403634 194868 403718
rect 193868 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 194868 403634
rect 193868 403366 194868 403398
rect 213868 403954 214868 403986
rect 213868 403718 213930 403954
rect 214166 403718 214250 403954
rect 214486 403718 214570 403954
rect 214806 403718 214868 403954
rect 213868 403634 214868 403718
rect 213868 403398 213930 403634
rect 214166 403398 214250 403634
rect 214486 403398 214570 403634
rect 214806 403398 214868 403634
rect 213868 403366 214868 403398
rect 233868 403954 234868 403986
rect 233868 403718 233930 403954
rect 234166 403718 234250 403954
rect 234486 403718 234570 403954
rect 234806 403718 234868 403954
rect 233868 403634 234868 403718
rect 233868 403398 233930 403634
rect 234166 403398 234250 403634
rect 234486 403398 234570 403634
rect 234806 403398 234868 403634
rect 233868 403366 234868 403398
rect 253868 403954 254868 403986
rect 253868 403718 253930 403954
rect 254166 403718 254250 403954
rect 254486 403718 254570 403954
rect 254806 403718 254868 403954
rect 253868 403634 254868 403718
rect 253868 403398 253930 403634
rect 254166 403398 254250 403634
rect 254486 403398 254570 403634
rect 254806 403398 254868 403634
rect 253868 403366 254868 403398
rect 273868 403954 274868 403986
rect 273868 403718 273930 403954
rect 274166 403718 274250 403954
rect 274486 403718 274570 403954
rect 274806 403718 274868 403954
rect 273868 403634 274868 403718
rect 273868 403398 273930 403634
rect 274166 403398 274250 403634
rect 274486 403398 274570 403634
rect 274806 403398 274868 403634
rect 273868 403366 274868 403398
rect 23868 399454 24868 399486
rect 23868 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 24868 399454
rect 23868 399134 24868 399218
rect 23868 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 24868 399134
rect 23868 398866 24868 398898
rect 43868 399454 44868 399486
rect 43868 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 44868 399454
rect 43868 399134 44868 399218
rect 43868 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 44868 399134
rect 43868 398866 44868 398898
rect 63868 399454 64868 399486
rect 63868 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 64868 399454
rect 63868 399134 64868 399218
rect 63868 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 64868 399134
rect 63868 398866 64868 398898
rect 83868 399454 84868 399486
rect 83868 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 84868 399454
rect 83868 399134 84868 399218
rect 83868 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 84868 399134
rect 83868 398866 84868 398898
rect 103868 399454 104868 399486
rect 103868 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 104868 399454
rect 103868 399134 104868 399218
rect 103868 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 104868 399134
rect 103868 398866 104868 398898
rect 123868 399454 124868 399486
rect 123868 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 124868 399454
rect 123868 399134 124868 399218
rect 123868 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 124868 399134
rect 123868 398866 124868 398898
rect 143868 399454 144868 399486
rect 143868 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 144868 399454
rect 143868 399134 144868 399218
rect 143868 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 144868 399134
rect 143868 398866 144868 398898
rect 163868 399454 164868 399486
rect 163868 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 164868 399454
rect 163868 399134 164868 399218
rect 163868 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 164868 399134
rect 163868 398866 164868 398898
rect 183868 399454 184868 399486
rect 183868 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 184868 399454
rect 183868 399134 184868 399218
rect 183868 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 184868 399134
rect 183868 398866 184868 398898
rect 203868 399454 204868 399486
rect 203868 399218 203930 399454
rect 204166 399218 204250 399454
rect 204486 399218 204570 399454
rect 204806 399218 204868 399454
rect 203868 399134 204868 399218
rect 203868 398898 203930 399134
rect 204166 398898 204250 399134
rect 204486 398898 204570 399134
rect 204806 398898 204868 399134
rect 203868 398866 204868 398898
rect 223868 399454 224868 399486
rect 223868 399218 223930 399454
rect 224166 399218 224250 399454
rect 224486 399218 224570 399454
rect 224806 399218 224868 399454
rect 223868 399134 224868 399218
rect 223868 398898 223930 399134
rect 224166 398898 224250 399134
rect 224486 398898 224570 399134
rect 224806 398898 224868 399134
rect 223868 398866 224868 398898
rect 243868 399454 244868 399486
rect 243868 399218 243930 399454
rect 244166 399218 244250 399454
rect 244486 399218 244570 399454
rect 244806 399218 244868 399454
rect 243868 399134 244868 399218
rect 243868 398898 243930 399134
rect 244166 398898 244250 399134
rect 244486 398898 244570 399134
rect 244806 398898 244868 399134
rect 243868 398866 244868 398898
rect 263868 399454 264868 399486
rect 263868 399218 263930 399454
rect 264166 399218 264250 399454
rect 264486 399218 264570 399454
rect 264806 399218 264868 399454
rect 263868 399134 264868 399218
rect 263868 398898 263930 399134
rect 264166 398898 264250 399134
rect 264486 398898 264570 399134
rect 264806 398898 264868 399134
rect 263868 398866 264868 398898
rect 283868 399454 284868 399486
rect 283868 399218 283930 399454
rect 284166 399218 284250 399454
rect 284486 399218 284570 399454
rect 284806 399218 284868 399454
rect 283868 399134 284868 399218
rect 283868 398898 283930 399134
rect 284166 398898 284250 399134
rect 284486 398898 284570 399134
rect 284806 398898 284868 399134
rect 283868 398866 284868 398898
rect 33868 367954 34868 367986
rect 33868 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 34868 367954
rect 33868 367634 34868 367718
rect 33868 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 34868 367634
rect 33868 367366 34868 367398
rect 53868 367954 54868 367986
rect 53868 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 54868 367954
rect 53868 367634 54868 367718
rect 53868 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 54868 367634
rect 53868 367366 54868 367398
rect 73868 367954 74868 367986
rect 73868 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 74868 367954
rect 73868 367634 74868 367718
rect 73868 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 74868 367634
rect 73868 367366 74868 367398
rect 93868 367954 94868 367986
rect 93868 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 94868 367954
rect 93868 367634 94868 367718
rect 93868 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 94868 367634
rect 93868 367366 94868 367398
rect 113868 367954 114868 367986
rect 113868 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 114868 367954
rect 113868 367634 114868 367718
rect 113868 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 114868 367634
rect 113868 367366 114868 367398
rect 133868 367954 134868 367986
rect 133868 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 134868 367954
rect 133868 367634 134868 367718
rect 133868 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 134868 367634
rect 133868 367366 134868 367398
rect 153868 367954 154868 367986
rect 153868 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 154868 367954
rect 153868 367634 154868 367718
rect 153868 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 154868 367634
rect 153868 367366 154868 367398
rect 173868 367954 174868 367986
rect 173868 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 174868 367954
rect 173868 367634 174868 367718
rect 173868 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 174868 367634
rect 173868 367366 174868 367398
rect 193868 367954 194868 367986
rect 193868 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 194868 367954
rect 193868 367634 194868 367718
rect 193868 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 194868 367634
rect 193868 367366 194868 367398
rect 213868 367954 214868 367986
rect 213868 367718 213930 367954
rect 214166 367718 214250 367954
rect 214486 367718 214570 367954
rect 214806 367718 214868 367954
rect 213868 367634 214868 367718
rect 213868 367398 213930 367634
rect 214166 367398 214250 367634
rect 214486 367398 214570 367634
rect 214806 367398 214868 367634
rect 213868 367366 214868 367398
rect 233868 367954 234868 367986
rect 233868 367718 233930 367954
rect 234166 367718 234250 367954
rect 234486 367718 234570 367954
rect 234806 367718 234868 367954
rect 233868 367634 234868 367718
rect 233868 367398 233930 367634
rect 234166 367398 234250 367634
rect 234486 367398 234570 367634
rect 234806 367398 234868 367634
rect 233868 367366 234868 367398
rect 253868 367954 254868 367986
rect 253868 367718 253930 367954
rect 254166 367718 254250 367954
rect 254486 367718 254570 367954
rect 254806 367718 254868 367954
rect 253868 367634 254868 367718
rect 253868 367398 253930 367634
rect 254166 367398 254250 367634
rect 254486 367398 254570 367634
rect 254806 367398 254868 367634
rect 253868 367366 254868 367398
rect 273868 367954 274868 367986
rect 273868 367718 273930 367954
rect 274166 367718 274250 367954
rect 274486 367718 274570 367954
rect 274806 367718 274868 367954
rect 273868 367634 274868 367718
rect 273868 367398 273930 367634
rect 274166 367398 274250 367634
rect 274486 367398 274570 367634
rect 274806 367398 274868 367634
rect 273868 367366 274868 367398
rect 23868 363454 24868 363486
rect 23868 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 24868 363454
rect 23868 363134 24868 363218
rect 23868 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 24868 363134
rect 23868 362866 24868 362898
rect 43868 363454 44868 363486
rect 43868 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 44868 363454
rect 43868 363134 44868 363218
rect 43868 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 44868 363134
rect 43868 362866 44868 362898
rect 63868 363454 64868 363486
rect 63868 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 64868 363454
rect 63868 363134 64868 363218
rect 63868 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 64868 363134
rect 63868 362866 64868 362898
rect 83868 363454 84868 363486
rect 83868 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 84868 363454
rect 83868 363134 84868 363218
rect 83868 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 84868 363134
rect 83868 362866 84868 362898
rect 103868 363454 104868 363486
rect 103868 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 104868 363454
rect 103868 363134 104868 363218
rect 103868 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 104868 363134
rect 103868 362866 104868 362898
rect 123868 363454 124868 363486
rect 123868 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 124868 363454
rect 123868 363134 124868 363218
rect 123868 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 124868 363134
rect 123868 362866 124868 362898
rect 143868 363454 144868 363486
rect 143868 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 144868 363454
rect 143868 363134 144868 363218
rect 143868 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 144868 363134
rect 143868 362866 144868 362898
rect 163868 363454 164868 363486
rect 163868 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 164868 363454
rect 163868 363134 164868 363218
rect 163868 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 164868 363134
rect 163868 362866 164868 362898
rect 183868 363454 184868 363486
rect 183868 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 184868 363454
rect 183868 363134 184868 363218
rect 183868 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 184868 363134
rect 183868 362866 184868 362898
rect 203868 363454 204868 363486
rect 203868 363218 203930 363454
rect 204166 363218 204250 363454
rect 204486 363218 204570 363454
rect 204806 363218 204868 363454
rect 203868 363134 204868 363218
rect 203868 362898 203930 363134
rect 204166 362898 204250 363134
rect 204486 362898 204570 363134
rect 204806 362898 204868 363134
rect 203868 362866 204868 362898
rect 223868 363454 224868 363486
rect 223868 363218 223930 363454
rect 224166 363218 224250 363454
rect 224486 363218 224570 363454
rect 224806 363218 224868 363454
rect 223868 363134 224868 363218
rect 223868 362898 223930 363134
rect 224166 362898 224250 363134
rect 224486 362898 224570 363134
rect 224806 362898 224868 363134
rect 223868 362866 224868 362898
rect 243868 363454 244868 363486
rect 243868 363218 243930 363454
rect 244166 363218 244250 363454
rect 244486 363218 244570 363454
rect 244806 363218 244868 363454
rect 243868 363134 244868 363218
rect 243868 362898 243930 363134
rect 244166 362898 244250 363134
rect 244486 362898 244570 363134
rect 244806 362898 244868 363134
rect 243868 362866 244868 362898
rect 263868 363454 264868 363486
rect 263868 363218 263930 363454
rect 264166 363218 264250 363454
rect 264486 363218 264570 363454
rect 264806 363218 264868 363454
rect 263868 363134 264868 363218
rect 263868 362898 263930 363134
rect 264166 362898 264250 363134
rect 264486 362898 264570 363134
rect 264806 362898 264868 363134
rect 263868 362866 264868 362898
rect 283868 363454 284868 363486
rect 283868 363218 283930 363454
rect 284166 363218 284250 363454
rect 284486 363218 284570 363454
rect 284806 363218 284868 363454
rect 283868 363134 284868 363218
rect 283868 362898 283930 363134
rect 284166 362898 284250 363134
rect 284486 362898 284570 363134
rect 284806 362898 284868 363134
rect 283868 362866 284868 362898
rect 21222 335310 22018 335370
rect 22694 335310 23306 335370
rect 21222 332893 21282 335310
rect 21219 332892 21285 332893
rect 21219 332828 21220 332892
rect 21284 332828 21285 332892
rect 21219 332827 21285 332828
rect 21222 202877 21282 332827
rect 22694 332213 22754 335310
rect 22691 332212 22757 332213
rect 22691 332148 22692 332212
rect 22756 332148 22757 332212
rect 22691 332147 22757 332148
rect 21403 207772 21469 207773
rect 21403 207708 21404 207772
rect 21468 207708 21469 207772
rect 21403 207707 21469 207708
rect 21406 206277 21466 207707
rect 22139 207636 22205 207637
rect 22139 207572 22140 207636
rect 22204 207572 22205 207636
rect 22139 207571 22205 207572
rect 22142 206413 22202 207571
rect 22139 206412 22205 206413
rect 22139 206348 22140 206412
rect 22204 206348 22205 206412
rect 22139 206347 22205 206348
rect 21403 206276 21469 206277
rect 21403 206212 21404 206276
rect 21468 206212 21469 206276
rect 21403 206211 21469 206212
rect 21955 203828 22021 203829
rect 21955 203764 21956 203828
rect 22020 203764 22021 203828
rect 21955 203763 22021 203764
rect 21219 202876 21285 202877
rect 21219 202812 21220 202876
rect 21284 202812 21285 202876
rect 21219 202811 21285 202812
rect 19931 200020 19997 200021
rect 19931 199956 19932 200020
rect 19996 199956 19997 200020
rect 19931 199955 19997 199956
rect 19563 110532 19629 110533
rect 19563 110468 19564 110532
rect 19628 110468 19629 110532
rect 19563 110467 19629 110468
rect 18459 21996 18525 21997
rect 18459 21932 18460 21996
rect 18524 21932 18525 21996
rect 18459 21931 18525 21932
rect 19566 21861 19626 110467
rect 19934 80205 19994 199955
rect 19931 80204 19997 80205
rect 19931 80140 19932 80204
rect 19996 80140 19997 80204
rect 19931 80139 19997 80140
rect 19794 57454 20414 76000
rect 21958 75853 22018 203763
rect 22694 202877 22754 332147
rect 285630 331397 285690 458083
rect 287651 457876 287717 457877
rect 287651 457812 287652 457876
rect 287716 457812 287717 457876
rect 287651 457811 287717 457812
rect 286179 444956 286245 444957
rect 286179 444892 286180 444956
rect 286244 444892 286245 444956
rect 286179 444891 286245 444892
rect 285627 331396 285693 331397
rect 285627 331332 285628 331396
rect 285692 331332 285693 331396
rect 285627 331331 285693 331332
rect 33868 295954 34868 295986
rect 33868 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 34868 295954
rect 33868 295634 34868 295718
rect 33868 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 34868 295634
rect 33868 295366 34868 295398
rect 53868 295954 54868 295986
rect 53868 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 54868 295954
rect 53868 295634 54868 295718
rect 53868 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 54868 295634
rect 53868 295366 54868 295398
rect 73868 295954 74868 295986
rect 73868 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 74868 295954
rect 73868 295634 74868 295718
rect 73868 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 74868 295634
rect 73868 295366 74868 295398
rect 93868 295954 94868 295986
rect 93868 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 94868 295954
rect 93868 295634 94868 295718
rect 93868 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 94868 295634
rect 93868 295366 94868 295398
rect 113868 295954 114868 295986
rect 113868 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 114868 295954
rect 113868 295634 114868 295718
rect 113868 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 114868 295634
rect 113868 295366 114868 295398
rect 133868 295954 134868 295986
rect 133868 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 134868 295954
rect 133868 295634 134868 295718
rect 133868 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 134868 295634
rect 133868 295366 134868 295398
rect 153868 295954 154868 295986
rect 153868 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 154868 295954
rect 153868 295634 154868 295718
rect 153868 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 154868 295634
rect 153868 295366 154868 295398
rect 173868 295954 174868 295986
rect 173868 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 174868 295954
rect 173868 295634 174868 295718
rect 173868 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 174868 295634
rect 173868 295366 174868 295398
rect 193868 295954 194868 295986
rect 193868 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 194868 295954
rect 193868 295634 194868 295718
rect 193868 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 194868 295634
rect 193868 295366 194868 295398
rect 213868 295954 214868 295986
rect 213868 295718 213930 295954
rect 214166 295718 214250 295954
rect 214486 295718 214570 295954
rect 214806 295718 214868 295954
rect 213868 295634 214868 295718
rect 213868 295398 213930 295634
rect 214166 295398 214250 295634
rect 214486 295398 214570 295634
rect 214806 295398 214868 295634
rect 213868 295366 214868 295398
rect 233868 295954 234868 295986
rect 233868 295718 233930 295954
rect 234166 295718 234250 295954
rect 234486 295718 234570 295954
rect 234806 295718 234868 295954
rect 233868 295634 234868 295718
rect 233868 295398 233930 295634
rect 234166 295398 234250 295634
rect 234486 295398 234570 295634
rect 234806 295398 234868 295634
rect 233868 295366 234868 295398
rect 253868 295954 254868 295986
rect 253868 295718 253930 295954
rect 254166 295718 254250 295954
rect 254486 295718 254570 295954
rect 254806 295718 254868 295954
rect 253868 295634 254868 295718
rect 253868 295398 253930 295634
rect 254166 295398 254250 295634
rect 254486 295398 254570 295634
rect 254806 295398 254868 295634
rect 253868 295366 254868 295398
rect 273868 295954 274868 295986
rect 273868 295718 273930 295954
rect 274166 295718 274250 295954
rect 274486 295718 274570 295954
rect 274806 295718 274868 295954
rect 273868 295634 274868 295718
rect 273868 295398 273930 295634
rect 274166 295398 274250 295634
rect 274486 295398 274570 295634
rect 274806 295398 274868 295634
rect 273868 295366 274868 295398
rect 23868 291454 24868 291486
rect 23868 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 24868 291454
rect 23868 291134 24868 291218
rect 23868 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 24868 291134
rect 23868 290866 24868 290898
rect 43868 291454 44868 291486
rect 43868 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 44868 291454
rect 43868 291134 44868 291218
rect 43868 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 44868 291134
rect 43868 290866 44868 290898
rect 63868 291454 64868 291486
rect 63868 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 64868 291454
rect 63868 291134 64868 291218
rect 63868 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 64868 291134
rect 63868 290866 64868 290898
rect 83868 291454 84868 291486
rect 83868 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 84868 291454
rect 83868 291134 84868 291218
rect 83868 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 84868 291134
rect 83868 290866 84868 290898
rect 103868 291454 104868 291486
rect 103868 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 104868 291454
rect 103868 291134 104868 291218
rect 103868 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 104868 291134
rect 103868 290866 104868 290898
rect 123868 291454 124868 291486
rect 123868 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 124868 291454
rect 123868 291134 124868 291218
rect 123868 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 124868 291134
rect 123868 290866 124868 290898
rect 143868 291454 144868 291486
rect 143868 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 144868 291454
rect 143868 291134 144868 291218
rect 143868 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 144868 291134
rect 143868 290866 144868 290898
rect 163868 291454 164868 291486
rect 163868 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 164868 291454
rect 163868 291134 164868 291218
rect 163868 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 164868 291134
rect 163868 290866 164868 290898
rect 183868 291454 184868 291486
rect 183868 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 184868 291454
rect 183868 291134 184868 291218
rect 183868 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 184868 291134
rect 183868 290866 184868 290898
rect 203868 291454 204868 291486
rect 203868 291218 203930 291454
rect 204166 291218 204250 291454
rect 204486 291218 204570 291454
rect 204806 291218 204868 291454
rect 203868 291134 204868 291218
rect 203868 290898 203930 291134
rect 204166 290898 204250 291134
rect 204486 290898 204570 291134
rect 204806 290898 204868 291134
rect 203868 290866 204868 290898
rect 223868 291454 224868 291486
rect 223868 291218 223930 291454
rect 224166 291218 224250 291454
rect 224486 291218 224570 291454
rect 224806 291218 224868 291454
rect 223868 291134 224868 291218
rect 223868 290898 223930 291134
rect 224166 290898 224250 291134
rect 224486 290898 224570 291134
rect 224806 290898 224868 291134
rect 223868 290866 224868 290898
rect 243868 291454 244868 291486
rect 243868 291218 243930 291454
rect 244166 291218 244250 291454
rect 244486 291218 244570 291454
rect 244806 291218 244868 291454
rect 243868 291134 244868 291218
rect 243868 290898 243930 291134
rect 244166 290898 244250 291134
rect 244486 290898 244570 291134
rect 244806 290898 244868 291134
rect 243868 290866 244868 290898
rect 263868 291454 264868 291486
rect 263868 291218 263930 291454
rect 264166 291218 264250 291454
rect 264486 291218 264570 291454
rect 264806 291218 264868 291454
rect 263868 291134 264868 291218
rect 263868 290898 263930 291134
rect 264166 290898 264250 291134
rect 264486 290898 264570 291134
rect 264806 290898 264868 291134
rect 263868 290866 264868 290898
rect 283868 291454 284868 291486
rect 283868 291218 283930 291454
rect 284166 291218 284250 291454
rect 284486 291218 284570 291454
rect 284806 291218 284868 291454
rect 283868 291134 284868 291218
rect 283868 290898 283930 291134
rect 284166 290898 284250 291134
rect 284486 290898 284570 291134
rect 284806 290898 284868 291134
rect 283868 290866 284868 290898
rect 33868 259954 34868 259986
rect 33868 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 34868 259954
rect 33868 259634 34868 259718
rect 33868 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 34868 259634
rect 33868 259366 34868 259398
rect 53868 259954 54868 259986
rect 53868 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 54868 259954
rect 53868 259634 54868 259718
rect 53868 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 54868 259634
rect 53868 259366 54868 259398
rect 73868 259954 74868 259986
rect 73868 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 74868 259954
rect 73868 259634 74868 259718
rect 73868 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 74868 259634
rect 73868 259366 74868 259398
rect 93868 259954 94868 259986
rect 93868 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 94868 259954
rect 93868 259634 94868 259718
rect 93868 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 94868 259634
rect 93868 259366 94868 259398
rect 113868 259954 114868 259986
rect 113868 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 114868 259954
rect 113868 259634 114868 259718
rect 113868 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 114868 259634
rect 113868 259366 114868 259398
rect 133868 259954 134868 259986
rect 133868 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 134868 259954
rect 133868 259634 134868 259718
rect 133868 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 134868 259634
rect 133868 259366 134868 259398
rect 153868 259954 154868 259986
rect 153868 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 154868 259954
rect 153868 259634 154868 259718
rect 153868 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 154868 259634
rect 153868 259366 154868 259398
rect 173868 259954 174868 259986
rect 173868 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 174868 259954
rect 173868 259634 174868 259718
rect 173868 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 174868 259634
rect 173868 259366 174868 259398
rect 193868 259954 194868 259986
rect 193868 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 194868 259954
rect 193868 259634 194868 259718
rect 193868 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 194868 259634
rect 193868 259366 194868 259398
rect 213868 259954 214868 259986
rect 213868 259718 213930 259954
rect 214166 259718 214250 259954
rect 214486 259718 214570 259954
rect 214806 259718 214868 259954
rect 213868 259634 214868 259718
rect 213868 259398 213930 259634
rect 214166 259398 214250 259634
rect 214486 259398 214570 259634
rect 214806 259398 214868 259634
rect 213868 259366 214868 259398
rect 233868 259954 234868 259986
rect 233868 259718 233930 259954
rect 234166 259718 234250 259954
rect 234486 259718 234570 259954
rect 234806 259718 234868 259954
rect 233868 259634 234868 259718
rect 233868 259398 233930 259634
rect 234166 259398 234250 259634
rect 234486 259398 234570 259634
rect 234806 259398 234868 259634
rect 233868 259366 234868 259398
rect 253868 259954 254868 259986
rect 253868 259718 253930 259954
rect 254166 259718 254250 259954
rect 254486 259718 254570 259954
rect 254806 259718 254868 259954
rect 253868 259634 254868 259718
rect 253868 259398 253930 259634
rect 254166 259398 254250 259634
rect 254486 259398 254570 259634
rect 254806 259398 254868 259634
rect 253868 259366 254868 259398
rect 273868 259954 274868 259986
rect 273868 259718 273930 259954
rect 274166 259718 274250 259954
rect 274486 259718 274570 259954
rect 274806 259718 274868 259954
rect 273868 259634 274868 259718
rect 273868 259398 273930 259634
rect 274166 259398 274250 259634
rect 274486 259398 274570 259634
rect 274806 259398 274868 259634
rect 273868 259366 274868 259398
rect 23868 255454 24868 255486
rect 23868 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 24868 255454
rect 23868 255134 24868 255218
rect 23868 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 24868 255134
rect 23868 254866 24868 254898
rect 43868 255454 44868 255486
rect 43868 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 44868 255454
rect 43868 255134 44868 255218
rect 43868 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 44868 255134
rect 43868 254866 44868 254898
rect 63868 255454 64868 255486
rect 63868 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 64868 255454
rect 63868 255134 64868 255218
rect 63868 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 64868 255134
rect 63868 254866 64868 254898
rect 83868 255454 84868 255486
rect 83868 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 84868 255454
rect 83868 255134 84868 255218
rect 83868 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 84868 255134
rect 83868 254866 84868 254898
rect 103868 255454 104868 255486
rect 103868 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 104868 255454
rect 103868 255134 104868 255218
rect 103868 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 104868 255134
rect 103868 254866 104868 254898
rect 123868 255454 124868 255486
rect 123868 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 124868 255454
rect 123868 255134 124868 255218
rect 123868 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 124868 255134
rect 123868 254866 124868 254898
rect 143868 255454 144868 255486
rect 143868 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 144868 255454
rect 143868 255134 144868 255218
rect 143868 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 144868 255134
rect 143868 254866 144868 254898
rect 163868 255454 164868 255486
rect 163868 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 164868 255454
rect 163868 255134 164868 255218
rect 163868 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 164868 255134
rect 163868 254866 164868 254898
rect 183868 255454 184868 255486
rect 183868 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 184868 255454
rect 183868 255134 184868 255218
rect 183868 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 184868 255134
rect 183868 254866 184868 254898
rect 203868 255454 204868 255486
rect 203868 255218 203930 255454
rect 204166 255218 204250 255454
rect 204486 255218 204570 255454
rect 204806 255218 204868 255454
rect 203868 255134 204868 255218
rect 203868 254898 203930 255134
rect 204166 254898 204250 255134
rect 204486 254898 204570 255134
rect 204806 254898 204868 255134
rect 203868 254866 204868 254898
rect 223868 255454 224868 255486
rect 223868 255218 223930 255454
rect 224166 255218 224250 255454
rect 224486 255218 224570 255454
rect 224806 255218 224868 255454
rect 223868 255134 224868 255218
rect 223868 254898 223930 255134
rect 224166 254898 224250 255134
rect 224486 254898 224570 255134
rect 224806 254898 224868 255134
rect 223868 254866 224868 254898
rect 243868 255454 244868 255486
rect 243868 255218 243930 255454
rect 244166 255218 244250 255454
rect 244486 255218 244570 255454
rect 244806 255218 244868 255454
rect 243868 255134 244868 255218
rect 243868 254898 243930 255134
rect 244166 254898 244250 255134
rect 244486 254898 244570 255134
rect 244806 254898 244868 255134
rect 243868 254866 244868 254898
rect 263868 255454 264868 255486
rect 263868 255218 263930 255454
rect 264166 255218 264250 255454
rect 264486 255218 264570 255454
rect 264806 255218 264868 255454
rect 263868 255134 264868 255218
rect 263868 254898 263930 255134
rect 264166 254898 264250 255134
rect 264486 254898 264570 255134
rect 264806 254898 264868 255134
rect 263868 254866 264868 254898
rect 283868 255454 284868 255486
rect 283868 255218 283930 255454
rect 284166 255218 284250 255454
rect 284486 255218 284570 255454
rect 284806 255218 284868 255454
rect 283868 255134 284868 255218
rect 283868 254898 283930 255134
rect 284166 254898 284250 255134
rect 284486 254898 284570 255134
rect 284806 254898 284868 255134
rect 283868 254866 284868 254898
rect 33868 223954 34868 223986
rect 33868 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 34868 223954
rect 33868 223634 34868 223718
rect 33868 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 34868 223634
rect 33868 223366 34868 223398
rect 53868 223954 54868 223986
rect 53868 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 54868 223954
rect 53868 223634 54868 223718
rect 53868 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 54868 223634
rect 53868 223366 54868 223398
rect 73868 223954 74868 223986
rect 73868 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 74868 223954
rect 73868 223634 74868 223718
rect 73868 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 74868 223634
rect 73868 223366 74868 223398
rect 93868 223954 94868 223986
rect 93868 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 94868 223954
rect 93868 223634 94868 223718
rect 93868 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 94868 223634
rect 93868 223366 94868 223398
rect 113868 223954 114868 223986
rect 113868 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 114868 223954
rect 113868 223634 114868 223718
rect 113868 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 114868 223634
rect 113868 223366 114868 223398
rect 133868 223954 134868 223986
rect 133868 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 134868 223954
rect 133868 223634 134868 223718
rect 133868 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 134868 223634
rect 133868 223366 134868 223398
rect 153868 223954 154868 223986
rect 153868 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 154868 223954
rect 153868 223634 154868 223718
rect 153868 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 154868 223634
rect 153868 223366 154868 223398
rect 173868 223954 174868 223986
rect 173868 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 174868 223954
rect 173868 223634 174868 223718
rect 173868 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 174868 223634
rect 173868 223366 174868 223398
rect 193868 223954 194868 223986
rect 193868 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 194868 223954
rect 193868 223634 194868 223718
rect 193868 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 194868 223634
rect 193868 223366 194868 223398
rect 213868 223954 214868 223986
rect 213868 223718 213930 223954
rect 214166 223718 214250 223954
rect 214486 223718 214570 223954
rect 214806 223718 214868 223954
rect 213868 223634 214868 223718
rect 213868 223398 213930 223634
rect 214166 223398 214250 223634
rect 214486 223398 214570 223634
rect 214806 223398 214868 223634
rect 213868 223366 214868 223398
rect 233868 223954 234868 223986
rect 233868 223718 233930 223954
rect 234166 223718 234250 223954
rect 234486 223718 234570 223954
rect 234806 223718 234868 223954
rect 233868 223634 234868 223718
rect 233868 223398 233930 223634
rect 234166 223398 234250 223634
rect 234486 223398 234570 223634
rect 234806 223398 234868 223634
rect 233868 223366 234868 223398
rect 253868 223954 254868 223986
rect 253868 223718 253930 223954
rect 254166 223718 254250 223954
rect 254486 223718 254570 223954
rect 254806 223718 254868 223954
rect 253868 223634 254868 223718
rect 253868 223398 253930 223634
rect 254166 223398 254250 223634
rect 254486 223398 254570 223634
rect 254806 223398 254868 223634
rect 253868 223366 254868 223398
rect 273868 223954 274868 223986
rect 273868 223718 273930 223954
rect 274166 223718 274250 223954
rect 274486 223718 274570 223954
rect 274806 223718 274868 223954
rect 273868 223634 274868 223718
rect 273868 223398 273930 223634
rect 274166 223398 274250 223634
rect 274486 223398 274570 223634
rect 274806 223398 274868 223634
rect 273868 223366 274868 223398
rect 23868 219454 24868 219486
rect 23868 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 24868 219454
rect 23868 219134 24868 219218
rect 23868 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 24868 219134
rect 23868 218866 24868 218898
rect 43868 219454 44868 219486
rect 43868 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 44868 219454
rect 43868 219134 44868 219218
rect 43868 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 44868 219134
rect 43868 218866 44868 218898
rect 63868 219454 64868 219486
rect 63868 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 64868 219454
rect 63868 219134 64868 219218
rect 63868 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 64868 219134
rect 63868 218866 64868 218898
rect 83868 219454 84868 219486
rect 83868 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 84868 219454
rect 83868 219134 84868 219218
rect 83868 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 84868 219134
rect 83868 218866 84868 218898
rect 103868 219454 104868 219486
rect 103868 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 104868 219454
rect 103868 219134 104868 219218
rect 103868 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 104868 219134
rect 103868 218866 104868 218898
rect 123868 219454 124868 219486
rect 123868 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 124868 219454
rect 123868 219134 124868 219218
rect 123868 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 124868 219134
rect 123868 218866 124868 218898
rect 143868 219454 144868 219486
rect 143868 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 144868 219454
rect 143868 219134 144868 219218
rect 143868 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 144868 219134
rect 143868 218866 144868 218898
rect 163868 219454 164868 219486
rect 163868 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 164868 219454
rect 163868 219134 164868 219218
rect 163868 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 164868 219134
rect 163868 218866 164868 218898
rect 183868 219454 184868 219486
rect 183868 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 184868 219454
rect 183868 219134 184868 219218
rect 183868 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 184868 219134
rect 183868 218866 184868 218898
rect 203868 219454 204868 219486
rect 203868 219218 203930 219454
rect 204166 219218 204250 219454
rect 204486 219218 204570 219454
rect 204806 219218 204868 219454
rect 203868 219134 204868 219218
rect 203868 218898 203930 219134
rect 204166 218898 204250 219134
rect 204486 218898 204570 219134
rect 204806 218898 204868 219134
rect 203868 218866 204868 218898
rect 223868 219454 224868 219486
rect 223868 219218 223930 219454
rect 224166 219218 224250 219454
rect 224486 219218 224570 219454
rect 224806 219218 224868 219454
rect 223868 219134 224868 219218
rect 223868 218898 223930 219134
rect 224166 218898 224250 219134
rect 224486 218898 224570 219134
rect 224806 218898 224868 219134
rect 223868 218866 224868 218898
rect 243868 219454 244868 219486
rect 243868 219218 243930 219454
rect 244166 219218 244250 219454
rect 244486 219218 244570 219454
rect 244806 219218 244868 219454
rect 243868 219134 244868 219218
rect 243868 218898 243930 219134
rect 244166 218898 244250 219134
rect 244486 218898 244570 219134
rect 244806 218898 244868 219134
rect 243868 218866 244868 218898
rect 263868 219454 264868 219486
rect 263868 219218 263930 219454
rect 264166 219218 264250 219454
rect 264486 219218 264570 219454
rect 264806 219218 264868 219454
rect 263868 219134 264868 219218
rect 263868 218898 263930 219134
rect 264166 218898 264250 219134
rect 264486 218898 264570 219134
rect 264806 218898 264868 219134
rect 263868 218866 264868 218898
rect 283868 219454 284868 219486
rect 283868 219218 283930 219454
rect 284166 219218 284250 219454
rect 284486 219218 284570 219454
rect 284806 219218 284868 219454
rect 283868 219134 284868 219218
rect 283868 218898 283930 219134
rect 284166 218898 284250 219134
rect 284486 218898 284570 219134
rect 284806 218898 284868 219134
rect 283868 218866 284868 218898
rect 22691 202876 22757 202877
rect 22691 202812 22692 202876
rect 22756 202812 22757 202876
rect 22691 202811 22757 202812
rect 22694 200130 22754 202811
rect 22694 200070 23306 200130
rect 21955 75852 22021 75853
rect 21955 75788 21956 75852
rect 22020 75788 22021 75852
rect 21955 75787 22021 75788
rect 23246 74357 23306 200070
rect 23868 183454 24868 183486
rect 23868 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 24868 183454
rect 23868 183134 24868 183218
rect 23868 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 24868 183134
rect 23868 182866 24868 182898
rect 43868 183454 44868 183486
rect 43868 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 44868 183454
rect 43868 183134 44868 183218
rect 43868 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 44868 183134
rect 43868 182866 44868 182898
rect 63868 183454 64868 183486
rect 63868 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 64868 183454
rect 63868 183134 64868 183218
rect 63868 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 64868 183134
rect 63868 182866 64868 182898
rect 83868 183454 84868 183486
rect 83868 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 84868 183454
rect 83868 183134 84868 183218
rect 83868 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 84868 183134
rect 83868 182866 84868 182898
rect 103868 183454 104868 183486
rect 103868 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 104868 183454
rect 103868 183134 104868 183218
rect 103868 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 104868 183134
rect 103868 182866 104868 182898
rect 123868 183454 124868 183486
rect 123868 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 124868 183454
rect 123868 183134 124868 183218
rect 123868 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 124868 183134
rect 123868 182866 124868 182898
rect 143868 183454 144868 183486
rect 143868 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 144868 183454
rect 143868 183134 144868 183218
rect 143868 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 144868 183134
rect 143868 182866 144868 182898
rect 163868 183454 164868 183486
rect 163868 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 164868 183454
rect 163868 183134 164868 183218
rect 163868 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 164868 183134
rect 163868 182866 164868 182898
rect 183868 183454 184868 183486
rect 183868 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 184868 183454
rect 183868 183134 184868 183218
rect 183868 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 184868 183134
rect 183868 182866 184868 182898
rect 203868 183454 204868 183486
rect 203868 183218 203930 183454
rect 204166 183218 204250 183454
rect 204486 183218 204570 183454
rect 204806 183218 204868 183454
rect 203868 183134 204868 183218
rect 203868 182898 203930 183134
rect 204166 182898 204250 183134
rect 204486 182898 204570 183134
rect 204806 182898 204868 183134
rect 203868 182866 204868 182898
rect 223868 183454 224868 183486
rect 223868 183218 223930 183454
rect 224166 183218 224250 183454
rect 224486 183218 224570 183454
rect 224806 183218 224868 183454
rect 223868 183134 224868 183218
rect 223868 182898 223930 183134
rect 224166 182898 224250 183134
rect 224486 182898 224570 183134
rect 224806 182898 224868 183134
rect 223868 182866 224868 182898
rect 243868 183454 244868 183486
rect 243868 183218 243930 183454
rect 244166 183218 244250 183454
rect 244486 183218 244570 183454
rect 244806 183218 244868 183454
rect 243868 183134 244868 183218
rect 243868 182898 243930 183134
rect 244166 182898 244250 183134
rect 244486 182898 244570 183134
rect 244806 182898 244868 183134
rect 243868 182866 244868 182898
rect 263868 183454 264868 183486
rect 263868 183218 263930 183454
rect 264166 183218 264250 183454
rect 264486 183218 264570 183454
rect 264806 183218 264868 183454
rect 263868 183134 264868 183218
rect 263868 182898 263930 183134
rect 264166 182898 264250 183134
rect 264486 182898 264570 183134
rect 264806 182898 264868 183134
rect 263868 182866 264868 182898
rect 283868 183454 284868 183486
rect 283868 183218 283930 183454
rect 284166 183218 284250 183454
rect 284486 183218 284570 183454
rect 284806 183218 284868 183454
rect 283868 183134 284868 183218
rect 283868 182898 283930 183134
rect 284166 182898 284250 183134
rect 284486 182898 284570 183134
rect 284806 182898 284868 183134
rect 283868 182866 284868 182898
rect 33868 151954 34868 151986
rect 33868 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 34868 151954
rect 33868 151634 34868 151718
rect 33868 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 34868 151634
rect 33868 151366 34868 151398
rect 53868 151954 54868 151986
rect 53868 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 54868 151954
rect 53868 151634 54868 151718
rect 53868 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 54868 151634
rect 53868 151366 54868 151398
rect 73868 151954 74868 151986
rect 73868 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 74868 151954
rect 73868 151634 74868 151718
rect 73868 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 74868 151634
rect 73868 151366 74868 151398
rect 93868 151954 94868 151986
rect 93868 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 94868 151954
rect 93868 151634 94868 151718
rect 93868 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 94868 151634
rect 93868 151366 94868 151398
rect 113868 151954 114868 151986
rect 113868 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 114868 151954
rect 113868 151634 114868 151718
rect 113868 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 114868 151634
rect 113868 151366 114868 151398
rect 133868 151954 134868 151986
rect 133868 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 134868 151954
rect 133868 151634 134868 151718
rect 133868 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 134868 151634
rect 133868 151366 134868 151398
rect 153868 151954 154868 151986
rect 153868 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 154868 151954
rect 153868 151634 154868 151718
rect 153868 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 154868 151634
rect 153868 151366 154868 151398
rect 173868 151954 174868 151986
rect 173868 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 174868 151954
rect 173868 151634 174868 151718
rect 173868 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 174868 151634
rect 173868 151366 174868 151398
rect 193868 151954 194868 151986
rect 193868 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 194868 151954
rect 193868 151634 194868 151718
rect 193868 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 194868 151634
rect 193868 151366 194868 151398
rect 213868 151954 214868 151986
rect 213868 151718 213930 151954
rect 214166 151718 214250 151954
rect 214486 151718 214570 151954
rect 214806 151718 214868 151954
rect 213868 151634 214868 151718
rect 213868 151398 213930 151634
rect 214166 151398 214250 151634
rect 214486 151398 214570 151634
rect 214806 151398 214868 151634
rect 213868 151366 214868 151398
rect 233868 151954 234868 151986
rect 233868 151718 233930 151954
rect 234166 151718 234250 151954
rect 234486 151718 234570 151954
rect 234806 151718 234868 151954
rect 233868 151634 234868 151718
rect 233868 151398 233930 151634
rect 234166 151398 234250 151634
rect 234486 151398 234570 151634
rect 234806 151398 234868 151634
rect 233868 151366 234868 151398
rect 253868 151954 254868 151986
rect 253868 151718 253930 151954
rect 254166 151718 254250 151954
rect 254486 151718 254570 151954
rect 254806 151718 254868 151954
rect 253868 151634 254868 151718
rect 253868 151398 253930 151634
rect 254166 151398 254250 151634
rect 254486 151398 254570 151634
rect 254806 151398 254868 151634
rect 253868 151366 254868 151398
rect 273868 151954 274868 151986
rect 273868 151718 273930 151954
rect 274166 151718 274250 151954
rect 274486 151718 274570 151954
rect 274806 151718 274868 151954
rect 273868 151634 274868 151718
rect 273868 151398 273930 151634
rect 274166 151398 274250 151634
rect 274486 151398 274570 151634
rect 274806 151398 274868 151634
rect 273868 151366 274868 151398
rect 23868 147454 24868 147486
rect 23868 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 24868 147454
rect 23868 147134 24868 147218
rect 23868 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 24868 147134
rect 23868 146866 24868 146898
rect 43868 147454 44868 147486
rect 43868 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 44868 147454
rect 43868 147134 44868 147218
rect 43868 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 44868 147134
rect 43868 146866 44868 146898
rect 63868 147454 64868 147486
rect 63868 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 64868 147454
rect 63868 147134 64868 147218
rect 63868 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 64868 147134
rect 63868 146866 64868 146898
rect 83868 147454 84868 147486
rect 83868 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 84868 147454
rect 83868 147134 84868 147218
rect 83868 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 84868 147134
rect 83868 146866 84868 146898
rect 103868 147454 104868 147486
rect 103868 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 104868 147454
rect 103868 147134 104868 147218
rect 103868 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 104868 147134
rect 103868 146866 104868 146898
rect 123868 147454 124868 147486
rect 123868 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 124868 147454
rect 123868 147134 124868 147218
rect 123868 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 124868 147134
rect 123868 146866 124868 146898
rect 143868 147454 144868 147486
rect 143868 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 144868 147454
rect 143868 147134 144868 147218
rect 143868 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 144868 147134
rect 143868 146866 144868 146898
rect 163868 147454 164868 147486
rect 163868 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 164868 147454
rect 163868 147134 164868 147218
rect 163868 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 164868 147134
rect 163868 146866 164868 146898
rect 183868 147454 184868 147486
rect 183868 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 184868 147454
rect 183868 147134 184868 147218
rect 183868 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 184868 147134
rect 183868 146866 184868 146898
rect 203868 147454 204868 147486
rect 203868 147218 203930 147454
rect 204166 147218 204250 147454
rect 204486 147218 204570 147454
rect 204806 147218 204868 147454
rect 203868 147134 204868 147218
rect 203868 146898 203930 147134
rect 204166 146898 204250 147134
rect 204486 146898 204570 147134
rect 204806 146898 204868 147134
rect 203868 146866 204868 146898
rect 223868 147454 224868 147486
rect 223868 147218 223930 147454
rect 224166 147218 224250 147454
rect 224486 147218 224570 147454
rect 224806 147218 224868 147454
rect 223868 147134 224868 147218
rect 223868 146898 223930 147134
rect 224166 146898 224250 147134
rect 224486 146898 224570 147134
rect 224806 146898 224868 147134
rect 223868 146866 224868 146898
rect 243868 147454 244868 147486
rect 243868 147218 243930 147454
rect 244166 147218 244250 147454
rect 244486 147218 244570 147454
rect 244806 147218 244868 147454
rect 243868 147134 244868 147218
rect 243868 146898 243930 147134
rect 244166 146898 244250 147134
rect 244486 146898 244570 147134
rect 244806 146898 244868 147134
rect 243868 146866 244868 146898
rect 263868 147454 264868 147486
rect 263868 147218 263930 147454
rect 264166 147218 264250 147454
rect 264486 147218 264570 147454
rect 264806 147218 264868 147454
rect 263868 147134 264868 147218
rect 263868 146898 263930 147134
rect 264166 146898 264250 147134
rect 264486 146898 264570 147134
rect 264806 146898 264868 147134
rect 263868 146866 264868 146898
rect 283868 147454 284868 147486
rect 283868 147218 283930 147454
rect 284166 147218 284250 147454
rect 284486 147218 284570 147454
rect 284806 147218 284868 147454
rect 283868 147134 284868 147218
rect 283868 146898 283930 147134
rect 284166 146898 284250 147134
rect 284486 146898 284570 147134
rect 284806 146898 284868 147134
rect 283868 146866 284868 146898
rect 33868 115954 34868 115986
rect 33868 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 34868 115954
rect 33868 115634 34868 115718
rect 33868 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 34868 115634
rect 33868 115366 34868 115398
rect 53868 115954 54868 115986
rect 53868 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 54868 115954
rect 53868 115634 54868 115718
rect 53868 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 54868 115634
rect 53868 115366 54868 115398
rect 73868 115954 74868 115986
rect 73868 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 74868 115954
rect 73868 115634 74868 115718
rect 73868 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 74868 115634
rect 73868 115366 74868 115398
rect 93868 115954 94868 115986
rect 93868 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 94868 115954
rect 93868 115634 94868 115718
rect 93868 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 94868 115634
rect 93868 115366 94868 115398
rect 113868 115954 114868 115986
rect 113868 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 114868 115954
rect 113868 115634 114868 115718
rect 113868 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 114868 115634
rect 113868 115366 114868 115398
rect 133868 115954 134868 115986
rect 133868 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 134868 115954
rect 133868 115634 134868 115718
rect 133868 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 134868 115634
rect 133868 115366 134868 115398
rect 153868 115954 154868 115986
rect 153868 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 154868 115954
rect 153868 115634 154868 115718
rect 153868 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 154868 115634
rect 153868 115366 154868 115398
rect 173868 115954 174868 115986
rect 173868 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 174868 115954
rect 173868 115634 174868 115718
rect 173868 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 174868 115634
rect 173868 115366 174868 115398
rect 193868 115954 194868 115986
rect 193868 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 194868 115954
rect 193868 115634 194868 115718
rect 193868 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 194868 115634
rect 193868 115366 194868 115398
rect 213868 115954 214868 115986
rect 213868 115718 213930 115954
rect 214166 115718 214250 115954
rect 214486 115718 214570 115954
rect 214806 115718 214868 115954
rect 213868 115634 214868 115718
rect 213868 115398 213930 115634
rect 214166 115398 214250 115634
rect 214486 115398 214570 115634
rect 214806 115398 214868 115634
rect 213868 115366 214868 115398
rect 233868 115954 234868 115986
rect 233868 115718 233930 115954
rect 234166 115718 234250 115954
rect 234486 115718 234570 115954
rect 234806 115718 234868 115954
rect 233868 115634 234868 115718
rect 233868 115398 233930 115634
rect 234166 115398 234250 115634
rect 234486 115398 234570 115634
rect 234806 115398 234868 115634
rect 233868 115366 234868 115398
rect 253868 115954 254868 115986
rect 253868 115718 253930 115954
rect 254166 115718 254250 115954
rect 254486 115718 254570 115954
rect 254806 115718 254868 115954
rect 253868 115634 254868 115718
rect 253868 115398 253930 115634
rect 254166 115398 254250 115634
rect 254486 115398 254570 115634
rect 254806 115398 254868 115634
rect 253868 115366 254868 115398
rect 273868 115954 274868 115986
rect 273868 115718 273930 115954
rect 274166 115718 274250 115954
rect 274486 115718 274570 115954
rect 274806 115718 274868 115954
rect 273868 115634 274868 115718
rect 273868 115398 273930 115634
rect 274166 115398 274250 115634
rect 274486 115398 274570 115634
rect 274806 115398 274868 115634
rect 273868 115366 274868 115398
rect 23868 111454 24868 111486
rect 23868 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 24868 111454
rect 23868 111134 24868 111218
rect 23868 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 24868 111134
rect 23868 110866 24868 110898
rect 43868 111454 44868 111486
rect 43868 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 44868 111454
rect 43868 111134 44868 111218
rect 43868 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 44868 111134
rect 43868 110866 44868 110898
rect 63868 111454 64868 111486
rect 63868 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 64868 111454
rect 63868 111134 64868 111218
rect 63868 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 64868 111134
rect 63868 110866 64868 110898
rect 83868 111454 84868 111486
rect 83868 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 84868 111454
rect 83868 111134 84868 111218
rect 83868 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 84868 111134
rect 83868 110866 84868 110898
rect 103868 111454 104868 111486
rect 103868 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 104868 111454
rect 103868 111134 104868 111218
rect 103868 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 104868 111134
rect 103868 110866 104868 110898
rect 123868 111454 124868 111486
rect 123868 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 124868 111454
rect 123868 111134 124868 111218
rect 123868 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 124868 111134
rect 123868 110866 124868 110898
rect 143868 111454 144868 111486
rect 143868 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 144868 111454
rect 143868 111134 144868 111218
rect 143868 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 144868 111134
rect 143868 110866 144868 110898
rect 163868 111454 164868 111486
rect 163868 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 164868 111454
rect 163868 111134 164868 111218
rect 163868 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 164868 111134
rect 163868 110866 164868 110898
rect 183868 111454 184868 111486
rect 183868 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 184868 111454
rect 183868 111134 184868 111218
rect 183868 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 184868 111134
rect 183868 110866 184868 110898
rect 203868 111454 204868 111486
rect 203868 111218 203930 111454
rect 204166 111218 204250 111454
rect 204486 111218 204570 111454
rect 204806 111218 204868 111454
rect 203868 111134 204868 111218
rect 203868 110898 203930 111134
rect 204166 110898 204250 111134
rect 204486 110898 204570 111134
rect 204806 110898 204868 111134
rect 203868 110866 204868 110898
rect 223868 111454 224868 111486
rect 223868 111218 223930 111454
rect 224166 111218 224250 111454
rect 224486 111218 224570 111454
rect 224806 111218 224868 111454
rect 223868 111134 224868 111218
rect 223868 110898 223930 111134
rect 224166 110898 224250 111134
rect 224486 110898 224570 111134
rect 224806 110898 224868 111134
rect 223868 110866 224868 110898
rect 243868 111454 244868 111486
rect 243868 111218 243930 111454
rect 244166 111218 244250 111454
rect 244486 111218 244570 111454
rect 244806 111218 244868 111454
rect 243868 111134 244868 111218
rect 243868 110898 243930 111134
rect 244166 110898 244250 111134
rect 244486 110898 244570 111134
rect 244806 110898 244868 111134
rect 243868 110866 244868 110898
rect 263868 111454 264868 111486
rect 263868 111218 263930 111454
rect 264166 111218 264250 111454
rect 264486 111218 264570 111454
rect 264806 111218 264868 111454
rect 263868 111134 264868 111218
rect 263868 110898 263930 111134
rect 264166 110898 264250 111134
rect 264486 110898 264570 111134
rect 264806 110898 264868 111134
rect 263868 110866 264868 110898
rect 283868 111454 284868 111486
rect 283868 111218 283930 111454
rect 284166 111218 284250 111454
rect 284486 111218 284570 111454
rect 284806 111218 284868 111454
rect 283868 111134 284868 111218
rect 283868 110898 283930 111134
rect 284166 110898 284250 111134
rect 284486 110898 284570 111134
rect 284806 110898 284868 111134
rect 283868 110866 284868 110898
rect 23611 80204 23677 80205
rect 23611 80140 23612 80204
rect 23676 80140 23677 80204
rect 23611 80139 23677 80140
rect 23614 74493 23674 80139
rect 23611 74492 23677 74493
rect 23611 74428 23612 74492
rect 23676 74428 23677 74492
rect 23611 74427 23677 74428
rect 23243 74356 23309 74357
rect 23243 74292 23244 74356
rect 23308 74292 23309 74356
rect 23243 74291 23309 74292
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19563 21860 19629 21861
rect 19563 21796 19564 21860
rect 19628 21796 19629 21860
rect 19563 21795 19629 21796
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 61954 24914 76000
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 66454 29414 76000
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 70954 33914 76000
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 75454 38414 76000
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 43954 42914 76000
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 48454 47414 76000
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 52954 51914 76000
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 76000
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 105294 70954 105914 76000
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 79568 43954 79888 43986
rect 79568 43718 79610 43954
rect 79846 43718 79888 43954
rect 79568 43634 79888 43718
rect 79568 43398 79610 43634
rect 79846 43398 79888 43634
rect 79568 43366 79888 43398
rect 64208 39454 64528 39486
rect 64208 39218 64250 39454
rect 64486 39218 64528 39454
rect 64208 39134 64528 39218
rect 64208 38898 64250 39134
rect 64486 38898 64528 39134
rect 64208 38866 64528 38898
rect 94928 39454 95248 39486
rect 94928 39218 94970 39454
rect 95206 39218 95248 39454
rect 94928 39134 95248 39218
rect 94928 38898 94970 39134
rect 95206 38898 95248 39134
rect 94928 38866 95248 38898
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 73794 3454 74414 22000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 7954 78914 22000
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 12454 83414 22000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 16954 87914 22000
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 21454 92414 22000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 76000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 76000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 76000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 76000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 76000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 76000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 76000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 76000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 76000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 76000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 76000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 76000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 76000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 76000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 76000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 76000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 76000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 76000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 76000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 76000
rect 286182 57221 286242 444891
rect 287654 345030 287714 457811
rect 287654 344970 288266 345030
rect 288206 332485 288266 344970
rect 288203 332484 288269 332485
rect 288203 332420 288204 332484
rect 288268 332420 288269 332484
rect 288203 332419 288269 332420
rect 287099 203556 287165 203557
rect 287099 203492 287100 203556
rect 287164 203492 287165 203556
rect 287099 203491 287165 203492
rect 287102 60077 287162 203491
rect 288206 202877 288266 332419
rect 287283 202876 287349 202877
rect 287283 202812 287284 202876
rect 287348 202812 287349 202876
rect 287283 202811 287349 202812
rect 288203 202876 288269 202877
rect 288203 202812 288204 202876
rect 288268 202812 288269 202876
rect 288203 202811 288269 202812
rect 287286 77893 287346 202811
rect 287283 77892 287349 77893
rect 287283 77828 287284 77892
rect 287348 77828 287349 77892
rect 287283 77827 287349 77828
rect 287099 60076 287165 60077
rect 287099 60012 287100 60076
rect 287164 60012 287165 60076
rect 287099 60011 287165 60012
rect 288390 57493 288450 585651
rect 291147 458964 291213 458965
rect 291147 458900 291148 458964
rect 291212 458900 291213 458964
rect 291147 458899 291213 458900
rect 289859 458828 289925 458829
rect 289859 458764 289860 458828
rect 289924 458764 289925 458828
rect 289859 458763 289925 458764
rect 288387 57492 288453 57493
rect 288387 57428 288388 57492
rect 288452 57428 288453 57492
rect 288387 57427 288453 57428
rect 289862 57357 289922 458763
rect 291150 60213 291210 458899
rect 291702 78029 291762 585651
rect 291699 78028 291765 78029
rect 291699 77964 291700 78028
rect 291764 77964 291765 78028
rect 291699 77963 291765 77964
rect 291147 60212 291213 60213
rect 291147 60148 291148 60212
rect 291212 60148 291213 60212
rect 291147 60147 291213 60148
rect 292622 59941 292682 586331
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 292619 59940 292685 59941
rect 292619 59876 292620 59940
rect 292684 59876 292685 59940
rect 292619 59875 292685 59876
rect 289859 57356 289925 57357
rect 289859 57292 289860 57356
rect 289924 57292 289925 57356
rect 289859 57291 289925 57292
rect 286179 57220 286245 57221
rect 286179 57156 286180 57220
rect 286244 57156 286245 57220
rect 286179 57155 286245 57156
rect 294294 56000 294914 79398
rect 295934 54501 295994 700299
rect 303294 700000 303914 700398
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 700000 339914 700398
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 700000 375914 700398
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 700000 411914 700398
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 700000 447914 700398
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 700000 483914 700398
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 700000 519914 700398
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 700000 555914 700398
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 313868 691954 314868 691986
rect 313868 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 314868 691954
rect 313868 691634 314868 691718
rect 313868 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 314868 691634
rect 313868 691366 314868 691398
rect 333868 691954 334868 691986
rect 333868 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 334868 691954
rect 333868 691634 334868 691718
rect 333868 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 334868 691634
rect 333868 691366 334868 691398
rect 353868 691954 354868 691986
rect 353868 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 354868 691954
rect 353868 691634 354868 691718
rect 353868 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 354868 691634
rect 353868 691366 354868 691398
rect 373868 691954 374868 691986
rect 373868 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 374868 691954
rect 373868 691634 374868 691718
rect 373868 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 374868 691634
rect 373868 691366 374868 691398
rect 393868 691954 394868 691986
rect 393868 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 394868 691954
rect 393868 691634 394868 691718
rect 393868 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 394868 691634
rect 393868 691366 394868 691398
rect 413868 691954 414868 691986
rect 413868 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 414868 691954
rect 413868 691634 414868 691718
rect 413868 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 414868 691634
rect 413868 691366 414868 691398
rect 433868 691954 434868 691986
rect 433868 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 434868 691954
rect 433868 691634 434868 691718
rect 433868 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 434868 691634
rect 433868 691366 434868 691398
rect 453868 691954 454868 691986
rect 453868 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 454868 691954
rect 453868 691634 454868 691718
rect 453868 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 454868 691634
rect 453868 691366 454868 691398
rect 473868 691954 474868 691986
rect 473868 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 474868 691954
rect 473868 691634 474868 691718
rect 473868 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 474868 691634
rect 473868 691366 474868 691398
rect 493868 691954 494868 691986
rect 493868 691718 493930 691954
rect 494166 691718 494250 691954
rect 494486 691718 494570 691954
rect 494806 691718 494868 691954
rect 493868 691634 494868 691718
rect 493868 691398 493930 691634
rect 494166 691398 494250 691634
rect 494486 691398 494570 691634
rect 494806 691398 494868 691634
rect 493868 691366 494868 691398
rect 513868 691954 514868 691986
rect 513868 691718 513930 691954
rect 514166 691718 514250 691954
rect 514486 691718 514570 691954
rect 514806 691718 514868 691954
rect 513868 691634 514868 691718
rect 513868 691398 513930 691634
rect 514166 691398 514250 691634
rect 514486 691398 514570 691634
rect 514806 691398 514868 691634
rect 513868 691366 514868 691398
rect 533868 691954 534868 691986
rect 533868 691718 533930 691954
rect 534166 691718 534250 691954
rect 534486 691718 534570 691954
rect 534806 691718 534868 691954
rect 533868 691634 534868 691718
rect 533868 691398 533930 691634
rect 534166 691398 534250 691634
rect 534486 691398 534570 691634
rect 534806 691398 534868 691634
rect 533868 691366 534868 691398
rect 553868 691954 554868 691986
rect 553868 691718 553930 691954
rect 554166 691718 554250 691954
rect 554486 691718 554570 691954
rect 554806 691718 554868 691954
rect 553868 691634 554868 691718
rect 553868 691398 553930 691634
rect 554166 691398 554250 691634
rect 554486 691398 554570 691634
rect 554806 691398 554868 691634
rect 553868 691366 554868 691398
rect 303868 687454 304868 687486
rect 303868 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 304868 687454
rect 303868 687134 304868 687218
rect 303868 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 304868 687134
rect 303868 686866 304868 686898
rect 323868 687454 324868 687486
rect 323868 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 324868 687454
rect 323868 687134 324868 687218
rect 323868 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 324868 687134
rect 323868 686866 324868 686898
rect 343868 687454 344868 687486
rect 343868 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 344868 687454
rect 343868 687134 344868 687218
rect 343868 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 344868 687134
rect 343868 686866 344868 686898
rect 363868 687454 364868 687486
rect 363868 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 364868 687454
rect 363868 687134 364868 687218
rect 363868 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 364868 687134
rect 363868 686866 364868 686898
rect 383868 687454 384868 687486
rect 383868 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 384868 687454
rect 383868 687134 384868 687218
rect 383868 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 384868 687134
rect 383868 686866 384868 686898
rect 403868 687454 404868 687486
rect 403868 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 404868 687454
rect 403868 687134 404868 687218
rect 403868 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 404868 687134
rect 403868 686866 404868 686898
rect 423868 687454 424868 687486
rect 423868 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 424868 687454
rect 423868 687134 424868 687218
rect 423868 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 424868 687134
rect 423868 686866 424868 686898
rect 443868 687454 444868 687486
rect 443868 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 444868 687454
rect 443868 687134 444868 687218
rect 443868 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 444868 687134
rect 443868 686866 444868 686898
rect 463868 687454 464868 687486
rect 463868 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 464868 687454
rect 463868 687134 464868 687218
rect 463868 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 464868 687134
rect 463868 686866 464868 686898
rect 483868 687454 484868 687486
rect 483868 687218 483930 687454
rect 484166 687218 484250 687454
rect 484486 687218 484570 687454
rect 484806 687218 484868 687454
rect 483868 687134 484868 687218
rect 483868 686898 483930 687134
rect 484166 686898 484250 687134
rect 484486 686898 484570 687134
rect 484806 686898 484868 687134
rect 483868 686866 484868 686898
rect 503868 687454 504868 687486
rect 503868 687218 503930 687454
rect 504166 687218 504250 687454
rect 504486 687218 504570 687454
rect 504806 687218 504868 687454
rect 503868 687134 504868 687218
rect 503868 686898 503930 687134
rect 504166 686898 504250 687134
rect 504486 686898 504570 687134
rect 504806 686898 504868 687134
rect 503868 686866 504868 686898
rect 523868 687454 524868 687486
rect 523868 687218 523930 687454
rect 524166 687218 524250 687454
rect 524486 687218 524570 687454
rect 524806 687218 524868 687454
rect 523868 687134 524868 687218
rect 523868 686898 523930 687134
rect 524166 686898 524250 687134
rect 524486 686898 524570 687134
rect 524806 686898 524868 687134
rect 523868 686866 524868 686898
rect 543868 687454 544868 687486
rect 543868 687218 543930 687454
rect 544166 687218 544250 687454
rect 544486 687218 544570 687454
rect 544806 687218 544868 687454
rect 543868 687134 544868 687218
rect 543868 686898 543930 687134
rect 544166 686898 544250 687134
rect 544486 686898 544570 687134
rect 544806 686898 544868 687134
rect 543868 686866 544868 686898
rect 563868 687454 564868 687486
rect 563868 687218 563930 687454
rect 564166 687218 564250 687454
rect 564486 687218 564570 687454
rect 564806 687218 564868 687454
rect 563868 687134 564868 687218
rect 563868 686898 563930 687134
rect 564166 686898 564250 687134
rect 564486 686898 564570 687134
rect 564806 686898 564868 687134
rect 563868 686866 564868 686898
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 313868 655954 314868 655986
rect 313868 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 314868 655954
rect 313868 655634 314868 655718
rect 313868 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 314868 655634
rect 313868 655366 314868 655398
rect 333868 655954 334868 655986
rect 333868 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 334868 655954
rect 333868 655634 334868 655718
rect 333868 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 334868 655634
rect 333868 655366 334868 655398
rect 353868 655954 354868 655986
rect 353868 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 354868 655954
rect 353868 655634 354868 655718
rect 353868 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 354868 655634
rect 353868 655366 354868 655398
rect 373868 655954 374868 655986
rect 373868 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 374868 655954
rect 373868 655634 374868 655718
rect 373868 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 374868 655634
rect 373868 655366 374868 655398
rect 393868 655954 394868 655986
rect 393868 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 394868 655954
rect 393868 655634 394868 655718
rect 393868 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 394868 655634
rect 393868 655366 394868 655398
rect 413868 655954 414868 655986
rect 413868 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 414868 655954
rect 413868 655634 414868 655718
rect 413868 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 414868 655634
rect 413868 655366 414868 655398
rect 433868 655954 434868 655986
rect 433868 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 434868 655954
rect 433868 655634 434868 655718
rect 433868 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 434868 655634
rect 433868 655366 434868 655398
rect 453868 655954 454868 655986
rect 453868 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 454868 655954
rect 453868 655634 454868 655718
rect 453868 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 454868 655634
rect 453868 655366 454868 655398
rect 473868 655954 474868 655986
rect 473868 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 474868 655954
rect 473868 655634 474868 655718
rect 473868 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 474868 655634
rect 473868 655366 474868 655398
rect 493868 655954 494868 655986
rect 493868 655718 493930 655954
rect 494166 655718 494250 655954
rect 494486 655718 494570 655954
rect 494806 655718 494868 655954
rect 493868 655634 494868 655718
rect 493868 655398 493930 655634
rect 494166 655398 494250 655634
rect 494486 655398 494570 655634
rect 494806 655398 494868 655634
rect 493868 655366 494868 655398
rect 513868 655954 514868 655986
rect 513868 655718 513930 655954
rect 514166 655718 514250 655954
rect 514486 655718 514570 655954
rect 514806 655718 514868 655954
rect 513868 655634 514868 655718
rect 513868 655398 513930 655634
rect 514166 655398 514250 655634
rect 514486 655398 514570 655634
rect 514806 655398 514868 655634
rect 513868 655366 514868 655398
rect 533868 655954 534868 655986
rect 533868 655718 533930 655954
rect 534166 655718 534250 655954
rect 534486 655718 534570 655954
rect 534806 655718 534868 655954
rect 533868 655634 534868 655718
rect 533868 655398 533930 655634
rect 534166 655398 534250 655634
rect 534486 655398 534570 655634
rect 534806 655398 534868 655634
rect 533868 655366 534868 655398
rect 553868 655954 554868 655986
rect 553868 655718 553930 655954
rect 554166 655718 554250 655954
rect 554486 655718 554570 655954
rect 554806 655718 554868 655954
rect 553868 655634 554868 655718
rect 553868 655398 553930 655634
rect 554166 655398 554250 655634
rect 554486 655398 554570 655634
rect 554806 655398 554868 655634
rect 553868 655366 554868 655398
rect 303868 651454 304868 651486
rect 303868 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 304868 651454
rect 303868 651134 304868 651218
rect 303868 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 304868 651134
rect 303868 650866 304868 650898
rect 323868 651454 324868 651486
rect 323868 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 324868 651454
rect 323868 651134 324868 651218
rect 323868 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 324868 651134
rect 323868 650866 324868 650898
rect 343868 651454 344868 651486
rect 343868 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 344868 651454
rect 343868 651134 344868 651218
rect 343868 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 344868 651134
rect 343868 650866 344868 650898
rect 363868 651454 364868 651486
rect 363868 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 364868 651454
rect 363868 651134 364868 651218
rect 363868 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 364868 651134
rect 363868 650866 364868 650898
rect 383868 651454 384868 651486
rect 383868 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 384868 651454
rect 383868 651134 384868 651218
rect 383868 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 384868 651134
rect 383868 650866 384868 650898
rect 403868 651454 404868 651486
rect 403868 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 404868 651454
rect 403868 651134 404868 651218
rect 403868 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 404868 651134
rect 403868 650866 404868 650898
rect 423868 651454 424868 651486
rect 423868 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 424868 651454
rect 423868 651134 424868 651218
rect 423868 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 424868 651134
rect 423868 650866 424868 650898
rect 443868 651454 444868 651486
rect 443868 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 444868 651454
rect 443868 651134 444868 651218
rect 443868 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 444868 651134
rect 443868 650866 444868 650898
rect 463868 651454 464868 651486
rect 463868 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 464868 651454
rect 463868 651134 464868 651218
rect 463868 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 464868 651134
rect 463868 650866 464868 650898
rect 483868 651454 484868 651486
rect 483868 651218 483930 651454
rect 484166 651218 484250 651454
rect 484486 651218 484570 651454
rect 484806 651218 484868 651454
rect 483868 651134 484868 651218
rect 483868 650898 483930 651134
rect 484166 650898 484250 651134
rect 484486 650898 484570 651134
rect 484806 650898 484868 651134
rect 483868 650866 484868 650898
rect 503868 651454 504868 651486
rect 503868 651218 503930 651454
rect 504166 651218 504250 651454
rect 504486 651218 504570 651454
rect 504806 651218 504868 651454
rect 503868 651134 504868 651218
rect 503868 650898 503930 651134
rect 504166 650898 504250 651134
rect 504486 650898 504570 651134
rect 504806 650898 504868 651134
rect 503868 650866 504868 650898
rect 523868 651454 524868 651486
rect 523868 651218 523930 651454
rect 524166 651218 524250 651454
rect 524486 651218 524570 651454
rect 524806 651218 524868 651454
rect 523868 651134 524868 651218
rect 523868 650898 523930 651134
rect 524166 650898 524250 651134
rect 524486 650898 524570 651134
rect 524806 650898 524868 651134
rect 523868 650866 524868 650898
rect 543868 651454 544868 651486
rect 543868 651218 543930 651454
rect 544166 651218 544250 651454
rect 544486 651218 544570 651454
rect 544806 651218 544868 651454
rect 543868 651134 544868 651218
rect 543868 650898 543930 651134
rect 544166 650898 544250 651134
rect 544486 650898 544570 651134
rect 544806 650898 544868 651134
rect 543868 650866 544868 650898
rect 563868 651454 564868 651486
rect 563868 651218 563930 651454
rect 564166 651218 564250 651454
rect 564486 651218 564570 651454
rect 564806 651218 564868 651454
rect 563868 651134 564868 651218
rect 563868 650898 563930 651134
rect 564166 650898 564250 651134
rect 564486 650898 564570 651134
rect 564806 650898 564868 651134
rect 563868 650866 564868 650898
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 313868 619954 314868 619986
rect 313868 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 314868 619954
rect 313868 619634 314868 619718
rect 313868 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 314868 619634
rect 313868 619366 314868 619398
rect 333868 619954 334868 619986
rect 333868 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 334868 619954
rect 333868 619634 334868 619718
rect 333868 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 334868 619634
rect 333868 619366 334868 619398
rect 353868 619954 354868 619986
rect 353868 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 354868 619954
rect 353868 619634 354868 619718
rect 353868 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 354868 619634
rect 353868 619366 354868 619398
rect 373868 619954 374868 619986
rect 373868 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 374868 619954
rect 373868 619634 374868 619718
rect 373868 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 374868 619634
rect 373868 619366 374868 619398
rect 393868 619954 394868 619986
rect 393868 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 394868 619954
rect 393868 619634 394868 619718
rect 393868 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 394868 619634
rect 393868 619366 394868 619398
rect 413868 619954 414868 619986
rect 413868 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 414868 619954
rect 413868 619634 414868 619718
rect 413868 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 414868 619634
rect 413868 619366 414868 619398
rect 433868 619954 434868 619986
rect 433868 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 434868 619954
rect 433868 619634 434868 619718
rect 433868 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 434868 619634
rect 433868 619366 434868 619398
rect 453868 619954 454868 619986
rect 453868 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 454868 619954
rect 453868 619634 454868 619718
rect 453868 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 454868 619634
rect 453868 619366 454868 619398
rect 473868 619954 474868 619986
rect 473868 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 474868 619954
rect 473868 619634 474868 619718
rect 473868 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 474868 619634
rect 473868 619366 474868 619398
rect 493868 619954 494868 619986
rect 493868 619718 493930 619954
rect 494166 619718 494250 619954
rect 494486 619718 494570 619954
rect 494806 619718 494868 619954
rect 493868 619634 494868 619718
rect 493868 619398 493930 619634
rect 494166 619398 494250 619634
rect 494486 619398 494570 619634
rect 494806 619398 494868 619634
rect 493868 619366 494868 619398
rect 513868 619954 514868 619986
rect 513868 619718 513930 619954
rect 514166 619718 514250 619954
rect 514486 619718 514570 619954
rect 514806 619718 514868 619954
rect 513868 619634 514868 619718
rect 513868 619398 513930 619634
rect 514166 619398 514250 619634
rect 514486 619398 514570 619634
rect 514806 619398 514868 619634
rect 513868 619366 514868 619398
rect 533868 619954 534868 619986
rect 533868 619718 533930 619954
rect 534166 619718 534250 619954
rect 534486 619718 534570 619954
rect 534806 619718 534868 619954
rect 533868 619634 534868 619718
rect 533868 619398 533930 619634
rect 534166 619398 534250 619634
rect 534486 619398 534570 619634
rect 534806 619398 534868 619634
rect 533868 619366 534868 619398
rect 553868 619954 554868 619986
rect 553868 619718 553930 619954
rect 554166 619718 554250 619954
rect 554486 619718 554570 619954
rect 554806 619718 554868 619954
rect 553868 619634 554868 619718
rect 553868 619398 553930 619634
rect 554166 619398 554250 619634
rect 554486 619398 554570 619634
rect 554806 619398 554868 619634
rect 553868 619366 554868 619398
rect 303868 615454 304868 615486
rect 303868 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 304868 615454
rect 303868 615134 304868 615218
rect 303868 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 304868 615134
rect 303868 614866 304868 614898
rect 323868 615454 324868 615486
rect 323868 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 324868 615454
rect 323868 615134 324868 615218
rect 323868 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 324868 615134
rect 323868 614866 324868 614898
rect 343868 615454 344868 615486
rect 343868 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 344868 615454
rect 343868 615134 344868 615218
rect 343868 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 344868 615134
rect 343868 614866 344868 614898
rect 363868 615454 364868 615486
rect 363868 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 364868 615454
rect 363868 615134 364868 615218
rect 363868 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 364868 615134
rect 363868 614866 364868 614898
rect 383868 615454 384868 615486
rect 383868 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 384868 615454
rect 383868 615134 384868 615218
rect 383868 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 384868 615134
rect 383868 614866 384868 614898
rect 403868 615454 404868 615486
rect 403868 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 404868 615454
rect 403868 615134 404868 615218
rect 403868 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 404868 615134
rect 403868 614866 404868 614898
rect 423868 615454 424868 615486
rect 423868 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 424868 615454
rect 423868 615134 424868 615218
rect 423868 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 424868 615134
rect 423868 614866 424868 614898
rect 443868 615454 444868 615486
rect 443868 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 444868 615454
rect 443868 615134 444868 615218
rect 443868 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 444868 615134
rect 443868 614866 444868 614898
rect 463868 615454 464868 615486
rect 463868 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 464868 615454
rect 463868 615134 464868 615218
rect 463868 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 464868 615134
rect 463868 614866 464868 614898
rect 483868 615454 484868 615486
rect 483868 615218 483930 615454
rect 484166 615218 484250 615454
rect 484486 615218 484570 615454
rect 484806 615218 484868 615454
rect 483868 615134 484868 615218
rect 483868 614898 483930 615134
rect 484166 614898 484250 615134
rect 484486 614898 484570 615134
rect 484806 614898 484868 615134
rect 483868 614866 484868 614898
rect 503868 615454 504868 615486
rect 503868 615218 503930 615454
rect 504166 615218 504250 615454
rect 504486 615218 504570 615454
rect 504806 615218 504868 615454
rect 503868 615134 504868 615218
rect 503868 614898 503930 615134
rect 504166 614898 504250 615134
rect 504486 614898 504570 615134
rect 504806 614898 504868 615134
rect 503868 614866 504868 614898
rect 523868 615454 524868 615486
rect 523868 615218 523930 615454
rect 524166 615218 524250 615454
rect 524486 615218 524570 615454
rect 524806 615218 524868 615454
rect 523868 615134 524868 615218
rect 523868 614898 523930 615134
rect 524166 614898 524250 615134
rect 524486 614898 524570 615134
rect 524806 614898 524868 615134
rect 523868 614866 524868 614898
rect 543868 615454 544868 615486
rect 543868 615218 543930 615454
rect 544166 615218 544250 615454
rect 544486 615218 544570 615454
rect 544806 615218 544868 615454
rect 543868 615134 544868 615218
rect 543868 614898 543930 615134
rect 544166 614898 544250 615134
rect 544486 614898 544570 615134
rect 544806 614898 544868 615134
rect 543868 614866 544868 614898
rect 563868 615454 564868 615486
rect 563868 615218 563930 615454
rect 564166 615218 564250 615454
rect 564486 615218 564570 615454
rect 564806 615218 564868 615454
rect 563868 615134 564868 615218
rect 563868 614898 563930 615134
rect 564166 614898 564250 615134
rect 564486 614898 564570 615134
rect 564806 614898 564868 615134
rect 563868 614866 564868 614898
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 569539 591020 569605 591021
rect 569539 590956 569540 591020
rect 569604 590956 569605 591020
rect 569539 590955 569605 590956
rect 303475 585988 303541 585989
rect 303475 585924 303476 585988
rect 303540 585924 303541 585988
rect 303475 585923 303541 585924
rect 299979 585852 300045 585853
rect 299979 585788 299980 585852
rect 300044 585788 300045 585852
rect 299979 585787 300045 585788
rect 298691 582996 298757 582997
rect 298691 582932 298692 582996
rect 298756 582932 298757 582996
rect 298691 582931 298757 582932
rect 297219 571980 297285 571981
rect 297219 571916 297220 571980
rect 297284 571916 297285 571980
rect 297219 571915 297285 571916
rect 297222 57221 297282 571915
rect 298694 459237 298754 582931
rect 298691 459236 298757 459237
rect 298691 459172 298692 459236
rect 298756 459172 298757 459236
rect 298691 459171 298757 459172
rect 298694 458285 298754 459171
rect 298691 458284 298757 458285
rect 298691 458220 298692 458284
rect 298756 458220 298757 458284
rect 298691 458219 298757 458220
rect 298691 317524 298757 317525
rect 298691 317460 298692 317524
rect 298756 317460 298757 317524
rect 298691 317459 298757 317460
rect 298694 189005 298754 317459
rect 298691 189004 298757 189005
rect 298691 188940 298692 189004
rect 298756 188940 298757 189004
rect 298691 188939 298757 188940
rect 298875 188868 298941 188869
rect 298875 188804 298876 188868
rect 298940 188804 298941 188868
rect 298875 188803 298941 188804
rect 298878 66877 298938 188803
rect 299243 185604 299309 185605
rect 299243 185540 299244 185604
rect 299308 185540 299309 185604
rect 299243 185539 299309 185540
rect 299246 79933 299306 185539
rect 299243 79932 299309 79933
rect 299243 79868 299244 79932
rect 299308 79868 299309 79932
rect 299243 79867 299309 79868
rect 299982 76533 300042 585787
rect 302003 583132 302069 583133
rect 302003 583068 302004 583132
rect 302068 583068 302069 583132
rect 302003 583067 302069 583068
rect 302006 461277 302066 583067
rect 302003 461276 302069 461277
rect 302003 461212 302004 461276
rect 302068 461212 302069 461276
rect 302003 461211 302069 461212
rect 300899 332620 300965 332621
rect 300899 332556 300900 332620
rect 300964 332556 300965 332620
rect 300899 332555 300965 332556
rect 300902 204781 300962 332555
rect 302006 315757 302066 461211
rect 303478 461005 303538 585923
rect 565859 585716 565925 585717
rect 565859 585652 565860 585716
rect 565924 585652 565925 585716
rect 565859 585651 565925 585652
rect 313868 547954 314868 547986
rect 313868 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 314868 547954
rect 313868 547634 314868 547718
rect 313868 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 314868 547634
rect 313868 547366 314868 547398
rect 333868 547954 334868 547986
rect 333868 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 334868 547954
rect 333868 547634 334868 547718
rect 333868 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 334868 547634
rect 333868 547366 334868 547398
rect 353868 547954 354868 547986
rect 353868 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 354868 547954
rect 353868 547634 354868 547718
rect 353868 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 354868 547634
rect 353868 547366 354868 547398
rect 373868 547954 374868 547986
rect 373868 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 374868 547954
rect 373868 547634 374868 547718
rect 373868 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 374868 547634
rect 373868 547366 374868 547398
rect 393868 547954 394868 547986
rect 393868 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 394868 547954
rect 393868 547634 394868 547718
rect 393868 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 394868 547634
rect 393868 547366 394868 547398
rect 413868 547954 414868 547986
rect 413868 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 414868 547954
rect 413868 547634 414868 547718
rect 413868 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 414868 547634
rect 413868 547366 414868 547398
rect 433868 547954 434868 547986
rect 433868 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 434868 547954
rect 433868 547634 434868 547718
rect 433868 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 434868 547634
rect 433868 547366 434868 547398
rect 453868 547954 454868 547986
rect 453868 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 454868 547954
rect 453868 547634 454868 547718
rect 453868 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 454868 547634
rect 453868 547366 454868 547398
rect 473868 547954 474868 547986
rect 473868 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 474868 547954
rect 473868 547634 474868 547718
rect 473868 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 474868 547634
rect 473868 547366 474868 547398
rect 493868 547954 494868 547986
rect 493868 547718 493930 547954
rect 494166 547718 494250 547954
rect 494486 547718 494570 547954
rect 494806 547718 494868 547954
rect 493868 547634 494868 547718
rect 493868 547398 493930 547634
rect 494166 547398 494250 547634
rect 494486 547398 494570 547634
rect 494806 547398 494868 547634
rect 493868 547366 494868 547398
rect 513868 547954 514868 547986
rect 513868 547718 513930 547954
rect 514166 547718 514250 547954
rect 514486 547718 514570 547954
rect 514806 547718 514868 547954
rect 513868 547634 514868 547718
rect 513868 547398 513930 547634
rect 514166 547398 514250 547634
rect 514486 547398 514570 547634
rect 514806 547398 514868 547634
rect 513868 547366 514868 547398
rect 533868 547954 534868 547986
rect 533868 547718 533930 547954
rect 534166 547718 534250 547954
rect 534486 547718 534570 547954
rect 534806 547718 534868 547954
rect 533868 547634 534868 547718
rect 533868 547398 533930 547634
rect 534166 547398 534250 547634
rect 534486 547398 534570 547634
rect 534806 547398 534868 547634
rect 533868 547366 534868 547398
rect 553868 547954 554868 547986
rect 553868 547718 553930 547954
rect 554166 547718 554250 547954
rect 554486 547718 554570 547954
rect 554806 547718 554868 547954
rect 553868 547634 554868 547718
rect 553868 547398 553930 547634
rect 554166 547398 554250 547634
rect 554486 547398 554570 547634
rect 554806 547398 554868 547634
rect 553868 547366 554868 547398
rect 303868 543454 304868 543486
rect 303868 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 304868 543454
rect 303868 543134 304868 543218
rect 303868 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 304868 543134
rect 303868 542866 304868 542898
rect 323868 543454 324868 543486
rect 323868 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 324868 543454
rect 323868 543134 324868 543218
rect 323868 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 324868 543134
rect 323868 542866 324868 542898
rect 343868 543454 344868 543486
rect 343868 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 344868 543454
rect 343868 543134 344868 543218
rect 343868 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 344868 543134
rect 343868 542866 344868 542898
rect 363868 543454 364868 543486
rect 363868 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 364868 543454
rect 363868 543134 364868 543218
rect 363868 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 364868 543134
rect 363868 542866 364868 542898
rect 383868 543454 384868 543486
rect 383868 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 384868 543454
rect 383868 543134 384868 543218
rect 383868 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 384868 543134
rect 383868 542866 384868 542898
rect 403868 543454 404868 543486
rect 403868 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 404868 543454
rect 403868 543134 404868 543218
rect 403868 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 404868 543134
rect 403868 542866 404868 542898
rect 423868 543454 424868 543486
rect 423868 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 424868 543454
rect 423868 543134 424868 543218
rect 423868 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 424868 543134
rect 423868 542866 424868 542898
rect 443868 543454 444868 543486
rect 443868 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 444868 543454
rect 443868 543134 444868 543218
rect 443868 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 444868 543134
rect 443868 542866 444868 542898
rect 463868 543454 464868 543486
rect 463868 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 464868 543454
rect 463868 543134 464868 543218
rect 463868 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 464868 543134
rect 463868 542866 464868 542898
rect 483868 543454 484868 543486
rect 483868 543218 483930 543454
rect 484166 543218 484250 543454
rect 484486 543218 484570 543454
rect 484806 543218 484868 543454
rect 483868 543134 484868 543218
rect 483868 542898 483930 543134
rect 484166 542898 484250 543134
rect 484486 542898 484570 543134
rect 484806 542898 484868 543134
rect 483868 542866 484868 542898
rect 503868 543454 504868 543486
rect 503868 543218 503930 543454
rect 504166 543218 504250 543454
rect 504486 543218 504570 543454
rect 504806 543218 504868 543454
rect 503868 543134 504868 543218
rect 503868 542898 503930 543134
rect 504166 542898 504250 543134
rect 504486 542898 504570 543134
rect 504806 542898 504868 543134
rect 503868 542866 504868 542898
rect 523868 543454 524868 543486
rect 523868 543218 523930 543454
rect 524166 543218 524250 543454
rect 524486 543218 524570 543454
rect 524806 543218 524868 543454
rect 523868 543134 524868 543218
rect 523868 542898 523930 543134
rect 524166 542898 524250 543134
rect 524486 542898 524570 543134
rect 524806 542898 524868 543134
rect 523868 542866 524868 542898
rect 543868 543454 544868 543486
rect 543868 543218 543930 543454
rect 544166 543218 544250 543454
rect 544486 543218 544570 543454
rect 544806 543218 544868 543454
rect 543868 543134 544868 543218
rect 543868 542898 543930 543134
rect 544166 542898 544250 543134
rect 544486 542898 544570 543134
rect 544806 542898 544868 543134
rect 543868 542866 544868 542898
rect 563868 543454 564868 543486
rect 563868 543218 563930 543454
rect 564166 543218 564250 543454
rect 564486 543218 564570 543454
rect 564806 543218 564868 543454
rect 563868 543134 564868 543218
rect 563868 542898 563930 543134
rect 564166 542898 564250 543134
rect 564486 542898 564570 543134
rect 564806 542898 564868 543134
rect 563868 542866 564868 542898
rect 313868 511954 314868 511986
rect 313868 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 314868 511954
rect 313868 511634 314868 511718
rect 313868 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 314868 511634
rect 313868 511366 314868 511398
rect 333868 511954 334868 511986
rect 333868 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 334868 511954
rect 333868 511634 334868 511718
rect 333868 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 334868 511634
rect 333868 511366 334868 511398
rect 353868 511954 354868 511986
rect 353868 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 354868 511954
rect 353868 511634 354868 511718
rect 353868 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 354868 511634
rect 353868 511366 354868 511398
rect 373868 511954 374868 511986
rect 373868 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 374868 511954
rect 373868 511634 374868 511718
rect 373868 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 374868 511634
rect 373868 511366 374868 511398
rect 393868 511954 394868 511986
rect 393868 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 394868 511954
rect 393868 511634 394868 511718
rect 393868 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 394868 511634
rect 393868 511366 394868 511398
rect 413868 511954 414868 511986
rect 413868 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 414868 511954
rect 413868 511634 414868 511718
rect 413868 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 414868 511634
rect 413868 511366 414868 511398
rect 433868 511954 434868 511986
rect 433868 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 434868 511954
rect 433868 511634 434868 511718
rect 433868 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 434868 511634
rect 433868 511366 434868 511398
rect 453868 511954 454868 511986
rect 453868 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 454868 511954
rect 453868 511634 454868 511718
rect 453868 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 454868 511634
rect 453868 511366 454868 511398
rect 473868 511954 474868 511986
rect 473868 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 474868 511954
rect 473868 511634 474868 511718
rect 473868 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 474868 511634
rect 473868 511366 474868 511398
rect 493868 511954 494868 511986
rect 493868 511718 493930 511954
rect 494166 511718 494250 511954
rect 494486 511718 494570 511954
rect 494806 511718 494868 511954
rect 493868 511634 494868 511718
rect 493868 511398 493930 511634
rect 494166 511398 494250 511634
rect 494486 511398 494570 511634
rect 494806 511398 494868 511634
rect 493868 511366 494868 511398
rect 513868 511954 514868 511986
rect 513868 511718 513930 511954
rect 514166 511718 514250 511954
rect 514486 511718 514570 511954
rect 514806 511718 514868 511954
rect 513868 511634 514868 511718
rect 513868 511398 513930 511634
rect 514166 511398 514250 511634
rect 514486 511398 514570 511634
rect 514806 511398 514868 511634
rect 513868 511366 514868 511398
rect 533868 511954 534868 511986
rect 533868 511718 533930 511954
rect 534166 511718 534250 511954
rect 534486 511718 534570 511954
rect 534806 511718 534868 511954
rect 533868 511634 534868 511718
rect 533868 511398 533930 511634
rect 534166 511398 534250 511634
rect 534486 511398 534570 511634
rect 534806 511398 534868 511634
rect 533868 511366 534868 511398
rect 553868 511954 554868 511986
rect 553868 511718 553930 511954
rect 554166 511718 554250 511954
rect 554486 511718 554570 511954
rect 554806 511718 554868 511954
rect 553868 511634 554868 511718
rect 553868 511398 553930 511634
rect 554166 511398 554250 511634
rect 554486 511398 554570 511634
rect 554806 511398 554868 511634
rect 553868 511366 554868 511398
rect 303868 507454 304868 507486
rect 303868 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 304868 507454
rect 303868 507134 304868 507218
rect 303868 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 304868 507134
rect 303868 506866 304868 506898
rect 323868 507454 324868 507486
rect 323868 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 324868 507454
rect 323868 507134 324868 507218
rect 323868 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 324868 507134
rect 323868 506866 324868 506898
rect 343868 507454 344868 507486
rect 343868 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 344868 507454
rect 343868 507134 344868 507218
rect 343868 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 344868 507134
rect 343868 506866 344868 506898
rect 363868 507454 364868 507486
rect 363868 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 364868 507454
rect 363868 507134 364868 507218
rect 363868 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 364868 507134
rect 363868 506866 364868 506898
rect 383868 507454 384868 507486
rect 383868 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 384868 507454
rect 383868 507134 384868 507218
rect 383868 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 384868 507134
rect 383868 506866 384868 506898
rect 403868 507454 404868 507486
rect 403868 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 404868 507454
rect 403868 507134 404868 507218
rect 403868 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 404868 507134
rect 403868 506866 404868 506898
rect 423868 507454 424868 507486
rect 423868 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 424868 507454
rect 423868 507134 424868 507218
rect 423868 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 424868 507134
rect 423868 506866 424868 506898
rect 443868 507454 444868 507486
rect 443868 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 444868 507454
rect 443868 507134 444868 507218
rect 443868 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 444868 507134
rect 443868 506866 444868 506898
rect 463868 507454 464868 507486
rect 463868 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 464868 507454
rect 463868 507134 464868 507218
rect 463868 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 464868 507134
rect 463868 506866 464868 506898
rect 483868 507454 484868 507486
rect 483868 507218 483930 507454
rect 484166 507218 484250 507454
rect 484486 507218 484570 507454
rect 484806 507218 484868 507454
rect 483868 507134 484868 507218
rect 483868 506898 483930 507134
rect 484166 506898 484250 507134
rect 484486 506898 484570 507134
rect 484806 506898 484868 507134
rect 483868 506866 484868 506898
rect 503868 507454 504868 507486
rect 503868 507218 503930 507454
rect 504166 507218 504250 507454
rect 504486 507218 504570 507454
rect 504806 507218 504868 507454
rect 503868 507134 504868 507218
rect 503868 506898 503930 507134
rect 504166 506898 504250 507134
rect 504486 506898 504570 507134
rect 504806 506898 504868 507134
rect 503868 506866 504868 506898
rect 523868 507454 524868 507486
rect 523868 507218 523930 507454
rect 524166 507218 524250 507454
rect 524486 507218 524570 507454
rect 524806 507218 524868 507454
rect 523868 507134 524868 507218
rect 523868 506898 523930 507134
rect 524166 506898 524250 507134
rect 524486 506898 524570 507134
rect 524806 506898 524868 507134
rect 523868 506866 524868 506898
rect 543868 507454 544868 507486
rect 543868 507218 543930 507454
rect 544166 507218 544250 507454
rect 544486 507218 544570 507454
rect 544806 507218 544868 507454
rect 543868 507134 544868 507218
rect 543868 506898 543930 507134
rect 544166 506898 544250 507134
rect 544486 506898 544570 507134
rect 544806 506898 544868 507134
rect 543868 506866 544868 506898
rect 563868 507454 564868 507486
rect 563868 507218 563930 507454
rect 564166 507218 564250 507454
rect 564486 507218 564570 507454
rect 564806 507218 564868 507454
rect 563868 507134 564868 507218
rect 563868 506898 563930 507134
rect 564166 506898 564250 507134
rect 564486 506898 564570 507134
rect 564806 506898 564868 507134
rect 563868 506866 564868 506898
rect 565862 480270 565922 585651
rect 568619 580276 568685 580277
rect 568619 580212 568620 580276
rect 568684 580212 568685 580276
rect 568619 580211 568685 580212
rect 567883 571980 567949 571981
rect 567883 571916 567884 571980
rect 567948 571916 567949 571980
rect 567883 571915 567949 571916
rect 565862 480210 566474 480270
rect 313868 475954 314868 475986
rect 313868 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 314868 475954
rect 313868 475634 314868 475718
rect 313868 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 314868 475634
rect 313868 475366 314868 475398
rect 333868 475954 334868 475986
rect 333868 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 334868 475954
rect 333868 475634 334868 475718
rect 333868 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 334868 475634
rect 333868 475366 334868 475398
rect 353868 475954 354868 475986
rect 353868 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 354868 475954
rect 353868 475634 354868 475718
rect 353868 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 354868 475634
rect 353868 475366 354868 475398
rect 373868 475954 374868 475986
rect 373868 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 374868 475954
rect 373868 475634 374868 475718
rect 373868 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 374868 475634
rect 373868 475366 374868 475398
rect 393868 475954 394868 475986
rect 393868 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 394868 475954
rect 393868 475634 394868 475718
rect 393868 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 394868 475634
rect 393868 475366 394868 475398
rect 413868 475954 414868 475986
rect 413868 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 414868 475954
rect 413868 475634 414868 475718
rect 413868 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 414868 475634
rect 413868 475366 414868 475398
rect 433868 475954 434868 475986
rect 433868 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 434868 475954
rect 433868 475634 434868 475718
rect 433868 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 434868 475634
rect 433868 475366 434868 475398
rect 453868 475954 454868 475986
rect 453868 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 454868 475954
rect 453868 475634 454868 475718
rect 453868 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 454868 475634
rect 453868 475366 454868 475398
rect 473868 475954 474868 475986
rect 473868 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 474868 475954
rect 473868 475634 474868 475718
rect 473868 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 474868 475634
rect 473868 475366 474868 475398
rect 493868 475954 494868 475986
rect 493868 475718 493930 475954
rect 494166 475718 494250 475954
rect 494486 475718 494570 475954
rect 494806 475718 494868 475954
rect 493868 475634 494868 475718
rect 493868 475398 493930 475634
rect 494166 475398 494250 475634
rect 494486 475398 494570 475634
rect 494806 475398 494868 475634
rect 493868 475366 494868 475398
rect 513868 475954 514868 475986
rect 513868 475718 513930 475954
rect 514166 475718 514250 475954
rect 514486 475718 514570 475954
rect 514806 475718 514868 475954
rect 513868 475634 514868 475718
rect 513868 475398 513930 475634
rect 514166 475398 514250 475634
rect 514486 475398 514570 475634
rect 514806 475398 514868 475634
rect 513868 475366 514868 475398
rect 533868 475954 534868 475986
rect 533868 475718 533930 475954
rect 534166 475718 534250 475954
rect 534486 475718 534570 475954
rect 534806 475718 534868 475954
rect 533868 475634 534868 475718
rect 533868 475398 533930 475634
rect 534166 475398 534250 475634
rect 534486 475398 534570 475634
rect 534806 475398 534868 475634
rect 533868 475366 534868 475398
rect 553868 475954 554868 475986
rect 553868 475718 553930 475954
rect 554166 475718 554250 475954
rect 554486 475718 554570 475954
rect 554806 475718 554868 475954
rect 553868 475634 554868 475718
rect 553868 475398 553930 475634
rect 554166 475398 554250 475634
rect 554486 475398 554570 475634
rect 554806 475398 554868 475634
rect 553868 475366 554868 475398
rect 303868 471454 304868 471486
rect 303868 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 304868 471454
rect 303868 471134 304868 471218
rect 303868 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 304868 471134
rect 303868 470866 304868 470898
rect 323868 471454 324868 471486
rect 323868 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 324868 471454
rect 323868 471134 324868 471218
rect 323868 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 324868 471134
rect 323868 470866 324868 470898
rect 343868 471454 344868 471486
rect 343868 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 344868 471454
rect 343868 471134 344868 471218
rect 343868 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 344868 471134
rect 343868 470866 344868 470898
rect 363868 471454 364868 471486
rect 363868 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 364868 471454
rect 363868 471134 364868 471218
rect 363868 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 364868 471134
rect 363868 470866 364868 470898
rect 383868 471454 384868 471486
rect 383868 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 384868 471454
rect 383868 471134 384868 471218
rect 383868 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 384868 471134
rect 383868 470866 384868 470898
rect 403868 471454 404868 471486
rect 403868 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 404868 471454
rect 403868 471134 404868 471218
rect 403868 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 404868 471134
rect 403868 470866 404868 470898
rect 423868 471454 424868 471486
rect 423868 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 424868 471454
rect 423868 471134 424868 471218
rect 423868 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 424868 471134
rect 423868 470866 424868 470898
rect 443868 471454 444868 471486
rect 443868 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 444868 471454
rect 443868 471134 444868 471218
rect 443868 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 444868 471134
rect 443868 470866 444868 470898
rect 463868 471454 464868 471486
rect 463868 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 464868 471454
rect 463868 471134 464868 471218
rect 463868 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 464868 471134
rect 463868 470866 464868 470898
rect 483868 471454 484868 471486
rect 483868 471218 483930 471454
rect 484166 471218 484250 471454
rect 484486 471218 484570 471454
rect 484806 471218 484868 471454
rect 483868 471134 484868 471218
rect 483868 470898 483930 471134
rect 484166 470898 484250 471134
rect 484486 470898 484570 471134
rect 484806 470898 484868 471134
rect 483868 470866 484868 470898
rect 503868 471454 504868 471486
rect 503868 471218 503930 471454
rect 504166 471218 504250 471454
rect 504486 471218 504570 471454
rect 504806 471218 504868 471454
rect 503868 471134 504868 471218
rect 503868 470898 503930 471134
rect 504166 470898 504250 471134
rect 504486 470898 504570 471134
rect 504806 470898 504868 471134
rect 503868 470866 504868 470898
rect 523868 471454 524868 471486
rect 523868 471218 523930 471454
rect 524166 471218 524250 471454
rect 524486 471218 524570 471454
rect 524806 471218 524868 471454
rect 523868 471134 524868 471218
rect 523868 470898 523930 471134
rect 524166 470898 524250 471134
rect 524486 470898 524570 471134
rect 524806 470898 524868 471134
rect 523868 470866 524868 470898
rect 543868 471454 544868 471486
rect 543868 471218 543930 471454
rect 544166 471218 544250 471454
rect 544486 471218 544570 471454
rect 544806 471218 544868 471454
rect 543868 471134 544868 471218
rect 543868 470898 543930 471134
rect 544166 470898 544250 471134
rect 544486 470898 544570 471134
rect 544806 470898 544868 471134
rect 543868 470866 544868 470898
rect 563868 471454 564868 471486
rect 563868 471218 563930 471454
rect 564166 471218 564250 471454
rect 564486 471218 564570 471454
rect 564806 471218 564868 471454
rect 563868 471134 564868 471218
rect 563868 470898 563930 471134
rect 564166 470898 564250 471134
rect 564486 470898 564570 471134
rect 564806 470898 564868 471134
rect 563868 470866 564868 470898
rect 303475 461004 303541 461005
rect 303475 460940 303476 461004
rect 303540 460940 303541 461004
rect 303475 460939 303541 460940
rect 303478 451290 303538 460939
rect 566414 458149 566474 480210
rect 567699 461140 567765 461141
rect 567699 461076 567700 461140
rect 567764 461076 567765 461140
rect 567699 461075 567765 461076
rect 566411 458148 566477 458149
rect 566411 458084 566412 458148
rect 566476 458084 566477 458148
rect 566411 458083 566477 458084
rect 302742 451230 303538 451290
rect 302742 332213 302802 451230
rect 313868 439954 314868 439986
rect 313868 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 314868 439954
rect 313868 439634 314868 439718
rect 313868 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 314868 439634
rect 313868 439366 314868 439398
rect 333868 439954 334868 439986
rect 333868 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 334868 439954
rect 333868 439634 334868 439718
rect 333868 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 334868 439634
rect 333868 439366 334868 439398
rect 353868 439954 354868 439986
rect 353868 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 354868 439954
rect 353868 439634 354868 439718
rect 353868 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 354868 439634
rect 353868 439366 354868 439398
rect 373868 439954 374868 439986
rect 373868 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 374868 439954
rect 373868 439634 374868 439718
rect 373868 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 374868 439634
rect 373868 439366 374868 439398
rect 393868 439954 394868 439986
rect 393868 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 394868 439954
rect 393868 439634 394868 439718
rect 393868 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 394868 439634
rect 393868 439366 394868 439398
rect 413868 439954 414868 439986
rect 413868 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 414868 439954
rect 413868 439634 414868 439718
rect 413868 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 414868 439634
rect 413868 439366 414868 439398
rect 433868 439954 434868 439986
rect 433868 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 434868 439954
rect 433868 439634 434868 439718
rect 433868 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 434868 439634
rect 433868 439366 434868 439398
rect 453868 439954 454868 439986
rect 453868 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 454868 439954
rect 453868 439634 454868 439718
rect 453868 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 454868 439634
rect 453868 439366 454868 439398
rect 473868 439954 474868 439986
rect 473868 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 474868 439954
rect 473868 439634 474868 439718
rect 473868 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 474868 439634
rect 473868 439366 474868 439398
rect 493868 439954 494868 439986
rect 493868 439718 493930 439954
rect 494166 439718 494250 439954
rect 494486 439718 494570 439954
rect 494806 439718 494868 439954
rect 493868 439634 494868 439718
rect 493868 439398 493930 439634
rect 494166 439398 494250 439634
rect 494486 439398 494570 439634
rect 494806 439398 494868 439634
rect 493868 439366 494868 439398
rect 513868 439954 514868 439986
rect 513868 439718 513930 439954
rect 514166 439718 514250 439954
rect 514486 439718 514570 439954
rect 514806 439718 514868 439954
rect 513868 439634 514868 439718
rect 513868 439398 513930 439634
rect 514166 439398 514250 439634
rect 514486 439398 514570 439634
rect 514806 439398 514868 439634
rect 513868 439366 514868 439398
rect 533868 439954 534868 439986
rect 533868 439718 533930 439954
rect 534166 439718 534250 439954
rect 534486 439718 534570 439954
rect 534806 439718 534868 439954
rect 533868 439634 534868 439718
rect 533868 439398 533930 439634
rect 534166 439398 534250 439634
rect 534486 439398 534570 439634
rect 534806 439398 534868 439634
rect 533868 439366 534868 439398
rect 553868 439954 554868 439986
rect 553868 439718 553930 439954
rect 554166 439718 554250 439954
rect 554486 439718 554570 439954
rect 554806 439718 554868 439954
rect 553868 439634 554868 439718
rect 553868 439398 553930 439634
rect 554166 439398 554250 439634
rect 554486 439398 554570 439634
rect 554806 439398 554868 439634
rect 553868 439366 554868 439398
rect 303868 435454 304868 435486
rect 303868 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 304868 435454
rect 303868 435134 304868 435218
rect 303868 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 304868 435134
rect 303868 434866 304868 434898
rect 323868 435454 324868 435486
rect 323868 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 324868 435454
rect 323868 435134 324868 435218
rect 323868 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 324868 435134
rect 323868 434866 324868 434898
rect 343868 435454 344868 435486
rect 343868 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 344868 435454
rect 343868 435134 344868 435218
rect 343868 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 344868 435134
rect 343868 434866 344868 434898
rect 363868 435454 364868 435486
rect 363868 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 364868 435454
rect 363868 435134 364868 435218
rect 363868 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 364868 435134
rect 363868 434866 364868 434898
rect 383868 435454 384868 435486
rect 383868 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 384868 435454
rect 383868 435134 384868 435218
rect 383868 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 384868 435134
rect 383868 434866 384868 434898
rect 403868 435454 404868 435486
rect 403868 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 404868 435454
rect 403868 435134 404868 435218
rect 403868 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 404868 435134
rect 403868 434866 404868 434898
rect 423868 435454 424868 435486
rect 423868 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 424868 435454
rect 423868 435134 424868 435218
rect 423868 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 424868 435134
rect 423868 434866 424868 434898
rect 443868 435454 444868 435486
rect 443868 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 444868 435454
rect 443868 435134 444868 435218
rect 443868 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 444868 435134
rect 443868 434866 444868 434898
rect 463868 435454 464868 435486
rect 463868 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 464868 435454
rect 463868 435134 464868 435218
rect 463868 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 464868 435134
rect 463868 434866 464868 434898
rect 483868 435454 484868 435486
rect 483868 435218 483930 435454
rect 484166 435218 484250 435454
rect 484486 435218 484570 435454
rect 484806 435218 484868 435454
rect 483868 435134 484868 435218
rect 483868 434898 483930 435134
rect 484166 434898 484250 435134
rect 484486 434898 484570 435134
rect 484806 434898 484868 435134
rect 483868 434866 484868 434898
rect 503868 435454 504868 435486
rect 503868 435218 503930 435454
rect 504166 435218 504250 435454
rect 504486 435218 504570 435454
rect 504806 435218 504868 435454
rect 503868 435134 504868 435218
rect 503868 434898 503930 435134
rect 504166 434898 504250 435134
rect 504486 434898 504570 435134
rect 504806 434898 504868 435134
rect 503868 434866 504868 434898
rect 523868 435454 524868 435486
rect 523868 435218 523930 435454
rect 524166 435218 524250 435454
rect 524486 435218 524570 435454
rect 524806 435218 524868 435454
rect 523868 435134 524868 435218
rect 523868 434898 523930 435134
rect 524166 434898 524250 435134
rect 524486 434898 524570 435134
rect 524806 434898 524868 435134
rect 523868 434866 524868 434898
rect 543868 435454 544868 435486
rect 543868 435218 543930 435454
rect 544166 435218 544250 435454
rect 544486 435218 544570 435454
rect 544806 435218 544868 435454
rect 543868 435134 544868 435218
rect 543868 434898 543930 435134
rect 544166 434898 544250 435134
rect 544486 434898 544570 435134
rect 544806 434898 544868 435134
rect 543868 434866 544868 434898
rect 563868 435454 564868 435486
rect 563868 435218 563930 435454
rect 564166 435218 564250 435454
rect 564486 435218 564570 435454
rect 564806 435218 564868 435454
rect 563868 435134 564868 435218
rect 563868 434898 563930 435134
rect 564166 434898 564250 435134
rect 564486 434898 564570 435134
rect 564806 434898 564868 435134
rect 563868 434866 564868 434898
rect 313868 403954 314868 403986
rect 313868 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 314868 403954
rect 313868 403634 314868 403718
rect 313868 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 314868 403634
rect 313868 403366 314868 403398
rect 333868 403954 334868 403986
rect 333868 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 334868 403954
rect 333868 403634 334868 403718
rect 333868 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 334868 403634
rect 333868 403366 334868 403398
rect 353868 403954 354868 403986
rect 353868 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 354868 403954
rect 353868 403634 354868 403718
rect 353868 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 354868 403634
rect 353868 403366 354868 403398
rect 373868 403954 374868 403986
rect 373868 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 374868 403954
rect 373868 403634 374868 403718
rect 373868 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 374868 403634
rect 373868 403366 374868 403398
rect 393868 403954 394868 403986
rect 393868 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 394868 403954
rect 393868 403634 394868 403718
rect 393868 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 394868 403634
rect 393868 403366 394868 403398
rect 413868 403954 414868 403986
rect 413868 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 414868 403954
rect 413868 403634 414868 403718
rect 413868 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 414868 403634
rect 413868 403366 414868 403398
rect 433868 403954 434868 403986
rect 433868 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 434868 403954
rect 433868 403634 434868 403718
rect 433868 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 434868 403634
rect 433868 403366 434868 403398
rect 453868 403954 454868 403986
rect 453868 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 454868 403954
rect 453868 403634 454868 403718
rect 453868 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 454868 403634
rect 453868 403366 454868 403398
rect 473868 403954 474868 403986
rect 473868 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 474868 403954
rect 473868 403634 474868 403718
rect 473868 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 474868 403634
rect 473868 403366 474868 403398
rect 493868 403954 494868 403986
rect 493868 403718 493930 403954
rect 494166 403718 494250 403954
rect 494486 403718 494570 403954
rect 494806 403718 494868 403954
rect 493868 403634 494868 403718
rect 493868 403398 493930 403634
rect 494166 403398 494250 403634
rect 494486 403398 494570 403634
rect 494806 403398 494868 403634
rect 493868 403366 494868 403398
rect 513868 403954 514868 403986
rect 513868 403718 513930 403954
rect 514166 403718 514250 403954
rect 514486 403718 514570 403954
rect 514806 403718 514868 403954
rect 513868 403634 514868 403718
rect 513868 403398 513930 403634
rect 514166 403398 514250 403634
rect 514486 403398 514570 403634
rect 514806 403398 514868 403634
rect 513868 403366 514868 403398
rect 533868 403954 534868 403986
rect 533868 403718 533930 403954
rect 534166 403718 534250 403954
rect 534486 403718 534570 403954
rect 534806 403718 534868 403954
rect 533868 403634 534868 403718
rect 533868 403398 533930 403634
rect 534166 403398 534250 403634
rect 534486 403398 534570 403634
rect 534806 403398 534868 403634
rect 533868 403366 534868 403398
rect 553868 403954 554868 403986
rect 553868 403718 553930 403954
rect 554166 403718 554250 403954
rect 554486 403718 554570 403954
rect 554806 403718 554868 403954
rect 553868 403634 554868 403718
rect 553868 403398 553930 403634
rect 554166 403398 554250 403634
rect 554486 403398 554570 403634
rect 554806 403398 554868 403634
rect 553868 403366 554868 403398
rect 303868 399454 304868 399486
rect 303868 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 304868 399454
rect 303868 399134 304868 399218
rect 303868 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 304868 399134
rect 303868 398866 304868 398898
rect 323868 399454 324868 399486
rect 323868 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 324868 399454
rect 323868 399134 324868 399218
rect 323868 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 324868 399134
rect 323868 398866 324868 398898
rect 343868 399454 344868 399486
rect 343868 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 344868 399454
rect 343868 399134 344868 399218
rect 343868 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 344868 399134
rect 343868 398866 344868 398898
rect 363868 399454 364868 399486
rect 363868 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 364868 399454
rect 363868 399134 364868 399218
rect 363868 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 364868 399134
rect 363868 398866 364868 398898
rect 383868 399454 384868 399486
rect 383868 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 384868 399454
rect 383868 399134 384868 399218
rect 383868 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 384868 399134
rect 383868 398866 384868 398898
rect 403868 399454 404868 399486
rect 403868 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 404868 399454
rect 403868 399134 404868 399218
rect 403868 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 404868 399134
rect 403868 398866 404868 398898
rect 423868 399454 424868 399486
rect 423868 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 424868 399454
rect 423868 399134 424868 399218
rect 423868 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 424868 399134
rect 423868 398866 424868 398898
rect 443868 399454 444868 399486
rect 443868 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 444868 399454
rect 443868 399134 444868 399218
rect 443868 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 444868 399134
rect 443868 398866 444868 398898
rect 463868 399454 464868 399486
rect 463868 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 464868 399454
rect 463868 399134 464868 399218
rect 463868 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 464868 399134
rect 463868 398866 464868 398898
rect 483868 399454 484868 399486
rect 483868 399218 483930 399454
rect 484166 399218 484250 399454
rect 484486 399218 484570 399454
rect 484806 399218 484868 399454
rect 483868 399134 484868 399218
rect 483868 398898 483930 399134
rect 484166 398898 484250 399134
rect 484486 398898 484570 399134
rect 484806 398898 484868 399134
rect 483868 398866 484868 398898
rect 503868 399454 504868 399486
rect 503868 399218 503930 399454
rect 504166 399218 504250 399454
rect 504486 399218 504570 399454
rect 504806 399218 504868 399454
rect 503868 399134 504868 399218
rect 503868 398898 503930 399134
rect 504166 398898 504250 399134
rect 504486 398898 504570 399134
rect 504806 398898 504868 399134
rect 503868 398866 504868 398898
rect 523868 399454 524868 399486
rect 523868 399218 523930 399454
rect 524166 399218 524250 399454
rect 524486 399218 524570 399454
rect 524806 399218 524868 399454
rect 523868 399134 524868 399218
rect 523868 398898 523930 399134
rect 524166 398898 524250 399134
rect 524486 398898 524570 399134
rect 524806 398898 524868 399134
rect 523868 398866 524868 398898
rect 543868 399454 544868 399486
rect 543868 399218 543930 399454
rect 544166 399218 544250 399454
rect 544486 399218 544570 399454
rect 544806 399218 544868 399454
rect 543868 399134 544868 399218
rect 543868 398898 543930 399134
rect 544166 398898 544250 399134
rect 544486 398898 544570 399134
rect 544806 398898 544868 399134
rect 543868 398866 544868 398898
rect 563868 399454 564868 399486
rect 563868 399218 563930 399454
rect 564166 399218 564250 399454
rect 564486 399218 564570 399454
rect 564806 399218 564868 399454
rect 563868 399134 564868 399218
rect 563868 398898 563930 399134
rect 564166 398898 564250 399134
rect 564486 398898 564570 399134
rect 564806 398898 564868 399134
rect 563868 398866 564868 398898
rect 313868 367954 314868 367986
rect 313868 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 314868 367954
rect 313868 367634 314868 367718
rect 313868 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 314868 367634
rect 313868 367366 314868 367398
rect 333868 367954 334868 367986
rect 333868 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 334868 367954
rect 333868 367634 334868 367718
rect 333868 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 334868 367634
rect 333868 367366 334868 367398
rect 353868 367954 354868 367986
rect 353868 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 354868 367954
rect 353868 367634 354868 367718
rect 353868 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 354868 367634
rect 353868 367366 354868 367398
rect 373868 367954 374868 367986
rect 373868 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 374868 367954
rect 373868 367634 374868 367718
rect 373868 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 374868 367634
rect 373868 367366 374868 367398
rect 393868 367954 394868 367986
rect 393868 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 394868 367954
rect 393868 367634 394868 367718
rect 393868 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 394868 367634
rect 393868 367366 394868 367398
rect 413868 367954 414868 367986
rect 413868 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 414868 367954
rect 413868 367634 414868 367718
rect 413868 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 414868 367634
rect 413868 367366 414868 367398
rect 433868 367954 434868 367986
rect 433868 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 434868 367954
rect 433868 367634 434868 367718
rect 433868 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 434868 367634
rect 433868 367366 434868 367398
rect 453868 367954 454868 367986
rect 453868 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 454868 367954
rect 453868 367634 454868 367718
rect 453868 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 454868 367634
rect 453868 367366 454868 367398
rect 473868 367954 474868 367986
rect 473868 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 474868 367954
rect 473868 367634 474868 367718
rect 473868 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 474868 367634
rect 473868 367366 474868 367398
rect 493868 367954 494868 367986
rect 493868 367718 493930 367954
rect 494166 367718 494250 367954
rect 494486 367718 494570 367954
rect 494806 367718 494868 367954
rect 493868 367634 494868 367718
rect 493868 367398 493930 367634
rect 494166 367398 494250 367634
rect 494486 367398 494570 367634
rect 494806 367398 494868 367634
rect 493868 367366 494868 367398
rect 513868 367954 514868 367986
rect 513868 367718 513930 367954
rect 514166 367718 514250 367954
rect 514486 367718 514570 367954
rect 514806 367718 514868 367954
rect 513868 367634 514868 367718
rect 513868 367398 513930 367634
rect 514166 367398 514250 367634
rect 514486 367398 514570 367634
rect 514806 367398 514868 367634
rect 513868 367366 514868 367398
rect 533868 367954 534868 367986
rect 533868 367718 533930 367954
rect 534166 367718 534250 367954
rect 534486 367718 534570 367954
rect 534806 367718 534868 367954
rect 533868 367634 534868 367718
rect 533868 367398 533930 367634
rect 534166 367398 534250 367634
rect 534486 367398 534570 367634
rect 534806 367398 534868 367634
rect 533868 367366 534868 367398
rect 553868 367954 554868 367986
rect 553868 367718 553930 367954
rect 554166 367718 554250 367954
rect 554486 367718 554570 367954
rect 554806 367718 554868 367954
rect 553868 367634 554868 367718
rect 553868 367398 553930 367634
rect 554166 367398 554250 367634
rect 554486 367398 554570 367634
rect 554806 367398 554868 367634
rect 553868 367366 554868 367398
rect 303868 363454 304868 363486
rect 303868 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 304868 363454
rect 303868 363134 304868 363218
rect 303868 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 304868 363134
rect 303868 362866 304868 362898
rect 323868 363454 324868 363486
rect 323868 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 324868 363454
rect 323868 363134 324868 363218
rect 323868 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 324868 363134
rect 323868 362866 324868 362898
rect 343868 363454 344868 363486
rect 343868 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 344868 363454
rect 343868 363134 344868 363218
rect 343868 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 344868 363134
rect 343868 362866 344868 362898
rect 363868 363454 364868 363486
rect 363868 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 364868 363454
rect 363868 363134 364868 363218
rect 363868 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 364868 363134
rect 363868 362866 364868 362898
rect 383868 363454 384868 363486
rect 383868 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 384868 363454
rect 383868 363134 384868 363218
rect 383868 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 384868 363134
rect 383868 362866 384868 362898
rect 403868 363454 404868 363486
rect 403868 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 404868 363454
rect 403868 363134 404868 363218
rect 403868 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 404868 363134
rect 403868 362866 404868 362898
rect 423868 363454 424868 363486
rect 423868 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 424868 363454
rect 423868 363134 424868 363218
rect 423868 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 424868 363134
rect 423868 362866 424868 362898
rect 443868 363454 444868 363486
rect 443868 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 444868 363454
rect 443868 363134 444868 363218
rect 443868 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 444868 363134
rect 443868 362866 444868 362898
rect 463868 363454 464868 363486
rect 463868 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 464868 363454
rect 463868 363134 464868 363218
rect 463868 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 464868 363134
rect 463868 362866 464868 362898
rect 483868 363454 484868 363486
rect 483868 363218 483930 363454
rect 484166 363218 484250 363454
rect 484486 363218 484570 363454
rect 484806 363218 484868 363454
rect 483868 363134 484868 363218
rect 483868 362898 483930 363134
rect 484166 362898 484250 363134
rect 484486 362898 484570 363134
rect 484806 362898 484868 363134
rect 483868 362866 484868 362898
rect 503868 363454 504868 363486
rect 503868 363218 503930 363454
rect 504166 363218 504250 363454
rect 504486 363218 504570 363454
rect 504806 363218 504868 363454
rect 503868 363134 504868 363218
rect 503868 362898 503930 363134
rect 504166 362898 504250 363134
rect 504486 362898 504570 363134
rect 504806 362898 504868 363134
rect 503868 362866 504868 362898
rect 523868 363454 524868 363486
rect 523868 363218 523930 363454
rect 524166 363218 524250 363454
rect 524486 363218 524570 363454
rect 524806 363218 524868 363454
rect 523868 363134 524868 363218
rect 523868 362898 523930 363134
rect 524166 362898 524250 363134
rect 524486 362898 524570 363134
rect 524806 362898 524868 363134
rect 523868 362866 524868 362898
rect 543868 363454 544868 363486
rect 543868 363218 543930 363454
rect 544166 363218 544250 363454
rect 544486 363218 544570 363454
rect 544806 363218 544868 363454
rect 543868 363134 544868 363218
rect 543868 362898 543930 363134
rect 544166 362898 544250 363134
rect 544486 362898 544570 363134
rect 544806 362898 544868 363134
rect 543868 362866 544868 362898
rect 563868 363454 564868 363486
rect 563868 363218 563930 363454
rect 564166 363218 564250 363454
rect 564486 363218 564570 363454
rect 564806 363218 564868 363454
rect 563868 363134 564868 363218
rect 563868 362898 563930 363134
rect 564166 362898 564250 363134
rect 564486 362898 564570 363134
rect 564806 362898 564868 363134
rect 563868 362866 564868 362898
rect 566414 335370 566474 458083
rect 565862 335310 566474 335370
rect 565862 332349 565922 335310
rect 565859 332348 565925 332349
rect 565859 332284 565860 332348
rect 565924 332284 565925 332348
rect 565859 332283 565925 332284
rect 302739 332212 302805 332213
rect 302739 332148 302740 332212
rect 302804 332148 302805 332212
rect 302739 332147 302805 332148
rect 302003 315756 302069 315757
rect 302003 315692 302004 315756
rect 302068 315692 302069 315756
rect 302003 315691 302069 315692
rect 302006 314805 302066 315691
rect 302003 314804 302069 314805
rect 302003 314740 302004 314804
rect 302068 314740 302069 314804
rect 302003 314739 302069 314740
rect 300899 204780 300965 204781
rect 300899 204716 300900 204780
rect 300964 204716 300965 204780
rect 300899 204715 300965 204716
rect 302003 204780 302069 204781
rect 302003 204716 302004 204780
rect 302068 204716 302069 204780
rect 302003 204715 302069 204716
rect 301451 186420 301517 186421
rect 301451 186356 301452 186420
rect 301516 186356 301517 186420
rect 301451 186355 301517 186356
rect 301454 161490 301514 186355
rect 300902 161430 301514 161490
rect 300902 158810 300962 161430
rect 300718 158750 300962 158810
rect 300718 80205 300778 158750
rect 300715 80204 300781 80205
rect 300715 80140 300716 80204
rect 300780 80140 300781 80204
rect 300715 80139 300781 80140
rect 299979 76532 300045 76533
rect 299979 76468 299980 76532
rect 300044 76468 300045 76532
rect 299979 76467 300045 76468
rect 298875 66876 298941 66877
rect 298875 66812 298876 66876
rect 298940 66812 298941 66876
rect 298875 66811 298941 66812
rect 302006 58581 302066 204715
rect 302742 201381 302802 332147
rect 313868 295954 314868 295986
rect 313868 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 314868 295954
rect 313868 295634 314868 295718
rect 313868 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 314868 295634
rect 313868 295366 314868 295398
rect 333868 295954 334868 295986
rect 333868 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 334868 295954
rect 333868 295634 334868 295718
rect 333868 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 334868 295634
rect 333868 295366 334868 295398
rect 353868 295954 354868 295986
rect 353868 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 354868 295954
rect 353868 295634 354868 295718
rect 353868 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 354868 295634
rect 353868 295366 354868 295398
rect 373868 295954 374868 295986
rect 373868 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 374868 295954
rect 373868 295634 374868 295718
rect 373868 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 374868 295634
rect 373868 295366 374868 295398
rect 393868 295954 394868 295986
rect 393868 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 394868 295954
rect 393868 295634 394868 295718
rect 393868 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 394868 295634
rect 393868 295366 394868 295398
rect 413868 295954 414868 295986
rect 413868 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 414868 295954
rect 413868 295634 414868 295718
rect 413868 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 414868 295634
rect 413868 295366 414868 295398
rect 433868 295954 434868 295986
rect 433868 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 434868 295954
rect 433868 295634 434868 295718
rect 433868 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 434868 295634
rect 433868 295366 434868 295398
rect 453868 295954 454868 295986
rect 453868 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 454868 295954
rect 453868 295634 454868 295718
rect 453868 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 454868 295634
rect 453868 295366 454868 295398
rect 473868 295954 474868 295986
rect 473868 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 474868 295954
rect 473868 295634 474868 295718
rect 473868 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 474868 295634
rect 473868 295366 474868 295398
rect 493868 295954 494868 295986
rect 493868 295718 493930 295954
rect 494166 295718 494250 295954
rect 494486 295718 494570 295954
rect 494806 295718 494868 295954
rect 493868 295634 494868 295718
rect 493868 295398 493930 295634
rect 494166 295398 494250 295634
rect 494486 295398 494570 295634
rect 494806 295398 494868 295634
rect 493868 295366 494868 295398
rect 513868 295954 514868 295986
rect 513868 295718 513930 295954
rect 514166 295718 514250 295954
rect 514486 295718 514570 295954
rect 514806 295718 514868 295954
rect 513868 295634 514868 295718
rect 513868 295398 513930 295634
rect 514166 295398 514250 295634
rect 514486 295398 514570 295634
rect 514806 295398 514868 295634
rect 513868 295366 514868 295398
rect 533868 295954 534868 295986
rect 533868 295718 533930 295954
rect 534166 295718 534250 295954
rect 534486 295718 534570 295954
rect 534806 295718 534868 295954
rect 533868 295634 534868 295718
rect 533868 295398 533930 295634
rect 534166 295398 534250 295634
rect 534486 295398 534570 295634
rect 534806 295398 534868 295634
rect 533868 295366 534868 295398
rect 553868 295954 554868 295986
rect 553868 295718 553930 295954
rect 554166 295718 554250 295954
rect 554486 295718 554570 295954
rect 554806 295718 554868 295954
rect 553868 295634 554868 295718
rect 553868 295398 553930 295634
rect 554166 295398 554250 295634
rect 554486 295398 554570 295634
rect 554806 295398 554868 295634
rect 553868 295366 554868 295398
rect 303868 291454 304868 291486
rect 303868 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 304868 291454
rect 303868 291134 304868 291218
rect 303868 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 304868 291134
rect 303868 290866 304868 290898
rect 323868 291454 324868 291486
rect 323868 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 324868 291454
rect 323868 291134 324868 291218
rect 323868 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 324868 291134
rect 323868 290866 324868 290898
rect 343868 291454 344868 291486
rect 343868 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 344868 291454
rect 343868 291134 344868 291218
rect 343868 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 344868 291134
rect 343868 290866 344868 290898
rect 363868 291454 364868 291486
rect 363868 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 364868 291454
rect 363868 291134 364868 291218
rect 363868 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 364868 291134
rect 363868 290866 364868 290898
rect 383868 291454 384868 291486
rect 383868 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 384868 291454
rect 383868 291134 384868 291218
rect 383868 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 384868 291134
rect 383868 290866 384868 290898
rect 403868 291454 404868 291486
rect 403868 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 404868 291454
rect 403868 291134 404868 291218
rect 403868 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 404868 291134
rect 403868 290866 404868 290898
rect 423868 291454 424868 291486
rect 423868 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 424868 291454
rect 423868 291134 424868 291218
rect 423868 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 424868 291134
rect 423868 290866 424868 290898
rect 443868 291454 444868 291486
rect 443868 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 444868 291454
rect 443868 291134 444868 291218
rect 443868 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 444868 291134
rect 443868 290866 444868 290898
rect 463868 291454 464868 291486
rect 463868 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 464868 291454
rect 463868 291134 464868 291218
rect 463868 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 464868 291134
rect 463868 290866 464868 290898
rect 483868 291454 484868 291486
rect 483868 291218 483930 291454
rect 484166 291218 484250 291454
rect 484486 291218 484570 291454
rect 484806 291218 484868 291454
rect 483868 291134 484868 291218
rect 483868 290898 483930 291134
rect 484166 290898 484250 291134
rect 484486 290898 484570 291134
rect 484806 290898 484868 291134
rect 483868 290866 484868 290898
rect 503868 291454 504868 291486
rect 503868 291218 503930 291454
rect 504166 291218 504250 291454
rect 504486 291218 504570 291454
rect 504806 291218 504868 291454
rect 503868 291134 504868 291218
rect 503868 290898 503930 291134
rect 504166 290898 504250 291134
rect 504486 290898 504570 291134
rect 504806 290898 504868 291134
rect 503868 290866 504868 290898
rect 523868 291454 524868 291486
rect 523868 291218 523930 291454
rect 524166 291218 524250 291454
rect 524486 291218 524570 291454
rect 524806 291218 524868 291454
rect 523868 291134 524868 291218
rect 523868 290898 523930 291134
rect 524166 290898 524250 291134
rect 524486 290898 524570 291134
rect 524806 290898 524868 291134
rect 523868 290866 524868 290898
rect 543868 291454 544868 291486
rect 543868 291218 543930 291454
rect 544166 291218 544250 291454
rect 544486 291218 544570 291454
rect 544806 291218 544868 291454
rect 543868 291134 544868 291218
rect 543868 290898 543930 291134
rect 544166 290898 544250 291134
rect 544486 290898 544570 291134
rect 544806 290898 544868 291134
rect 543868 290866 544868 290898
rect 563868 291454 564868 291486
rect 563868 291218 563930 291454
rect 564166 291218 564250 291454
rect 564486 291218 564570 291454
rect 564806 291218 564868 291454
rect 563868 291134 564868 291218
rect 563868 290898 563930 291134
rect 564166 290898 564250 291134
rect 564486 290898 564570 291134
rect 564806 290898 564868 291134
rect 563868 290866 564868 290898
rect 313868 259954 314868 259986
rect 313868 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 314868 259954
rect 313868 259634 314868 259718
rect 313868 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 314868 259634
rect 313868 259366 314868 259398
rect 333868 259954 334868 259986
rect 333868 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 334868 259954
rect 333868 259634 334868 259718
rect 333868 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 334868 259634
rect 333868 259366 334868 259398
rect 353868 259954 354868 259986
rect 353868 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 354868 259954
rect 353868 259634 354868 259718
rect 353868 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 354868 259634
rect 353868 259366 354868 259398
rect 373868 259954 374868 259986
rect 373868 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 374868 259954
rect 373868 259634 374868 259718
rect 373868 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 374868 259634
rect 373868 259366 374868 259398
rect 393868 259954 394868 259986
rect 393868 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 394868 259954
rect 393868 259634 394868 259718
rect 393868 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 394868 259634
rect 393868 259366 394868 259398
rect 413868 259954 414868 259986
rect 413868 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 414868 259954
rect 413868 259634 414868 259718
rect 413868 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 414868 259634
rect 413868 259366 414868 259398
rect 433868 259954 434868 259986
rect 433868 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 434868 259954
rect 433868 259634 434868 259718
rect 433868 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 434868 259634
rect 433868 259366 434868 259398
rect 453868 259954 454868 259986
rect 453868 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 454868 259954
rect 453868 259634 454868 259718
rect 453868 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 454868 259634
rect 453868 259366 454868 259398
rect 473868 259954 474868 259986
rect 473868 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 474868 259954
rect 473868 259634 474868 259718
rect 473868 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 474868 259634
rect 473868 259366 474868 259398
rect 493868 259954 494868 259986
rect 493868 259718 493930 259954
rect 494166 259718 494250 259954
rect 494486 259718 494570 259954
rect 494806 259718 494868 259954
rect 493868 259634 494868 259718
rect 493868 259398 493930 259634
rect 494166 259398 494250 259634
rect 494486 259398 494570 259634
rect 494806 259398 494868 259634
rect 493868 259366 494868 259398
rect 513868 259954 514868 259986
rect 513868 259718 513930 259954
rect 514166 259718 514250 259954
rect 514486 259718 514570 259954
rect 514806 259718 514868 259954
rect 513868 259634 514868 259718
rect 513868 259398 513930 259634
rect 514166 259398 514250 259634
rect 514486 259398 514570 259634
rect 514806 259398 514868 259634
rect 513868 259366 514868 259398
rect 533868 259954 534868 259986
rect 533868 259718 533930 259954
rect 534166 259718 534250 259954
rect 534486 259718 534570 259954
rect 534806 259718 534868 259954
rect 533868 259634 534868 259718
rect 533868 259398 533930 259634
rect 534166 259398 534250 259634
rect 534486 259398 534570 259634
rect 534806 259398 534868 259634
rect 533868 259366 534868 259398
rect 553868 259954 554868 259986
rect 553868 259718 553930 259954
rect 554166 259718 554250 259954
rect 554486 259718 554570 259954
rect 554806 259718 554868 259954
rect 553868 259634 554868 259718
rect 553868 259398 553930 259634
rect 554166 259398 554250 259634
rect 554486 259398 554570 259634
rect 554806 259398 554868 259634
rect 553868 259366 554868 259398
rect 303868 255454 304868 255486
rect 303868 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 304868 255454
rect 303868 255134 304868 255218
rect 303868 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 304868 255134
rect 303868 254866 304868 254898
rect 323868 255454 324868 255486
rect 323868 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 324868 255454
rect 323868 255134 324868 255218
rect 323868 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 324868 255134
rect 323868 254866 324868 254898
rect 343868 255454 344868 255486
rect 343868 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 344868 255454
rect 343868 255134 344868 255218
rect 343868 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 344868 255134
rect 343868 254866 344868 254898
rect 363868 255454 364868 255486
rect 363868 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 364868 255454
rect 363868 255134 364868 255218
rect 363868 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 364868 255134
rect 363868 254866 364868 254898
rect 383868 255454 384868 255486
rect 383868 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 384868 255454
rect 383868 255134 384868 255218
rect 383868 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 384868 255134
rect 383868 254866 384868 254898
rect 403868 255454 404868 255486
rect 403868 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 404868 255454
rect 403868 255134 404868 255218
rect 403868 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 404868 255134
rect 403868 254866 404868 254898
rect 423868 255454 424868 255486
rect 423868 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 424868 255454
rect 423868 255134 424868 255218
rect 423868 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 424868 255134
rect 423868 254866 424868 254898
rect 443868 255454 444868 255486
rect 443868 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 444868 255454
rect 443868 255134 444868 255218
rect 443868 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 444868 255134
rect 443868 254866 444868 254898
rect 463868 255454 464868 255486
rect 463868 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 464868 255454
rect 463868 255134 464868 255218
rect 463868 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 464868 255134
rect 463868 254866 464868 254898
rect 483868 255454 484868 255486
rect 483868 255218 483930 255454
rect 484166 255218 484250 255454
rect 484486 255218 484570 255454
rect 484806 255218 484868 255454
rect 483868 255134 484868 255218
rect 483868 254898 483930 255134
rect 484166 254898 484250 255134
rect 484486 254898 484570 255134
rect 484806 254898 484868 255134
rect 483868 254866 484868 254898
rect 503868 255454 504868 255486
rect 503868 255218 503930 255454
rect 504166 255218 504250 255454
rect 504486 255218 504570 255454
rect 504806 255218 504868 255454
rect 503868 255134 504868 255218
rect 503868 254898 503930 255134
rect 504166 254898 504250 255134
rect 504486 254898 504570 255134
rect 504806 254898 504868 255134
rect 503868 254866 504868 254898
rect 523868 255454 524868 255486
rect 523868 255218 523930 255454
rect 524166 255218 524250 255454
rect 524486 255218 524570 255454
rect 524806 255218 524868 255454
rect 523868 255134 524868 255218
rect 523868 254898 523930 255134
rect 524166 254898 524250 255134
rect 524486 254898 524570 255134
rect 524806 254898 524868 255134
rect 523868 254866 524868 254898
rect 543868 255454 544868 255486
rect 543868 255218 543930 255454
rect 544166 255218 544250 255454
rect 544486 255218 544570 255454
rect 544806 255218 544868 255454
rect 543868 255134 544868 255218
rect 543868 254898 543930 255134
rect 544166 254898 544250 255134
rect 544486 254898 544570 255134
rect 544806 254898 544868 255134
rect 543868 254866 544868 254898
rect 563868 255454 564868 255486
rect 563868 255218 563930 255454
rect 564166 255218 564250 255454
rect 564486 255218 564570 255454
rect 564806 255218 564868 255454
rect 563868 255134 564868 255218
rect 563868 254898 563930 255134
rect 564166 254898 564250 255134
rect 564486 254898 564570 255134
rect 564806 254898 564868 255134
rect 563868 254866 564868 254898
rect 313868 223954 314868 223986
rect 313868 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 314868 223954
rect 313868 223634 314868 223718
rect 313868 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 314868 223634
rect 313868 223366 314868 223398
rect 333868 223954 334868 223986
rect 333868 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 334868 223954
rect 333868 223634 334868 223718
rect 333868 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 334868 223634
rect 333868 223366 334868 223398
rect 353868 223954 354868 223986
rect 353868 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 354868 223954
rect 353868 223634 354868 223718
rect 353868 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 354868 223634
rect 353868 223366 354868 223398
rect 373868 223954 374868 223986
rect 373868 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 374868 223954
rect 373868 223634 374868 223718
rect 373868 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 374868 223634
rect 373868 223366 374868 223398
rect 393868 223954 394868 223986
rect 393868 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 394868 223954
rect 393868 223634 394868 223718
rect 393868 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 394868 223634
rect 393868 223366 394868 223398
rect 413868 223954 414868 223986
rect 413868 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 414868 223954
rect 413868 223634 414868 223718
rect 413868 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 414868 223634
rect 413868 223366 414868 223398
rect 433868 223954 434868 223986
rect 433868 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 434868 223954
rect 433868 223634 434868 223718
rect 433868 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 434868 223634
rect 433868 223366 434868 223398
rect 453868 223954 454868 223986
rect 453868 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 454868 223954
rect 453868 223634 454868 223718
rect 453868 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 454868 223634
rect 453868 223366 454868 223398
rect 473868 223954 474868 223986
rect 473868 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 474868 223954
rect 473868 223634 474868 223718
rect 473868 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 474868 223634
rect 473868 223366 474868 223398
rect 493868 223954 494868 223986
rect 493868 223718 493930 223954
rect 494166 223718 494250 223954
rect 494486 223718 494570 223954
rect 494806 223718 494868 223954
rect 493868 223634 494868 223718
rect 493868 223398 493930 223634
rect 494166 223398 494250 223634
rect 494486 223398 494570 223634
rect 494806 223398 494868 223634
rect 493868 223366 494868 223398
rect 513868 223954 514868 223986
rect 513868 223718 513930 223954
rect 514166 223718 514250 223954
rect 514486 223718 514570 223954
rect 514806 223718 514868 223954
rect 513868 223634 514868 223718
rect 513868 223398 513930 223634
rect 514166 223398 514250 223634
rect 514486 223398 514570 223634
rect 514806 223398 514868 223634
rect 513868 223366 514868 223398
rect 533868 223954 534868 223986
rect 533868 223718 533930 223954
rect 534166 223718 534250 223954
rect 534486 223718 534570 223954
rect 534806 223718 534868 223954
rect 533868 223634 534868 223718
rect 533868 223398 533930 223634
rect 534166 223398 534250 223634
rect 534486 223398 534570 223634
rect 534806 223398 534868 223634
rect 533868 223366 534868 223398
rect 553868 223954 554868 223986
rect 553868 223718 553930 223954
rect 554166 223718 554250 223954
rect 554486 223718 554570 223954
rect 554806 223718 554868 223954
rect 553868 223634 554868 223718
rect 553868 223398 553930 223634
rect 554166 223398 554250 223634
rect 554486 223398 554570 223634
rect 554806 223398 554868 223634
rect 553868 223366 554868 223398
rect 303868 219454 304868 219486
rect 303868 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 304868 219454
rect 303868 219134 304868 219218
rect 303868 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 304868 219134
rect 303868 218866 304868 218898
rect 323868 219454 324868 219486
rect 323868 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 324868 219454
rect 323868 219134 324868 219218
rect 323868 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 324868 219134
rect 323868 218866 324868 218898
rect 343868 219454 344868 219486
rect 343868 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 344868 219454
rect 343868 219134 344868 219218
rect 343868 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 344868 219134
rect 343868 218866 344868 218898
rect 363868 219454 364868 219486
rect 363868 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 364868 219454
rect 363868 219134 364868 219218
rect 363868 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 364868 219134
rect 363868 218866 364868 218898
rect 383868 219454 384868 219486
rect 383868 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 384868 219454
rect 383868 219134 384868 219218
rect 383868 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 384868 219134
rect 383868 218866 384868 218898
rect 403868 219454 404868 219486
rect 403868 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 404868 219454
rect 403868 219134 404868 219218
rect 403868 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 404868 219134
rect 403868 218866 404868 218898
rect 423868 219454 424868 219486
rect 423868 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 424868 219454
rect 423868 219134 424868 219218
rect 423868 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 424868 219134
rect 423868 218866 424868 218898
rect 443868 219454 444868 219486
rect 443868 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 444868 219454
rect 443868 219134 444868 219218
rect 443868 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 444868 219134
rect 443868 218866 444868 218898
rect 463868 219454 464868 219486
rect 463868 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 464868 219454
rect 463868 219134 464868 219218
rect 463868 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 464868 219134
rect 463868 218866 464868 218898
rect 483868 219454 484868 219486
rect 483868 219218 483930 219454
rect 484166 219218 484250 219454
rect 484486 219218 484570 219454
rect 484806 219218 484868 219454
rect 483868 219134 484868 219218
rect 483868 218898 483930 219134
rect 484166 218898 484250 219134
rect 484486 218898 484570 219134
rect 484806 218898 484868 219134
rect 483868 218866 484868 218898
rect 503868 219454 504868 219486
rect 503868 219218 503930 219454
rect 504166 219218 504250 219454
rect 504486 219218 504570 219454
rect 504806 219218 504868 219454
rect 503868 219134 504868 219218
rect 503868 218898 503930 219134
rect 504166 218898 504250 219134
rect 504486 218898 504570 219134
rect 504806 218898 504868 219134
rect 503868 218866 504868 218898
rect 523868 219454 524868 219486
rect 523868 219218 523930 219454
rect 524166 219218 524250 219454
rect 524486 219218 524570 219454
rect 524806 219218 524868 219454
rect 523868 219134 524868 219218
rect 523868 218898 523930 219134
rect 524166 218898 524250 219134
rect 524486 218898 524570 219134
rect 524806 218898 524868 219134
rect 523868 218866 524868 218898
rect 543868 219454 544868 219486
rect 543868 219218 543930 219454
rect 544166 219218 544250 219454
rect 544486 219218 544570 219454
rect 544806 219218 544868 219454
rect 543868 219134 544868 219218
rect 543868 218898 543930 219134
rect 544166 218898 544250 219134
rect 544486 218898 544570 219134
rect 544806 218898 544868 219134
rect 543868 218866 544868 218898
rect 563868 219454 564868 219486
rect 563868 219218 563930 219454
rect 564166 219218 564250 219454
rect 564486 219218 564570 219454
rect 564806 219218 564868 219454
rect 563868 219134 564868 219218
rect 563868 218898 563930 219134
rect 564166 218898 564250 219134
rect 564486 218898 564570 219134
rect 564806 218898 564868 219134
rect 563868 218866 564868 218898
rect 302739 201380 302805 201381
rect 302739 201316 302740 201380
rect 302804 201316 302805 201380
rect 302739 201315 302805 201316
rect 302742 200130 302802 201315
rect 302742 200070 303538 200130
rect 303478 59261 303538 200070
rect 565862 187645 565922 332283
rect 567702 315757 567762 461075
rect 567886 459373 567946 571915
rect 568622 463589 568682 580211
rect 568619 463588 568685 463589
rect 568619 463524 568620 463588
rect 568684 463524 568685 463588
rect 568619 463523 568685 463524
rect 567883 459372 567949 459373
rect 567883 459308 567884 459372
rect 567948 459308 567949 459372
rect 567883 459307 567949 459308
rect 568435 336700 568501 336701
rect 568435 336636 568436 336700
rect 568500 336636 568501 336700
rect 568435 336635 568501 336636
rect 567699 315756 567765 315757
rect 567699 315692 567700 315756
rect 567764 315692 567765 315756
rect 567699 315691 567765 315692
rect 567702 209790 567762 315691
rect 568438 314669 568498 336635
rect 568435 314668 568501 314669
rect 568435 314604 568436 314668
rect 568500 314604 568501 314668
rect 568435 314603 568501 314604
rect 567334 209730 567762 209790
rect 567334 204373 567394 209730
rect 567331 204372 567397 204373
rect 567331 204308 567332 204372
rect 567396 204308 567397 204372
rect 567331 204307 567397 204308
rect 567334 202890 567394 204307
rect 566966 202830 567394 202890
rect 565859 187644 565925 187645
rect 565859 187580 565860 187644
rect 565924 187580 565925 187644
rect 565859 187579 565925 187580
rect 303868 183454 304868 183486
rect 303868 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 304868 183454
rect 303868 183134 304868 183218
rect 303868 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 304868 183134
rect 303868 182866 304868 182898
rect 323868 183454 324868 183486
rect 323868 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 324868 183454
rect 323868 183134 324868 183218
rect 323868 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 324868 183134
rect 323868 182866 324868 182898
rect 343868 183454 344868 183486
rect 343868 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 344868 183454
rect 343868 183134 344868 183218
rect 343868 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 344868 183134
rect 343868 182866 344868 182898
rect 363868 183454 364868 183486
rect 363868 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 364868 183454
rect 363868 183134 364868 183218
rect 363868 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 364868 183134
rect 363868 182866 364868 182898
rect 383868 183454 384868 183486
rect 383868 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 384868 183454
rect 383868 183134 384868 183218
rect 383868 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 384868 183134
rect 383868 182866 384868 182898
rect 403868 183454 404868 183486
rect 403868 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 404868 183454
rect 403868 183134 404868 183218
rect 403868 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 404868 183134
rect 403868 182866 404868 182898
rect 423868 183454 424868 183486
rect 423868 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 424868 183454
rect 423868 183134 424868 183218
rect 423868 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 424868 183134
rect 423868 182866 424868 182898
rect 443868 183454 444868 183486
rect 443868 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 444868 183454
rect 443868 183134 444868 183218
rect 443868 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 444868 183134
rect 443868 182866 444868 182898
rect 463868 183454 464868 183486
rect 463868 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 464868 183454
rect 463868 183134 464868 183218
rect 463868 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 464868 183134
rect 463868 182866 464868 182898
rect 483868 183454 484868 183486
rect 483868 183218 483930 183454
rect 484166 183218 484250 183454
rect 484486 183218 484570 183454
rect 484806 183218 484868 183454
rect 483868 183134 484868 183218
rect 483868 182898 483930 183134
rect 484166 182898 484250 183134
rect 484486 182898 484570 183134
rect 484806 182898 484868 183134
rect 483868 182866 484868 182898
rect 503868 183454 504868 183486
rect 503868 183218 503930 183454
rect 504166 183218 504250 183454
rect 504486 183218 504570 183454
rect 504806 183218 504868 183454
rect 503868 183134 504868 183218
rect 503868 182898 503930 183134
rect 504166 182898 504250 183134
rect 504486 182898 504570 183134
rect 504806 182898 504868 183134
rect 503868 182866 504868 182898
rect 523868 183454 524868 183486
rect 523868 183218 523930 183454
rect 524166 183218 524250 183454
rect 524486 183218 524570 183454
rect 524806 183218 524868 183454
rect 523868 183134 524868 183218
rect 523868 182898 523930 183134
rect 524166 182898 524250 183134
rect 524486 182898 524570 183134
rect 524806 182898 524868 183134
rect 523868 182866 524868 182898
rect 543868 183454 544868 183486
rect 543868 183218 543930 183454
rect 544166 183218 544250 183454
rect 544486 183218 544570 183454
rect 544806 183218 544868 183454
rect 543868 183134 544868 183218
rect 543868 182898 543930 183134
rect 544166 182898 544250 183134
rect 544486 182898 544570 183134
rect 544806 182898 544868 183134
rect 543868 182866 544868 182898
rect 563868 183454 564868 183486
rect 563868 183218 563930 183454
rect 564166 183218 564250 183454
rect 564486 183218 564570 183454
rect 564806 183218 564868 183454
rect 563868 183134 564868 183218
rect 563868 182898 563930 183134
rect 564166 182898 564250 183134
rect 564486 182898 564570 183134
rect 564806 182898 564868 183134
rect 563868 182866 564868 182898
rect 313868 151954 314868 151986
rect 313868 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 314868 151954
rect 313868 151634 314868 151718
rect 313868 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 314868 151634
rect 313868 151366 314868 151398
rect 333868 151954 334868 151986
rect 333868 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 334868 151954
rect 333868 151634 334868 151718
rect 333868 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 334868 151634
rect 333868 151366 334868 151398
rect 353868 151954 354868 151986
rect 353868 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 354868 151954
rect 353868 151634 354868 151718
rect 353868 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 354868 151634
rect 353868 151366 354868 151398
rect 373868 151954 374868 151986
rect 373868 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 374868 151954
rect 373868 151634 374868 151718
rect 373868 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 374868 151634
rect 373868 151366 374868 151398
rect 393868 151954 394868 151986
rect 393868 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 394868 151954
rect 393868 151634 394868 151718
rect 393868 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 394868 151634
rect 393868 151366 394868 151398
rect 413868 151954 414868 151986
rect 413868 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 414868 151954
rect 413868 151634 414868 151718
rect 413868 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 414868 151634
rect 413868 151366 414868 151398
rect 433868 151954 434868 151986
rect 433868 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 434868 151954
rect 433868 151634 434868 151718
rect 433868 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 434868 151634
rect 433868 151366 434868 151398
rect 453868 151954 454868 151986
rect 453868 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 454868 151954
rect 453868 151634 454868 151718
rect 453868 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 454868 151634
rect 453868 151366 454868 151398
rect 473868 151954 474868 151986
rect 473868 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 474868 151954
rect 473868 151634 474868 151718
rect 473868 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 474868 151634
rect 473868 151366 474868 151398
rect 493868 151954 494868 151986
rect 493868 151718 493930 151954
rect 494166 151718 494250 151954
rect 494486 151718 494570 151954
rect 494806 151718 494868 151954
rect 493868 151634 494868 151718
rect 493868 151398 493930 151634
rect 494166 151398 494250 151634
rect 494486 151398 494570 151634
rect 494806 151398 494868 151634
rect 493868 151366 494868 151398
rect 513868 151954 514868 151986
rect 513868 151718 513930 151954
rect 514166 151718 514250 151954
rect 514486 151718 514570 151954
rect 514806 151718 514868 151954
rect 513868 151634 514868 151718
rect 513868 151398 513930 151634
rect 514166 151398 514250 151634
rect 514486 151398 514570 151634
rect 514806 151398 514868 151634
rect 513868 151366 514868 151398
rect 533868 151954 534868 151986
rect 533868 151718 533930 151954
rect 534166 151718 534250 151954
rect 534486 151718 534570 151954
rect 534806 151718 534868 151954
rect 533868 151634 534868 151718
rect 533868 151398 533930 151634
rect 534166 151398 534250 151634
rect 534486 151398 534570 151634
rect 534806 151398 534868 151634
rect 533868 151366 534868 151398
rect 553868 151954 554868 151986
rect 553868 151718 553930 151954
rect 554166 151718 554250 151954
rect 554486 151718 554570 151954
rect 554806 151718 554868 151954
rect 553868 151634 554868 151718
rect 553868 151398 553930 151634
rect 554166 151398 554250 151634
rect 554486 151398 554570 151634
rect 554806 151398 554868 151634
rect 553868 151366 554868 151398
rect 303868 147454 304868 147486
rect 303868 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 304868 147454
rect 303868 147134 304868 147218
rect 303868 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 304868 147134
rect 303868 146866 304868 146898
rect 323868 147454 324868 147486
rect 323868 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 324868 147454
rect 323868 147134 324868 147218
rect 323868 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 324868 147134
rect 323868 146866 324868 146898
rect 343868 147454 344868 147486
rect 343868 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 344868 147454
rect 343868 147134 344868 147218
rect 343868 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 344868 147134
rect 343868 146866 344868 146898
rect 363868 147454 364868 147486
rect 363868 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 364868 147454
rect 363868 147134 364868 147218
rect 363868 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 364868 147134
rect 363868 146866 364868 146898
rect 383868 147454 384868 147486
rect 383868 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 384868 147454
rect 383868 147134 384868 147218
rect 383868 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 384868 147134
rect 383868 146866 384868 146898
rect 403868 147454 404868 147486
rect 403868 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 404868 147454
rect 403868 147134 404868 147218
rect 403868 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 404868 147134
rect 403868 146866 404868 146898
rect 423868 147454 424868 147486
rect 423868 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 424868 147454
rect 423868 147134 424868 147218
rect 423868 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 424868 147134
rect 423868 146866 424868 146898
rect 443868 147454 444868 147486
rect 443868 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 444868 147454
rect 443868 147134 444868 147218
rect 443868 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 444868 147134
rect 443868 146866 444868 146898
rect 463868 147454 464868 147486
rect 463868 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 464868 147454
rect 463868 147134 464868 147218
rect 463868 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 464868 147134
rect 463868 146866 464868 146898
rect 483868 147454 484868 147486
rect 483868 147218 483930 147454
rect 484166 147218 484250 147454
rect 484486 147218 484570 147454
rect 484806 147218 484868 147454
rect 483868 147134 484868 147218
rect 483868 146898 483930 147134
rect 484166 146898 484250 147134
rect 484486 146898 484570 147134
rect 484806 146898 484868 147134
rect 483868 146866 484868 146898
rect 503868 147454 504868 147486
rect 503868 147218 503930 147454
rect 504166 147218 504250 147454
rect 504486 147218 504570 147454
rect 504806 147218 504868 147454
rect 503868 147134 504868 147218
rect 503868 146898 503930 147134
rect 504166 146898 504250 147134
rect 504486 146898 504570 147134
rect 504806 146898 504868 147134
rect 503868 146866 504868 146898
rect 523868 147454 524868 147486
rect 523868 147218 523930 147454
rect 524166 147218 524250 147454
rect 524486 147218 524570 147454
rect 524806 147218 524868 147454
rect 523868 147134 524868 147218
rect 523868 146898 523930 147134
rect 524166 146898 524250 147134
rect 524486 146898 524570 147134
rect 524806 146898 524868 147134
rect 523868 146866 524868 146898
rect 543868 147454 544868 147486
rect 543868 147218 543930 147454
rect 544166 147218 544250 147454
rect 544486 147218 544570 147454
rect 544806 147218 544868 147454
rect 543868 147134 544868 147218
rect 543868 146898 543930 147134
rect 544166 146898 544250 147134
rect 544486 146898 544570 147134
rect 544806 146898 544868 147134
rect 543868 146866 544868 146898
rect 563868 147454 564868 147486
rect 563868 147218 563930 147454
rect 564166 147218 564250 147454
rect 564486 147218 564570 147454
rect 564806 147218 564868 147454
rect 563868 147134 564868 147218
rect 563868 146898 563930 147134
rect 564166 146898 564250 147134
rect 564486 146898 564570 147134
rect 564806 146898 564868 147134
rect 563868 146866 564868 146898
rect 313868 115954 314868 115986
rect 313868 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 314868 115954
rect 313868 115634 314868 115718
rect 313868 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 314868 115634
rect 313868 115366 314868 115398
rect 333868 115954 334868 115986
rect 333868 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 334868 115954
rect 333868 115634 334868 115718
rect 333868 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 334868 115634
rect 333868 115366 334868 115398
rect 353868 115954 354868 115986
rect 353868 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 354868 115954
rect 353868 115634 354868 115718
rect 353868 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 354868 115634
rect 353868 115366 354868 115398
rect 373868 115954 374868 115986
rect 373868 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 374868 115954
rect 373868 115634 374868 115718
rect 373868 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 374868 115634
rect 373868 115366 374868 115398
rect 393868 115954 394868 115986
rect 393868 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 394868 115954
rect 393868 115634 394868 115718
rect 393868 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 394868 115634
rect 393868 115366 394868 115398
rect 413868 115954 414868 115986
rect 413868 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 414868 115954
rect 413868 115634 414868 115718
rect 413868 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 414868 115634
rect 413868 115366 414868 115398
rect 433868 115954 434868 115986
rect 433868 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 434868 115954
rect 433868 115634 434868 115718
rect 433868 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 434868 115634
rect 433868 115366 434868 115398
rect 453868 115954 454868 115986
rect 453868 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 454868 115954
rect 453868 115634 454868 115718
rect 453868 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 454868 115634
rect 453868 115366 454868 115398
rect 473868 115954 474868 115986
rect 473868 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 474868 115954
rect 473868 115634 474868 115718
rect 473868 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 474868 115634
rect 473868 115366 474868 115398
rect 493868 115954 494868 115986
rect 493868 115718 493930 115954
rect 494166 115718 494250 115954
rect 494486 115718 494570 115954
rect 494806 115718 494868 115954
rect 493868 115634 494868 115718
rect 493868 115398 493930 115634
rect 494166 115398 494250 115634
rect 494486 115398 494570 115634
rect 494806 115398 494868 115634
rect 493868 115366 494868 115398
rect 513868 115954 514868 115986
rect 513868 115718 513930 115954
rect 514166 115718 514250 115954
rect 514486 115718 514570 115954
rect 514806 115718 514868 115954
rect 513868 115634 514868 115718
rect 513868 115398 513930 115634
rect 514166 115398 514250 115634
rect 514486 115398 514570 115634
rect 514806 115398 514868 115634
rect 513868 115366 514868 115398
rect 533868 115954 534868 115986
rect 533868 115718 533930 115954
rect 534166 115718 534250 115954
rect 534486 115718 534570 115954
rect 534806 115718 534868 115954
rect 533868 115634 534868 115718
rect 533868 115398 533930 115634
rect 534166 115398 534250 115634
rect 534486 115398 534570 115634
rect 534806 115398 534868 115634
rect 533868 115366 534868 115398
rect 553868 115954 554868 115986
rect 553868 115718 553930 115954
rect 554166 115718 554250 115954
rect 554486 115718 554570 115954
rect 554806 115718 554868 115954
rect 553868 115634 554868 115718
rect 553868 115398 553930 115634
rect 554166 115398 554250 115634
rect 554486 115398 554570 115634
rect 554806 115398 554868 115634
rect 553868 115366 554868 115398
rect 303868 111454 304868 111486
rect 303868 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 304868 111454
rect 303868 111134 304868 111218
rect 303868 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 304868 111134
rect 303868 110866 304868 110898
rect 323868 111454 324868 111486
rect 323868 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 324868 111454
rect 323868 111134 324868 111218
rect 323868 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 324868 111134
rect 323868 110866 324868 110898
rect 343868 111454 344868 111486
rect 343868 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 344868 111454
rect 343868 111134 344868 111218
rect 343868 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 344868 111134
rect 343868 110866 344868 110898
rect 363868 111454 364868 111486
rect 363868 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 364868 111454
rect 363868 111134 364868 111218
rect 363868 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 364868 111134
rect 363868 110866 364868 110898
rect 383868 111454 384868 111486
rect 383868 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 384868 111454
rect 383868 111134 384868 111218
rect 383868 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 384868 111134
rect 383868 110866 384868 110898
rect 403868 111454 404868 111486
rect 403868 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 404868 111454
rect 403868 111134 404868 111218
rect 403868 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 404868 111134
rect 403868 110866 404868 110898
rect 423868 111454 424868 111486
rect 423868 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 424868 111454
rect 423868 111134 424868 111218
rect 423868 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 424868 111134
rect 423868 110866 424868 110898
rect 443868 111454 444868 111486
rect 443868 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 444868 111454
rect 443868 111134 444868 111218
rect 443868 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 444868 111134
rect 443868 110866 444868 110898
rect 463868 111454 464868 111486
rect 463868 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 464868 111454
rect 463868 111134 464868 111218
rect 463868 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 464868 111134
rect 463868 110866 464868 110898
rect 483868 111454 484868 111486
rect 483868 111218 483930 111454
rect 484166 111218 484250 111454
rect 484486 111218 484570 111454
rect 484806 111218 484868 111454
rect 483868 111134 484868 111218
rect 483868 110898 483930 111134
rect 484166 110898 484250 111134
rect 484486 110898 484570 111134
rect 484806 110898 484868 111134
rect 483868 110866 484868 110898
rect 503868 111454 504868 111486
rect 503868 111218 503930 111454
rect 504166 111218 504250 111454
rect 504486 111218 504570 111454
rect 504806 111218 504868 111454
rect 503868 111134 504868 111218
rect 503868 110898 503930 111134
rect 504166 110898 504250 111134
rect 504486 110898 504570 111134
rect 504806 110898 504868 111134
rect 503868 110866 504868 110898
rect 523868 111454 524868 111486
rect 523868 111218 523930 111454
rect 524166 111218 524250 111454
rect 524486 111218 524570 111454
rect 524806 111218 524868 111454
rect 523868 111134 524868 111218
rect 523868 110898 523930 111134
rect 524166 110898 524250 111134
rect 524486 110898 524570 111134
rect 524806 110898 524868 111134
rect 523868 110866 524868 110898
rect 543868 111454 544868 111486
rect 543868 111218 543930 111454
rect 544166 111218 544250 111454
rect 544486 111218 544570 111454
rect 544806 111218 544868 111454
rect 543868 111134 544868 111218
rect 543868 110898 543930 111134
rect 544166 110898 544250 111134
rect 544486 110898 544570 111134
rect 544806 110898 544868 111134
rect 543868 110866 544868 110898
rect 563868 111454 564868 111486
rect 563868 111218 563930 111454
rect 564166 111218 564250 111454
rect 564486 111218 564570 111454
rect 564806 111218 564868 111454
rect 563868 111134 564868 111218
rect 563868 110898 563930 111134
rect 564166 110898 564250 111134
rect 564486 110898 564570 111134
rect 564806 110898 564868 111134
rect 563868 110866 564868 110898
rect 303659 80204 303725 80205
rect 303659 80140 303660 80204
rect 303724 80140 303725 80204
rect 303659 80139 303725 80140
rect 303662 61437 303722 80139
rect 303659 61436 303725 61437
rect 303659 61372 303660 61436
rect 303724 61372 303725 61436
rect 303659 61371 303725 61372
rect 303475 59260 303541 59261
rect 303475 59196 303476 59260
rect 303540 59196 303541 59260
rect 303475 59195 303541 59196
rect 302003 58580 302069 58581
rect 302003 58516 302004 58580
rect 302068 58516 302069 58580
rect 302003 58515 302069 58516
rect 297219 57220 297285 57221
rect 297219 57156 297220 57220
rect 297284 57156 297285 57220
rect 297219 57155 297285 57156
rect 295931 54500 295997 54501
rect 295931 54436 295932 54500
rect 295996 54436 295997 54500
rect 295931 54435 295997 54436
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 213868 43954 214868 43986
rect 213868 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 214868 43954
rect 213868 43634 214868 43718
rect 213868 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 214868 43634
rect 213868 43366 214868 43398
rect 233868 43954 234868 43986
rect 233868 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 234868 43954
rect 233868 43634 234868 43718
rect 233868 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 234868 43634
rect 233868 43366 234868 43398
rect 253868 43954 254868 43986
rect 253868 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 254868 43954
rect 253868 43634 254868 43718
rect 253868 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 254868 43634
rect 253868 43366 254868 43398
rect 273868 43954 274868 43986
rect 273868 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 274868 43954
rect 273868 43634 274868 43718
rect 273868 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 274868 43634
rect 273868 43366 274868 43398
rect 293868 43954 294868 43986
rect 293868 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 294868 43954
rect 293868 43634 294868 43718
rect 293868 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 294868 43634
rect 293868 43366 294868 43398
rect 313868 43954 314868 43986
rect 313868 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 314868 43954
rect 313868 43634 314868 43718
rect 313868 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 314868 43634
rect 313868 43366 314868 43398
rect 333868 43954 334868 43986
rect 333868 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 334868 43954
rect 333868 43634 334868 43718
rect 333868 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 334868 43634
rect 333868 43366 334868 43398
rect 353868 43954 354868 43986
rect 353868 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 354868 43954
rect 353868 43634 354868 43718
rect 353868 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 354868 43634
rect 353868 43366 354868 43398
rect 373868 43954 374868 43986
rect 373868 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 374868 43954
rect 373868 43634 374868 43718
rect 373868 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 374868 43634
rect 373868 43366 374868 43398
rect 393868 43954 394868 43986
rect 393868 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 394868 43954
rect 393868 43634 394868 43718
rect 393868 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 394868 43634
rect 393868 43366 394868 43398
rect 402294 43954 402914 76000
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 203868 39454 204868 39486
rect 203868 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 204868 39454
rect 203868 39134 204868 39218
rect 203868 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 204868 39134
rect 203868 38866 204868 38898
rect 223868 39454 224868 39486
rect 223868 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 224868 39454
rect 223868 39134 224868 39218
rect 223868 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 224868 39134
rect 223868 38866 224868 38898
rect 243868 39454 244868 39486
rect 243868 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 244868 39454
rect 243868 39134 244868 39218
rect 243868 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 244868 39134
rect 243868 38866 244868 38898
rect 263868 39454 264868 39486
rect 263868 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 264868 39454
rect 263868 39134 264868 39218
rect 263868 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 264868 39134
rect 263868 38866 264868 38898
rect 283868 39454 284868 39486
rect 283868 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 284868 39454
rect 283868 39134 284868 39218
rect 283868 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 284868 39134
rect 283868 38866 284868 38898
rect 303868 39454 304868 39486
rect 303868 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 304868 39454
rect 303868 39134 304868 39218
rect 303868 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 304868 39134
rect 303868 38866 304868 38898
rect 323868 39454 324868 39486
rect 323868 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 324868 39454
rect 323868 39134 324868 39218
rect 323868 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 324868 39134
rect 323868 38866 324868 38898
rect 343868 39454 344868 39486
rect 343868 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 344868 39454
rect 343868 39134 344868 39218
rect 343868 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 344868 39134
rect 343868 38866 344868 38898
rect 363868 39454 364868 39486
rect 363868 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 364868 39454
rect 363868 39134 364868 39218
rect 363868 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 364868 39134
rect 363868 38866 364868 38898
rect 383868 39454 384868 39486
rect 383868 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 384868 39454
rect 383868 39134 384868 39218
rect 383868 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 384868 39134
rect 383868 38866 384868 38898
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 22000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 217794 3454 218414 22000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7954 222914 22000
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 12454 227414 22000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 16954 231914 22000
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 21454 236414 22000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 253794 3454 254414 22000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 7954 258914 22000
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 12454 263414 22000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 22000
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 21454 272414 22000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 289794 3454 290414 22000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 22000
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 22000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 22000
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 22000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 325794 3454 326414 22000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 7954 330914 22000
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 12454 335414 22000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 16954 339914 22000
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 21454 344414 22000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 361794 3454 362414 22000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 7954 366914 22000
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 12454 371414 22000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 16954 375914 22000
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 21454 380414 22000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 397794 3454 398414 22000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 48454 407414 76000
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 52954 411914 76000
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 57454 416414 76000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 61954 420914 76000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 76000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 70954 429914 76000
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 75454 434414 76000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 43954 438914 76000
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 48454 443414 76000
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 52954 447914 76000
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 57454 452414 76000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 76000
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 66454 461414 76000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 70954 465914 76000
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 75454 470414 76000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 43954 474914 76000
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 48454 479414 76000
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 52954 483914 76000
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 57454 488414 76000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 61954 492914 76000
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 66454 497414 76000
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 70954 501914 76000
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 75454 506414 76000
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 43954 510914 76000
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 48454 515414 76000
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 52954 519914 76000
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 57454 524414 76000
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 61954 528914 76000
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 66454 533414 76000
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 70954 537914 76000
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 75454 542414 76000
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 43954 546914 76000
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 48454 551414 76000
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 52954 555914 76000
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 57454 560414 76000
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 61954 564914 76000
rect 565862 75853 565922 187579
rect 565859 75852 565925 75853
rect 565859 75788 565860 75852
rect 565924 75788 565925 75852
rect 565859 75787 565925 75788
rect 566966 74493 567026 202830
rect 566963 74492 567029 74493
rect 566963 74428 566964 74492
rect 567028 74428 567029 74492
rect 566963 74427 567029 74428
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 66454 569414 76000
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 569542 22133 569602 590955
rect 570091 585852 570157 585853
rect 570091 585788 570092 585852
rect 570156 585788 570157 585852
rect 570091 585787 570157 585788
rect 570094 76669 570154 585787
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 571379 458828 571445 458829
rect 571379 458764 571380 458828
rect 571444 458764 571445 458828
rect 571379 458763 571445 458764
rect 570459 418300 570525 418301
rect 570459 418236 570460 418300
rect 570524 418236 570525 418300
rect 570459 418235 570525 418236
rect 570091 76668 570157 76669
rect 570091 76604 570092 76668
rect 570156 76604 570157 76668
rect 570091 76603 570157 76604
rect 570462 75989 570522 418235
rect 571382 76533 571442 458763
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 571379 76532 571445 76533
rect 571379 76468 571380 76532
rect 571444 76468 571445 76532
rect 571379 76467 571445 76468
rect 570459 75988 570525 75989
rect 570459 75924 570460 75988
rect 570524 75924 570525 75988
rect 570459 75923 570525 75924
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 569539 22132 569605 22133
rect 569539 22068 569540 22132
rect 569604 22068 569605 22132
rect 569539 22067 569605 22068
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 33930 691718 34166 691954
rect 34250 691718 34486 691954
rect 34570 691718 34806 691954
rect 33930 691398 34166 691634
rect 34250 691398 34486 691634
rect 34570 691398 34806 691634
rect 53930 691718 54166 691954
rect 54250 691718 54486 691954
rect 54570 691718 54806 691954
rect 53930 691398 54166 691634
rect 54250 691398 54486 691634
rect 54570 691398 54806 691634
rect 73930 691718 74166 691954
rect 74250 691718 74486 691954
rect 74570 691718 74806 691954
rect 73930 691398 74166 691634
rect 74250 691398 74486 691634
rect 74570 691398 74806 691634
rect 93930 691718 94166 691954
rect 94250 691718 94486 691954
rect 94570 691718 94806 691954
rect 93930 691398 94166 691634
rect 94250 691398 94486 691634
rect 94570 691398 94806 691634
rect 113930 691718 114166 691954
rect 114250 691718 114486 691954
rect 114570 691718 114806 691954
rect 113930 691398 114166 691634
rect 114250 691398 114486 691634
rect 114570 691398 114806 691634
rect 133930 691718 134166 691954
rect 134250 691718 134486 691954
rect 134570 691718 134806 691954
rect 133930 691398 134166 691634
rect 134250 691398 134486 691634
rect 134570 691398 134806 691634
rect 153930 691718 154166 691954
rect 154250 691718 154486 691954
rect 154570 691718 154806 691954
rect 153930 691398 154166 691634
rect 154250 691398 154486 691634
rect 154570 691398 154806 691634
rect 173930 691718 174166 691954
rect 174250 691718 174486 691954
rect 174570 691718 174806 691954
rect 173930 691398 174166 691634
rect 174250 691398 174486 691634
rect 174570 691398 174806 691634
rect 193930 691718 194166 691954
rect 194250 691718 194486 691954
rect 194570 691718 194806 691954
rect 193930 691398 194166 691634
rect 194250 691398 194486 691634
rect 194570 691398 194806 691634
rect 213930 691718 214166 691954
rect 214250 691718 214486 691954
rect 214570 691718 214806 691954
rect 213930 691398 214166 691634
rect 214250 691398 214486 691634
rect 214570 691398 214806 691634
rect 233930 691718 234166 691954
rect 234250 691718 234486 691954
rect 234570 691718 234806 691954
rect 233930 691398 234166 691634
rect 234250 691398 234486 691634
rect 234570 691398 234806 691634
rect 253930 691718 254166 691954
rect 254250 691718 254486 691954
rect 254570 691718 254806 691954
rect 253930 691398 254166 691634
rect 254250 691398 254486 691634
rect 254570 691398 254806 691634
rect 273930 691718 274166 691954
rect 274250 691718 274486 691954
rect 274570 691718 274806 691954
rect 273930 691398 274166 691634
rect 274250 691398 274486 691634
rect 274570 691398 274806 691634
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 23930 687218 24166 687454
rect 24250 687218 24486 687454
rect 24570 687218 24806 687454
rect 23930 686898 24166 687134
rect 24250 686898 24486 687134
rect 24570 686898 24806 687134
rect 43930 687218 44166 687454
rect 44250 687218 44486 687454
rect 44570 687218 44806 687454
rect 43930 686898 44166 687134
rect 44250 686898 44486 687134
rect 44570 686898 44806 687134
rect 63930 687218 64166 687454
rect 64250 687218 64486 687454
rect 64570 687218 64806 687454
rect 63930 686898 64166 687134
rect 64250 686898 64486 687134
rect 64570 686898 64806 687134
rect 83930 687218 84166 687454
rect 84250 687218 84486 687454
rect 84570 687218 84806 687454
rect 83930 686898 84166 687134
rect 84250 686898 84486 687134
rect 84570 686898 84806 687134
rect 103930 687218 104166 687454
rect 104250 687218 104486 687454
rect 104570 687218 104806 687454
rect 103930 686898 104166 687134
rect 104250 686898 104486 687134
rect 104570 686898 104806 687134
rect 123930 687218 124166 687454
rect 124250 687218 124486 687454
rect 124570 687218 124806 687454
rect 123930 686898 124166 687134
rect 124250 686898 124486 687134
rect 124570 686898 124806 687134
rect 143930 687218 144166 687454
rect 144250 687218 144486 687454
rect 144570 687218 144806 687454
rect 143930 686898 144166 687134
rect 144250 686898 144486 687134
rect 144570 686898 144806 687134
rect 163930 687218 164166 687454
rect 164250 687218 164486 687454
rect 164570 687218 164806 687454
rect 163930 686898 164166 687134
rect 164250 686898 164486 687134
rect 164570 686898 164806 687134
rect 183930 687218 184166 687454
rect 184250 687218 184486 687454
rect 184570 687218 184806 687454
rect 183930 686898 184166 687134
rect 184250 686898 184486 687134
rect 184570 686898 184806 687134
rect 203930 687218 204166 687454
rect 204250 687218 204486 687454
rect 204570 687218 204806 687454
rect 203930 686898 204166 687134
rect 204250 686898 204486 687134
rect 204570 686898 204806 687134
rect 223930 687218 224166 687454
rect 224250 687218 224486 687454
rect 224570 687218 224806 687454
rect 223930 686898 224166 687134
rect 224250 686898 224486 687134
rect 224570 686898 224806 687134
rect 243930 687218 244166 687454
rect 244250 687218 244486 687454
rect 244570 687218 244806 687454
rect 243930 686898 244166 687134
rect 244250 686898 244486 687134
rect 244570 686898 244806 687134
rect 263930 687218 264166 687454
rect 264250 687218 264486 687454
rect 264570 687218 264806 687454
rect 263930 686898 264166 687134
rect 264250 686898 264486 687134
rect 264570 686898 264806 687134
rect 283930 687218 284166 687454
rect 284250 687218 284486 687454
rect 284570 687218 284806 687454
rect 283930 686898 284166 687134
rect 284250 686898 284486 687134
rect 284570 686898 284806 687134
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 33930 655718 34166 655954
rect 34250 655718 34486 655954
rect 34570 655718 34806 655954
rect 33930 655398 34166 655634
rect 34250 655398 34486 655634
rect 34570 655398 34806 655634
rect 53930 655718 54166 655954
rect 54250 655718 54486 655954
rect 54570 655718 54806 655954
rect 53930 655398 54166 655634
rect 54250 655398 54486 655634
rect 54570 655398 54806 655634
rect 73930 655718 74166 655954
rect 74250 655718 74486 655954
rect 74570 655718 74806 655954
rect 73930 655398 74166 655634
rect 74250 655398 74486 655634
rect 74570 655398 74806 655634
rect 93930 655718 94166 655954
rect 94250 655718 94486 655954
rect 94570 655718 94806 655954
rect 93930 655398 94166 655634
rect 94250 655398 94486 655634
rect 94570 655398 94806 655634
rect 113930 655718 114166 655954
rect 114250 655718 114486 655954
rect 114570 655718 114806 655954
rect 113930 655398 114166 655634
rect 114250 655398 114486 655634
rect 114570 655398 114806 655634
rect 133930 655718 134166 655954
rect 134250 655718 134486 655954
rect 134570 655718 134806 655954
rect 133930 655398 134166 655634
rect 134250 655398 134486 655634
rect 134570 655398 134806 655634
rect 153930 655718 154166 655954
rect 154250 655718 154486 655954
rect 154570 655718 154806 655954
rect 153930 655398 154166 655634
rect 154250 655398 154486 655634
rect 154570 655398 154806 655634
rect 173930 655718 174166 655954
rect 174250 655718 174486 655954
rect 174570 655718 174806 655954
rect 173930 655398 174166 655634
rect 174250 655398 174486 655634
rect 174570 655398 174806 655634
rect 193930 655718 194166 655954
rect 194250 655718 194486 655954
rect 194570 655718 194806 655954
rect 193930 655398 194166 655634
rect 194250 655398 194486 655634
rect 194570 655398 194806 655634
rect 213930 655718 214166 655954
rect 214250 655718 214486 655954
rect 214570 655718 214806 655954
rect 213930 655398 214166 655634
rect 214250 655398 214486 655634
rect 214570 655398 214806 655634
rect 233930 655718 234166 655954
rect 234250 655718 234486 655954
rect 234570 655718 234806 655954
rect 233930 655398 234166 655634
rect 234250 655398 234486 655634
rect 234570 655398 234806 655634
rect 253930 655718 254166 655954
rect 254250 655718 254486 655954
rect 254570 655718 254806 655954
rect 253930 655398 254166 655634
rect 254250 655398 254486 655634
rect 254570 655398 254806 655634
rect 273930 655718 274166 655954
rect 274250 655718 274486 655954
rect 274570 655718 274806 655954
rect 273930 655398 274166 655634
rect 274250 655398 274486 655634
rect 274570 655398 274806 655634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 23930 651218 24166 651454
rect 24250 651218 24486 651454
rect 24570 651218 24806 651454
rect 23930 650898 24166 651134
rect 24250 650898 24486 651134
rect 24570 650898 24806 651134
rect 43930 651218 44166 651454
rect 44250 651218 44486 651454
rect 44570 651218 44806 651454
rect 43930 650898 44166 651134
rect 44250 650898 44486 651134
rect 44570 650898 44806 651134
rect 63930 651218 64166 651454
rect 64250 651218 64486 651454
rect 64570 651218 64806 651454
rect 63930 650898 64166 651134
rect 64250 650898 64486 651134
rect 64570 650898 64806 651134
rect 83930 651218 84166 651454
rect 84250 651218 84486 651454
rect 84570 651218 84806 651454
rect 83930 650898 84166 651134
rect 84250 650898 84486 651134
rect 84570 650898 84806 651134
rect 103930 651218 104166 651454
rect 104250 651218 104486 651454
rect 104570 651218 104806 651454
rect 103930 650898 104166 651134
rect 104250 650898 104486 651134
rect 104570 650898 104806 651134
rect 123930 651218 124166 651454
rect 124250 651218 124486 651454
rect 124570 651218 124806 651454
rect 123930 650898 124166 651134
rect 124250 650898 124486 651134
rect 124570 650898 124806 651134
rect 143930 651218 144166 651454
rect 144250 651218 144486 651454
rect 144570 651218 144806 651454
rect 143930 650898 144166 651134
rect 144250 650898 144486 651134
rect 144570 650898 144806 651134
rect 163930 651218 164166 651454
rect 164250 651218 164486 651454
rect 164570 651218 164806 651454
rect 163930 650898 164166 651134
rect 164250 650898 164486 651134
rect 164570 650898 164806 651134
rect 183930 651218 184166 651454
rect 184250 651218 184486 651454
rect 184570 651218 184806 651454
rect 183930 650898 184166 651134
rect 184250 650898 184486 651134
rect 184570 650898 184806 651134
rect 203930 651218 204166 651454
rect 204250 651218 204486 651454
rect 204570 651218 204806 651454
rect 203930 650898 204166 651134
rect 204250 650898 204486 651134
rect 204570 650898 204806 651134
rect 223930 651218 224166 651454
rect 224250 651218 224486 651454
rect 224570 651218 224806 651454
rect 223930 650898 224166 651134
rect 224250 650898 224486 651134
rect 224570 650898 224806 651134
rect 243930 651218 244166 651454
rect 244250 651218 244486 651454
rect 244570 651218 244806 651454
rect 243930 650898 244166 651134
rect 244250 650898 244486 651134
rect 244570 650898 244806 651134
rect 263930 651218 264166 651454
rect 264250 651218 264486 651454
rect 264570 651218 264806 651454
rect 263930 650898 264166 651134
rect 264250 650898 264486 651134
rect 264570 650898 264806 651134
rect 283930 651218 284166 651454
rect 284250 651218 284486 651454
rect 284570 651218 284806 651454
rect 283930 650898 284166 651134
rect 284250 650898 284486 651134
rect 284570 650898 284806 651134
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 33930 619718 34166 619954
rect 34250 619718 34486 619954
rect 34570 619718 34806 619954
rect 33930 619398 34166 619634
rect 34250 619398 34486 619634
rect 34570 619398 34806 619634
rect 53930 619718 54166 619954
rect 54250 619718 54486 619954
rect 54570 619718 54806 619954
rect 53930 619398 54166 619634
rect 54250 619398 54486 619634
rect 54570 619398 54806 619634
rect 73930 619718 74166 619954
rect 74250 619718 74486 619954
rect 74570 619718 74806 619954
rect 73930 619398 74166 619634
rect 74250 619398 74486 619634
rect 74570 619398 74806 619634
rect 93930 619718 94166 619954
rect 94250 619718 94486 619954
rect 94570 619718 94806 619954
rect 93930 619398 94166 619634
rect 94250 619398 94486 619634
rect 94570 619398 94806 619634
rect 113930 619718 114166 619954
rect 114250 619718 114486 619954
rect 114570 619718 114806 619954
rect 113930 619398 114166 619634
rect 114250 619398 114486 619634
rect 114570 619398 114806 619634
rect 133930 619718 134166 619954
rect 134250 619718 134486 619954
rect 134570 619718 134806 619954
rect 133930 619398 134166 619634
rect 134250 619398 134486 619634
rect 134570 619398 134806 619634
rect 153930 619718 154166 619954
rect 154250 619718 154486 619954
rect 154570 619718 154806 619954
rect 153930 619398 154166 619634
rect 154250 619398 154486 619634
rect 154570 619398 154806 619634
rect 173930 619718 174166 619954
rect 174250 619718 174486 619954
rect 174570 619718 174806 619954
rect 173930 619398 174166 619634
rect 174250 619398 174486 619634
rect 174570 619398 174806 619634
rect 193930 619718 194166 619954
rect 194250 619718 194486 619954
rect 194570 619718 194806 619954
rect 193930 619398 194166 619634
rect 194250 619398 194486 619634
rect 194570 619398 194806 619634
rect 213930 619718 214166 619954
rect 214250 619718 214486 619954
rect 214570 619718 214806 619954
rect 213930 619398 214166 619634
rect 214250 619398 214486 619634
rect 214570 619398 214806 619634
rect 233930 619718 234166 619954
rect 234250 619718 234486 619954
rect 234570 619718 234806 619954
rect 233930 619398 234166 619634
rect 234250 619398 234486 619634
rect 234570 619398 234806 619634
rect 253930 619718 254166 619954
rect 254250 619718 254486 619954
rect 254570 619718 254806 619954
rect 253930 619398 254166 619634
rect 254250 619398 254486 619634
rect 254570 619398 254806 619634
rect 273930 619718 274166 619954
rect 274250 619718 274486 619954
rect 274570 619718 274806 619954
rect 273930 619398 274166 619634
rect 274250 619398 274486 619634
rect 274570 619398 274806 619634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 23930 615218 24166 615454
rect 24250 615218 24486 615454
rect 24570 615218 24806 615454
rect 23930 614898 24166 615134
rect 24250 614898 24486 615134
rect 24570 614898 24806 615134
rect 43930 615218 44166 615454
rect 44250 615218 44486 615454
rect 44570 615218 44806 615454
rect 43930 614898 44166 615134
rect 44250 614898 44486 615134
rect 44570 614898 44806 615134
rect 63930 615218 64166 615454
rect 64250 615218 64486 615454
rect 64570 615218 64806 615454
rect 63930 614898 64166 615134
rect 64250 614898 64486 615134
rect 64570 614898 64806 615134
rect 83930 615218 84166 615454
rect 84250 615218 84486 615454
rect 84570 615218 84806 615454
rect 83930 614898 84166 615134
rect 84250 614898 84486 615134
rect 84570 614898 84806 615134
rect 103930 615218 104166 615454
rect 104250 615218 104486 615454
rect 104570 615218 104806 615454
rect 103930 614898 104166 615134
rect 104250 614898 104486 615134
rect 104570 614898 104806 615134
rect 123930 615218 124166 615454
rect 124250 615218 124486 615454
rect 124570 615218 124806 615454
rect 123930 614898 124166 615134
rect 124250 614898 124486 615134
rect 124570 614898 124806 615134
rect 143930 615218 144166 615454
rect 144250 615218 144486 615454
rect 144570 615218 144806 615454
rect 143930 614898 144166 615134
rect 144250 614898 144486 615134
rect 144570 614898 144806 615134
rect 163930 615218 164166 615454
rect 164250 615218 164486 615454
rect 164570 615218 164806 615454
rect 163930 614898 164166 615134
rect 164250 614898 164486 615134
rect 164570 614898 164806 615134
rect 183930 615218 184166 615454
rect 184250 615218 184486 615454
rect 184570 615218 184806 615454
rect 183930 614898 184166 615134
rect 184250 614898 184486 615134
rect 184570 614898 184806 615134
rect 203930 615218 204166 615454
rect 204250 615218 204486 615454
rect 204570 615218 204806 615454
rect 203930 614898 204166 615134
rect 204250 614898 204486 615134
rect 204570 614898 204806 615134
rect 223930 615218 224166 615454
rect 224250 615218 224486 615454
rect 224570 615218 224806 615454
rect 223930 614898 224166 615134
rect 224250 614898 224486 615134
rect 224570 614898 224806 615134
rect 243930 615218 244166 615454
rect 244250 615218 244486 615454
rect 244570 615218 244806 615454
rect 243930 614898 244166 615134
rect 244250 614898 244486 615134
rect 244570 614898 244806 615134
rect 263930 615218 264166 615454
rect 264250 615218 264486 615454
rect 264570 615218 264806 615454
rect 263930 614898 264166 615134
rect 264250 614898 264486 615134
rect 264570 614898 264806 615134
rect 283930 615218 284166 615454
rect 284250 615218 284486 615454
rect 284570 615218 284806 615454
rect 283930 614898 284166 615134
rect 284250 614898 284486 615134
rect 284570 614898 284806 615134
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 33930 547718 34166 547954
rect 34250 547718 34486 547954
rect 34570 547718 34806 547954
rect 33930 547398 34166 547634
rect 34250 547398 34486 547634
rect 34570 547398 34806 547634
rect 53930 547718 54166 547954
rect 54250 547718 54486 547954
rect 54570 547718 54806 547954
rect 53930 547398 54166 547634
rect 54250 547398 54486 547634
rect 54570 547398 54806 547634
rect 73930 547718 74166 547954
rect 74250 547718 74486 547954
rect 74570 547718 74806 547954
rect 73930 547398 74166 547634
rect 74250 547398 74486 547634
rect 74570 547398 74806 547634
rect 93930 547718 94166 547954
rect 94250 547718 94486 547954
rect 94570 547718 94806 547954
rect 93930 547398 94166 547634
rect 94250 547398 94486 547634
rect 94570 547398 94806 547634
rect 113930 547718 114166 547954
rect 114250 547718 114486 547954
rect 114570 547718 114806 547954
rect 113930 547398 114166 547634
rect 114250 547398 114486 547634
rect 114570 547398 114806 547634
rect 133930 547718 134166 547954
rect 134250 547718 134486 547954
rect 134570 547718 134806 547954
rect 133930 547398 134166 547634
rect 134250 547398 134486 547634
rect 134570 547398 134806 547634
rect 153930 547718 154166 547954
rect 154250 547718 154486 547954
rect 154570 547718 154806 547954
rect 153930 547398 154166 547634
rect 154250 547398 154486 547634
rect 154570 547398 154806 547634
rect 173930 547718 174166 547954
rect 174250 547718 174486 547954
rect 174570 547718 174806 547954
rect 173930 547398 174166 547634
rect 174250 547398 174486 547634
rect 174570 547398 174806 547634
rect 193930 547718 194166 547954
rect 194250 547718 194486 547954
rect 194570 547718 194806 547954
rect 193930 547398 194166 547634
rect 194250 547398 194486 547634
rect 194570 547398 194806 547634
rect 213930 547718 214166 547954
rect 214250 547718 214486 547954
rect 214570 547718 214806 547954
rect 213930 547398 214166 547634
rect 214250 547398 214486 547634
rect 214570 547398 214806 547634
rect 233930 547718 234166 547954
rect 234250 547718 234486 547954
rect 234570 547718 234806 547954
rect 233930 547398 234166 547634
rect 234250 547398 234486 547634
rect 234570 547398 234806 547634
rect 253930 547718 254166 547954
rect 254250 547718 254486 547954
rect 254570 547718 254806 547954
rect 253930 547398 254166 547634
rect 254250 547398 254486 547634
rect 254570 547398 254806 547634
rect 273930 547718 274166 547954
rect 274250 547718 274486 547954
rect 274570 547718 274806 547954
rect 273930 547398 274166 547634
rect 274250 547398 274486 547634
rect 274570 547398 274806 547634
rect 23930 543218 24166 543454
rect 24250 543218 24486 543454
rect 24570 543218 24806 543454
rect 23930 542898 24166 543134
rect 24250 542898 24486 543134
rect 24570 542898 24806 543134
rect 43930 543218 44166 543454
rect 44250 543218 44486 543454
rect 44570 543218 44806 543454
rect 43930 542898 44166 543134
rect 44250 542898 44486 543134
rect 44570 542898 44806 543134
rect 63930 543218 64166 543454
rect 64250 543218 64486 543454
rect 64570 543218 64806 543454
rect 63930 542898 64166 543134
rect 64250 542898 64486 543134
rect 64570 542898 64806 543134
rect 83930 543218 84166 543454
rect 84250 543218 84486 543454
rect 84570 543218 84806 543454
rect 83930 542898 84166 543134
rect 84250 542898 84486 543134
rect 84570 542898 84806 543134
rect 103930 543218 104166 543454
rect 104250 543218 104486 543454
rect 104570 543218 104806 543454
rect 103930 542898 104166 543134
rect 104250 542898 104486 543134
rect 104570 542898 104806 543134
rect 123930 543218 124166 543454
rect 124250 543218 124486 543454
rect 124570 543218 124806 543454
rect 123930 542898 124166 543134
rect 124250 542898 124486 543134
rect 124570 542898 124806 543134
rect 143930 543218 144166 543454
rect 144250 543218 144486 543454
rect 144570 543218 144806 543454
rect 143930 542898 144166 543134
rect 144250 542898 144486 543134
rect 144570 542898 144806 543134
rect 163930 543218 164166 543454
rect 164250 543218 164486 543454
rect 164570 543218 164806 543454
rect 163930 542898 164166 543134
rect 164250 542898 164486 543134
rect 164570 542898 164806 543134
rect 183930 543218 184166 543454
rect 184250 543218 184486 543454
rect 184570 543218 184806 543454
rect 183930 542898 184166 543134
rect 184250 542898 184486 543134
rect 184570 542898 184806 543134
rect 203930 543218 204166 543454
rect 204250 543218 204486 543454
rect 204570 543218 204806 543454
rect 203930 542898 204166 543134
rect 204250 542898 204486 543134
rect 204570 542898 204806 543134
rect 223930 543218 224166 543454
rect 224250 543218 224486 543454
rect 224570 543218 224806 543454
rect 223930 542898 224166 543134
rect 224250 542898 224486 543134
rect 224570 542898 224806 543134
rect 243930 543218 244166 543454
rect 244250 543218 244486 543454
rect 244570 543218 244806 543454
rect 243930 542898 244166 543134
rect 244250 542898 244486 543134
rect 244570 542898 244806 543134
rect 263930 543218 264166 543454
rect 264250 543218 264486 543454
rect 264570 543218 264806 543454
rect 263930 542898 264166 543134
rect 264250 542898 264486 543134
rect 264570 542898 264806 543134
rect 283930 543218 284166 543454
rect 284250 543218 284486 543454
rect 284570 543218 284806 543454
rect 283930 542898 284166 543134
rect 284250 542898 284486 543134
rect 284570 542898 284806 543134
rect 33930 511718 34166 511954
rect 34250 511718 34486 511954
rect 34570 511718 34806 511954
rect 33930 511398 34166 511634
rect 34250 511398 34486 511634
rect 34570 511398 34806 511634
rect 53930 511718 54166 511954
rect 54250 511718 54486 511954
rect 54570 511718 54806 511954
rect 53930 511398 54166 511634
rect 54250 511398 54486 511634
rect 54570 511398 54806 511634
rect 73930 511718 74166 511954
rect 74250 511718 74486 511954
rect 74570 511718 74806 511954
rect 73930 511398 74166 511634
rect 74250 511398 74486 511634
rect 74570 511398 74806 511634
rect 93930 511718 94166 511954
rect 94250 511718 94486 511954
rect 94570 511718 94806 511954
rect 93930 511398 94166 511634
rect 94250 511398 94486 511634
rect 94570 511398 94806 511634
rect 113930 511718 114166 511954
rect 114250 511718 114486 511954
rect 114570 511718 114806 511954
rect 113930 511398 114166 511634
rect 114250 511398 114486 511634
rect 114570 511398 114806 511634
rect 133930 511718 134166 511954
rect 134250 511718 134486 511954
rect 134570 511718 134806 511954
rect 133930 511398 134166 511634
rect 134250 511398 134486 511634
rect 134570 511398 134806 511634
rect 153930 511718 154166 511954
rect 154250 511718 154486 511954
rect 154570 511718 154806 511954
rect 153930 511398 154166 511634
rect 154250 511398 154486 511634
rect 154570 511398 154806 511634
rect 173930 511718 174166 511954
rect 174250 511718 174486 511954
rect 174570 511718 174806 511954
rect 173930 511398 174166 511634
rect 174250 511398 174486 511634
rect 174570 511398 174806 511634
rect 193930 511718 194166 511954
rect 194250 511718 194486 511954
rect 194570 511718 194806 511954
rect 193930 511398 194166 511634
rect 194250 511398 194486 511634
rect 194570 511398 194806 511634
rect 213930 511718 214166 511954
rect 214250 511718 214486 511954
rect 214570 511718 214806 511954
rect 213930 511398 214166 511634
rect 214250 511398 214486 511634
rect 214570 511398 214806 511634
rect 233930 511718 234166 511954
rect 234250 511718 234486 511954
rect 234570 511718 234806 511954
rect 233930 511398 234166 511634
rect 234250 511398 234486 511634
rect 234570 511398 234806 511634
rect 253930 511718 254166 511954
rect 254250 511718 254486 511954
rect 254570 511718 254806 511954
rect 253930 511398 254166 511634
rect 254250 511398 254486 511634
rect 254570 511398 254806 511634
rect 273930 511718 274166 511954
rect 274250 511718 274486 511954
rect 274570 511718 274806 511954
rect 273930 511398 274166 511634
rect 274250 511398 274486 511634
rect 274570 511398 274806 511634
rect 23930 507218 24166 507454
rect 24250 507218 24486 507454
rect 24570 507218 24806 507454
rect 23930 506898 24166 507134
rect 24250 506898 24486 507134
rect 24570 506898 24806 507134
rect 43930 507218 44166 507454
rect 44250 507218 44486 507454
rect 44570 507218 44806 507454
rect 43930 506898 44166 507134
rect 44250 506898 44486 507134
rect 44570 506898 44806 507134
rect 63930 507218 64166 507454
rect 64250 507218 64486 507454
rect 64570 507218 64806 507454
rect 63930 506898 64166 507134
rect 64250 506898 64486 507134
rect 64570 506898 64806 507134
rect 83930 507218 84166 507454
rect 84250 507218 84486 507454
rect 84570 507218 84806 507454
rect 83930 506898 84166 507134
rect 84250 506898 84486 507134
rect 84570 506898 84806 507134
rect 103930 507218 104166 507454
rect 104250 507218 104486 507454
rect 104570 507218 104806 507454
rect 103930 506898 104166 507134
rect 104250 506898 104486 507134
rect 104570 506898 104806 507134
rect 123930 507218 124166 507454
rect 124250 507218 124486 507454
rect 124570 507218 124806 507454
rect 123930 506898 124166 507134
rect 124250 506898 124486 507134
rect 124570 506898 124806 507134
rect 143930 507218 144166 507454
rect 144250 507218 144486 507454
rect 144570 507218 144806 507454
rect 143930 506898 144166 507134
rect 144250 506898 144486 507134
rect 144570 506898 144806 507134
rect 163930 507218 164166 507454
rect 164250 507218 164486 507454
rect 164570 507218 164806 507454
rect 163930 506898 164166 507134
rect 164250 506898 164486 507134
rect 164570 506898 164806 507134
rect 183930 507218 184166 507454
rect 184250 507218 184486 507454
rect 184570 507218 184806 507454
rect 183930 506898 184166 507134
rect 184250 506898 184486 507134
rect 184570 506898 184806 507134
rect 203930 507218 204166 507454
rect 204250 507218 204486 507454
rect 204570 507218 204806 507454
rect 203930 506898 204166 507134
rect 204250 506898 204486 507134
rect 204570 506898 204806 507134
rect 223930 507218 224166 507454
rect 224250 507218 224486 507454
rect 224570 507218 224806 507454
rect 223930 506898 224166 507134
rect 224250 506898 224486 507134
rect 224570 506898 224806 507134
rect 243930 507218 244166 507454
rect 244250 507218 244486 507454
rect 244570 507218 244806 507454
rect 243930 506898 244166 507134
rect 244250 506898 244486 507134
rect 244570 506898 244806 507134
rect 263930 507218 264166 507454
rect 264250 507218 264486 507454
rect 264570 507218 264806 507454
rect 263930 506898 264166 507134
rect 264250 506898 264486 507134
rect 264570 506898 264806 507134
rect 283930 507218 284166 507454
rect 284250 507218 284486 507454
rect 284570 507218 284806 507454
rect 283930 506898 284166 507134
rect 284250 506898 284486 507134
rect 284570 506898 284806 507134
rect 33930 475718 34166 475954
rect 34250 475718 34486 475954
rect 34570 475718 34806 475954
rect 33930 475398 34166 475634
rect 34250 475398 34486 475634
rect 34570 475398 34806 475634
rect 53930 475718 54166 475954
rect 54250 475718 54486 475954
rect 54570 475718 54806 475954
rect 53930 475398 54166 475634
rect 54250 475398 54486 475634
rect 54570 475398 54806 475634
rect 73930 475718 74166 475954
rect 74250 475718 74486 475954
rect 74570 475718 74806 475954
rect 73930 475398 74166 475634
rect 74250 475398 74486 475634
rect 74570 475398 74806 475634
rect 93930 475718 94166 475954
rect 94250 475718 94486 475954
rect 94570 475718 94806 475954
rect 93930 475398 94166 475634
rect 94250 475398 94486 475634
rect 94570 475398 94806 475634
rect 113930 475718 114166 475954
rect 114250 475718 114486 475954
rect 114570 475718 114806 475954
rect 113930 475398 114166 475634
rect 114250 475398 114486 475634
rect 114570 475398 114806 475634
rect 133930 475718 134166 475954
rect 134250 475718 134486 475954
rect 134570 475718 134806 475954
rect 133930 475398 134166 475634
rect 134250 475398 134486 475634
rect 134570 475398 134806 475634
rect 153930 475718 154166 475954
rect 154250 475718 154486 475954
rect 154570 475718 154806 475954
rect 153930 475398 154166 475634
rect 154250 475398 154486 475634
rect 154570 475398 154806 475634
rect 173930 475718 174166 475954
rect 174250 475718 174486 475954
rect 174570 475718 174806 475954
rect 173930 475398 174166 475634
rect 174250 475398 174486 475634
rect 174570 475398 174806 475634
rect 193930 475718 194166 475954
rect 194250 475718 194486 475954
rect 194570 475718 194806 475954
rect 193930 475398 194166 475634
rect 194250 475398 194486 475634
rect 194570 475398 194806 475634
rect 213930 475718 214166 475954
rect 214250 475718 214486 475954
rect 214570 475718 214806 475954
rect 213930 475398 214166 475634
rect 214250 475398 214486 475634
rect 214570 475398 214806 475634
rect 233930 475718 234166 475954
rect 234250 475718 234486 475954
rect 234570 475718 234806 475954
rect 233930 475398 234166 475634
rect 234250 475398 234486 475634
rect 234570 475398 234806 475634
rect 253930 475718 254166 475954
rect 254250 475718 254486 475954
rect 254570 475718 254806 475954
rect 253930 475398 254166 475634
rect 254250 475398 254486 475634
rect 254570 475398 254806 475634
rect 273930 475718 274166 475954
rect 274250 475718 274486 475954
rect 274570 475718 274806 475954
rect 273930 475398 274166 475634
rect 274250 475398 274486 475634
rect 274570 475398 274806 475634
rect 23930 471218 24166 471454
rect 24250 471218 24486 471454
rect 24570 471218 24806 471454
rect 23930 470898 24166 471134
rect 24250 470898 24486 471134
rect 24570 470898 24806 471134
rect 43930 471218 44166 471454
rect 44250 471218 44486 471454
rect 44570 471218 44806 471454
rect 43930 470898 44166 471134
rect 44250 470898 44486 471134
rect 44570 470898 44806 471134
rect 63930 471218 64166 471454
rect 64250 471218 64486 471454
rect 64570 471218 64806 471454
rect 63930 470898 64166 471134
rect 64250 470898 64486 471134
rect 64570 470898 64806 471134
rect 83930 471218 84166 471454
rect 84250 471218 84486 471454
rect 84570 471218 84806 471454
rect 83930 470898 84166 471134
rect 84250 470898 84486 471134
rect 84570 470898 84806 471134
rect 103930 471218 104166 471454
rect 104250 471218 104486 471454
rect 104570 471218 104806 471454
rect 103930 470898 104166 471134
rect 104250 470898 104486 471134
rect 104570 470898 104806 471134
rect 123930 471218 124166 471454
rect 124250 471218 124486 471454
rect 124570 471218 124806 471454
rect 123930 470898 124166 471134
rect 124250 470898 124486 471134
rect 124570 470898 124806 471134
rect 143930 471218 144166 471454
rect 144250 471218 144486 471454
rect 144570 471218 144806 471454
rect 143930 470898 144166 471134
rect 144250 470898 144486 471134
rect 144570 470898 144806 471134
rect 163930 471218 164166 471454
rect 164250 471218 164486 471454
rect 164570 471218 164806 471454
rect 163930 470898 164166 471134
rect 164250 470898 164486 471134
rect 164570 470898 164806 471134
rect 183930 471218 184166 471454
rect 184250 471218 184486 471454
rect 184570 471218 184806 471454
rect 183930 470898 184166 471134
rect 184250 470898 184486 471134
rect 184570 470898 184806 471134
rect 203930 471218 204166 471454
rect 204250 471218 204486 471454
rect 204570 471218 204806 471454
rect 203930 470898 204166 471134
rect 204250 470898 204486 471134
rect 204570 470898 204806 471134
rect 223930 471218 224166 471454
rect 224250 471218 224486 471454
rect 224570 471218 224806 471454
rect 223930 470898 224166 471134
rect 224250 470898 224486 471134
rect 224570 470898 224806 471134
rect 243930 471218 244166 471454
rect 244250 471218 244486 471454
rect 244570 471218 244806 471454
rect 243930 470898 244166 471134
rect 244250 470898 244486 471134
rect 244570 470898 244806 471134
rect 263930 471218 264166 471454
rect 264250 471218 264486 471454
rect 264570 471218 264806 471454
rect 263930 470898 264166 471134
rect 264250 470898 264486 471134
rect 264570 470898 264806 471134
rect 283930 471218 284166 471454
rect 284250 471218 284486 471454
rect 284570 471218 284806 471454
rect 283930 470898 284166 471134
rect 284250 470898 284486 471134
rect 284570 470898 284806 471134
rect 33930 439718 34166 439954
rect 34250 439718 34486 439954
rect 34570 439718 34806 439954
rect 33930 439398 34166 439634
rect 34250 439398 34486 439634
rect 34570 439398 34806 439634
rect 53930 439718 54166 439954
rect 54250 439718 54486 439954
rect 54570 439718 54806 439954
rect 53930 439398 54166 439634
rect 54250 439398 54486 439634
rect 54570 439398 54806 439634
rect 73930 439718 74166 439954
rect 74250 439718 74486 439954
rect 74570 439718 74806 439954
rect 73930 439398 74166 439634
rect 74250 439398 74486 439634
rect 74570 439398 74806 439634
rect 93930 439718 94166 439954
rect 94250 439718 94486 439954
rect 94570 439718 94806 439954
rect 93930 439398 94166 439634
rect 94250 439398 94486 439634
rect 94570 439398 94806 439634
rect 113930 439718 114166 439954
rect 114250 439718 114486 439954
rect 114570 439718 114806 439954
rect 113930 439398 114166 439634
rect 114250 439398 114486 439634
rect 114570 439398 114806 439634
rect 133930 439718 134166 439954
rect 134250 439718 134486 439954
rect 134570 439718 134806 439954
rect 133930 439398 134166 439634
rect 134250 439398 134486 439634
rect 134570 439398 134806 439634
rect 153930 439718 154166 439954
rect 154250 439718 154486 439954
rect 154570 439718 154806 439954
rect 153930 439398 154166 439634
rect 154250 439398 154486 439634
rect 154570 439398 154806 439634
rect 173930 439718 174166 439954
rect 174250 439718 174486 439954
rect 174570 439718 174806 439954
rect 173930 439398 174166 439634
rect 174250 439398 174486 439634
rect 174570 439398 174806 439634
rect 193930 439718 194166 439954
rect 194250 439718 194486 439954
rect 194570 439718 194806 439954
rect 193930 439398 194166 439634
rect 194250 439398 194486 439634
rect 194570 439398 194806 439634
rect 213930 439718 214166 439954
rect 214250 439718 214486 439954
rect 214570 439718 214806 439954
rect 213930 439398 214166 439634
rect 214250 439398 214486 439634
rect 214570 439398 214806 439634
rect 233930 439718 234166 439954
rect 234250 439718 234486 439954
rect 234570 439718 234806 439954
rect 233930 439398 234166 439634
rect 234250 439398 234486 439634
rect 234570 439398 234806 439634
rect 253930 439718 254166 439954
rect 254250 439718 254486 439954
rect 254570 439718 254806 439954
rect 253930 439398 254166 439634
rect 254250 439398 254486 439634
rect 254570 439398 254806 439634
rect 273930 439718 274166 439954
rect 274250 439718 274486 439954
rect 274570 439718 274806 439954
rect 273930 439398 274166 439634
rect 274250 439398 274486 439634
rect 274570 439398 274806 439634
rect 23930 435218 24166 435454
rect 24250 435218 24486 435454
rect 24570 435218 24806 435454
rect 23930 434898 24166 435134
rect 24250 434898 24486 435134
rect 24570 434898 24806 435134
rect 43930 435218 44166 435454
rect 44250 435218 44486 435454
rect 44570 435218 44806 435454
rect 43930 434898 44166 435134
rect 44250 434898 44486 435134
rect 44570 434898 44806 435134
rect 63930 435218 64166 435454
rect 64250 435218 64486 435454
rect 64570 435218 64806 435454
rect 63930 434898 64166 435134
rect 64250 434898 64486 435134
rect 64570 434898 64806 435134
rect 83930 435218 84166 435454
rect 84250 435218 84486 435454
rect 84570 435218 84806 435454
rect 83930 434898 84166 435134
rect 84250 434898 84486 435134
rect 84570 434898 84806 435134
rect 103930 435218 104166 435454
rect 104250 435218 104486 435454
rect 104570 435218 104806 435454
rect 103930 434898 104166 435134
rect 104250 434898 104486 435134
rect 104570 434898 104806 435134
rect 123930 435218 124166 435454
rect 124250 435218 124486 435454
rect 124570 435218 124806 435454
rect 123930 434898 124166 435134
rect 124250 434898 124486 435134
rect 124570 434898 124806 435134
rect 143930 435218 144166 435454
rect 144250 435218 144486 435454
rect 144570 435218 144806 435454
rect 143930 434898 144166 435134
rect 144250 434898 144486 435134
rect 144570 434898 144806 435134
rect 163930 435218 164166 435454
rect 164250 435218 164486 435454
rect 164570 435218 164806 435454
rect 163930 434898 164166 435134
rect 164250 434898 164486 435134
rect 164570 434898 164806 435134
rect 183930 435218 184166 435454
rect 184250 435218 184486 435454
rect 184570 435218 184806 435454
rect 183930 434898 184166 435134
rect 184250 434898 184486 435134
rect 184570 434898 184806 435134
rect 203930 435218 204166 435454
rect 204250 435218 204486 435454
rect 204570 435218 204806 435454
rect 203930 434898 204166 435134
rect 204250 434898 204486 435134
rect 204570 434898 204806 435134
rect 223930 435218 224166 435454
rect 224250 435218 224486 435454
rect 224570 435218 224806 435454
rect 223930 434898 224166 435134
rect 224250 434898 224486 435134
rect 224570 434898 224806 435134
rect 243930 435218 244166 435454
rect 244250 435218 244486 435454
rect 244570 435218 244806 435454
rect 243930 434898 244166 435134
rect 244250 434898 244486 435134
rect 244570 434898 244806 435134
rect 263930 435218 264166 435454
rect 264250 435218 264486 435454
rect 264570 435218 264806 435454
rect 263930 434898 264166 435134
rect 264250 434898 264486 435134
rect 264570 434898 264806 435134
rect 283930 435218 284166 435454
rect 284250 435218 284486 435454
rect 284570 435218 284806 435454
rect 283930 434898 284166 435134
rect 284250 434898 284486 435134
rect 284570 434898 284806 435134
rect 33930 403718 34166 403954
rect 34250 403718 34486 403954
rect 34570 403718 34806 403954
rect 33930 403398 34166 403634
rect 34250 403398 34486 403634
rect 34570 403398 34806 403634
rect 53930 403718 54166 403954
rect 54250 403718 54486 403954
rect 54570 403718 54806 403954
rect 53930 403398 54166 403634
rect 54250 403398 54486 403634
rect 54570 403398 54806 403634
rect 73930 403718 74166 403954
rect 74250 403718 74486 403954
rect 74570 403718 74806 403954
rect 73930 403398 74166 403634
rect 74250 403398 74486 403634
rect 74570 403398 74806 403634
rect 93930 403718 94166 403954
rect 94250 403718 94486 403954
rect 94570 403718 94806 403954
rect 93930 403398 94166 403634
rect 94250 403398 94486 403634
rect 94570 403398 94806 403634
rect 113930 403718 114166 403954
rect 114250 403718 114486 403954
rect 114570 403718 114806 403954
rect 113930 403398 114166 403634
rect 114250 403398 114486 403634
rect 114570 403398 114806 403634
rect 133930 403718 134166 403954
rect 134250 403718 134486 403954
rect 134570 403718 134806 403954
rect 133930 403398 134166 403634
rect 134250 403398 134486 403634
rect 134570 403398 134806 403634
rect 153930 403718 154166 403954
rect 154250 403718 154486 403954
rect 154570 403718 154806 403954
rect 153930 403398 154166 403634
rect 154250 403398 154486 403634
rect 154570 403398 154806 403634
rect 173930 403718 174166 403954
rect 174250 403718 174486 403954
rect 174570 403718 174806 403954
rect 173930 403398 174166 403634
rect 174250 403398 174486 403634
rect 174570 403398 174806 403634
rect 193930 403718 194166 403954
rect 194250 403718 194486 403954
rect 194570 403718 194806 403954
rect 193930 403398 194166 403634
rect 194250 403398 194486 403634
rect 194570 403398 194806 403634
rect 213930 403718 214166 403954
rect 214250 403718 214486 403954
rect 214570 403718 214806 403954
rect 213930 403398 214166 403634
rect 214250 403398 214486 403634
rect 214570 403398 214806 403634
rect 233930 403718 234166 403954
rect 234250 403718 234486 403954
rect 234570 403718 234806 403954
rect 233930 403398 234166 403634
rect 234250 403398 234486 403634
rect 234570 403398 234806 403634
rect 253930 403718 254166 403954
rect 254250 403718 254486 403954
rect 254570 403718 254806 403954
rect 253930 403398 254166 403634
rect 254250 403398 254486 403634
rect 254570 403398 254806 403634
rect 273930 403718 274166 403954
rect 274250 403718 274486 403954
rect 274570 403718 274806 403954
rect 273930 403398 274166 403634
rect 274250 403398 274486 403634
rect 274570 403398 274806 403634
rect 23930 399218 24166 399454
rect 24250 399218 24486 399454
rect 24570 399218 24806 399454
rect 23930 398898 24166 399134
rect 24250 398898 24486 399134
rect 24570 398898 24806 399134
rect 43930 399218 44166 399454
rect 44250 399218 44486 399454
rect 44570 399218 44806 399454
rect 43930 398898 44166 399134
rect 44250 398898 44486 399134
rect 44570 398898 44806 399134
rect 63930 399218 64166 399454
rect 64250 399218 64486 399454
rect 64570 399218 64806 399454
rect 63930 398898 64166 399134
rect 64250 398898 64486 399134
rect 64570 398898 64806 399134
rect 83930 399218 84166 399454
rect 84250 399218 84486 399454
rect 84570 399218 84806 399454
rect 83930 398898 84166 399134
rect 84250 398898 84486 399134
rect 84570 398898 84806 399134
rect 103930 399218 104166 399454
rect 104250 399218 104486 399454
rect 104570 399218 104806 399454
rect 103930 398898 104166 399134
rect 104250 398898 104486 399134
rect 104570 398898 104806 399134
rect 123930 399218 124166 399454
rect 124250 399218 124486 399454
rect 124570 399218 124806 399454
rect 123930 398898 124166 399134
rect 124250 398898 124486 399134
rect 124570 398898 124806 399134
rect 143930 399218 144166 399454
rect 144250 399218 144486 399454
rect 144570 399218 144806 399454
rect 143930 398898 144166 399134
rect 144250 398898 144486 399134
rect 144570 398898 144806 399134
rect 163930 399218 164166 399454
rect 164250 399218 164486 399454
rect 164570 399218 164806 399454
rect 163930 398898 164166 399134
rect 164250 398898 164486 399134
rect 164570 398898 164806 399134
rect 183930 399218 184166 399454
rect 184250 399218 184486 399454
rect 184570 399218 184806 399454
rect 183930 398898 184166 399134
rect 184250 398898 184486 399134
rect 184570 398898 184806 399134
rect 203930 399218 204166 399454
rect 204250 399218 204486 399454
rect 204570 399218 204806 399454
rect 203930 398898 204166 399134
rect 204250 398898 204486 399134
rect 204570 398898 204806 399134
rect 223930 399218 224166 399454
rect 224250 399218 224486 399454
rect 224570 399218 224806 399454
rect 223930 398898 224166 399134
rect 224250 398898 224486 399134
rect 224570 398898 224806 399134
rect 243930 399218 244166 399454
rect 244250 399218 244486 399454
rect 244570 399218 244806 399454
rect 243930 398898 244166 399134
rect 244250 398898 244486 399134
rect 244570 398898 244806 399134
rect 263930 399218 264166 399454
rect 264250 399218 264486 399454
rect 264570 399218 264806 399454
rect 263930 398898 264166 399134
rect 264250 398898 264486 399134
rect 264570 398898 264806 399134
rect 283930 399218 284166 399454
rect 284250 399218 284486 399454
rect 284570 399218 284806 399454
rect 283930 398898 284166 399134
rect 284250 398898 284486 399134
rect 284570 398898 284806 399134
rect 33930 367718 34166 367954
rect 34250 367718 34486 367954
rect 34570 367718 34806 367954
rect 33930 367398 34166 367634
rect 34250 367398 34486 367634
rect 34570 367398 34806 367634
rect 53930 367718 54166 367954
rect 54250 367718 54486 367954
rect 54570 367718 54806 367954
rect 53930 367398 54166 367634
rect 54250 367398 54486 367634
rect 54570 367398 54806 367634
rect 73930 367718 74166 367954
rect 74250 367718 74486 367954
rect 74570 367718 74806 367954
rect 73930 367398 74166 367634
rect 74250 367398 74486 367634
rect 74570 367398 74806 367634
rect 93930 367718 94166 367954
rect 94250 367718 94486 367954
rect 94570 367718 94806 367954
rect 93930 367398 94166 367634
rect 94250 367398 94486 367634
rect 94570 367398 94806 367634
rect 113930 367718 114166 367954
rect 114250 367718 114486 367954
rect 114570 367718 114806 367954
rect 113930 367398 114166 367634
rect 114250 367398 114486 367634
rect 114570 367398 114806 367634
rect 133930 367718 134166 367954
rect 134250 367718 134486 367954
rect 134570 367718 134806 367954
rect 133930 367398 134166 367634
rect 134250 367398 134486 367634
rect 134570 367398 134806 367634
rect 153930 367718 154166 367954
rect 154250 367718 154486 367954
rect 154570 367718 154806 367954
rect 153930 367398 154166 367634
rect 154250 367398 154486 367634
rect 154570 367398 154806 367634
rect 173930 367718 174166 367954
rect 174250 367718 174486 367954
rect 174570 367718 174806 367954
rect 173930 367398 174166 367634
rect 174250 367398 174486 367634
rect 174570 367398 174806 367634
rect 193930 367718 194166 367954
rect 194250 367718 194486 367954
rect 194570 367718 194806 367954
rect 193930 367398 194166 367634
rect 194250 367398 194486 367634
rect 194570 367398 194806 367634
rect 213930 367718 214166 367954
rect 214250 367718 214486 367954
rect 214570 367718 214806 367954
rect 213930 367398 214166 367634
rect 214250 367398 214486 367634
rect 214570 367398 214806 367634
rect 233930 367718 234166 367954
rect 234250 367718 234486 367954
rect 234570 367718 234806 367954
rect 233930 367398 234166 367634
rect 234250 367398 234486 367634
rect 234570 367398 234806 367634
rect 253930 367718 254166 367954
rect 254250 367718 254486 367954
rect 254570 367718 254806 367954
rect 253930 367398 254166 367634
rect 254250 367398 254486 367634
rect 254570 367398 254806 367634
rect 273930 367718 274166 367954
rect 274250 367718 274486 367954
rect 274570 367718 274806 367954
rect 273930 367398 274166 367634
rect 274250 367398 274486 367634
rect 274570 367398 274806 367634
rect 23930 363218 24166 363454
rect 24250 363218 24486 363454
rect 24570 363218 24806 363454
rect 23930 362898 24166 363134
rect 24250 362898 24486 363134
rect 24570 362898 24806 363134
rect 43930 363218 44166 363454
rect 44250 363218 44486 363454
rect 44570 363218 44806 363454
rect 43930 362898 44166 363134
rect 44250 362898 44486 363134
rect 44570 362898 44806 363134
rect 63930 363218 64166 363454
rect 64250 363218 64486 363454
rect 64570 363218 64806 363454
rect 63930 362898 64166 363134
rect 64250 362898 64486 363134
rect 64570 362898 64806 363134
rect 83930 363218 84166 363454
rect 84250 363218 84486 363454
rect 84570 363218 84806 363454
rect 83930 362898 84166 363134
rect 84250 362898 84486 363134
rect 84570 362898 84806 363134
rect 103930 363218 104166 363454
rect 104250 363218 104486 363454
rect 104570 363218 104806 363454
rect 103930 362898 104166 363134
rect 104250 362898 104486 363134
rect 104570 362898 104806 363134
rect 123930 363218 124166 363454
rect 124250 363218 124486 363454
rect 124570 363218 124806 363454
rect 123930 362898 124166 363134
rect 124250 362898 124486 363134
rect 124570 362898 124806 363134
rect 143930 363218 144166 363454
rect 144250 363218 144486 363454
rect 144570 363218 144806 363454
rect 143930 362898 144166 363134
rect 144250 362898 144486 363134
rect 144570 362898 144806 363134
rect 163930 363218 164166 363454
rect 164250 363218 164486 363454
rect 164570 363218 164806 363454
rect 163930 362898 164166 363134
rect 164250 362898 164486 363134
rect 164570 362898 164806 363134
rect 183930 363218 184166 363454
rect 184250 363218 184486 363454
rect 184570 363218 184806 363454
rect 183930 362898 184166 363134
rect 184250 362898 184486 363134
rect 184570 362898 184806 363134
rect 203930 363218 204166 363454
rect 204250 363218 204486 363454
rect 204570 363218 204806 363454
rect 203930 362898 204166 363134
rect 204250 362898 204486 363134
rect 204570 362898 204806 363134
rect 223930 363218 224166 363454
rect 224250 363218 224486 363454
rect 224570 363218 224806 363454
rect 223930 362898 224166 363134
rect 224250 362898 224486 363134
rect 224570 362898 224806 363134
rect 243930 363218 244166 363454
rect 244250 363218 244486 363454
rect 244570 363218 244806 363454
rect 243930 362898 244166 363134
rect 244250 362898 244486 363134
rect 244570 362898 244806 363134
rect 263930 363218 264166 363454
rect 264250 363218 264486 363454
rect 264570 363218 264806 363454
rect 263930 362898 264166 363134
rect 264250 362898 264486 363134
rect 264570 362898 264806 363134
rect 283930 363218 284166 363454
rect 284250 363218 284486 363454
rect 284570 363218 284806 363454
rect 283930 362898 284166 363134
rect 284250 362898 284486 363134
rect 284570 362898 284806 363134
rect 33930 295718 34166 295954
rect 34250 295718 34486 295954
rect 34570 295718 34806 295954
rect 33930 295398 34166 295634
rect 34250 295398 34486 295634
rect 34570 295398 34806 295634
rect 53930 295718 54166 295954
rect 54250 295718 54486 295954
rect 54570 295718 54806 295954
rect 53930 295398 54166 295634
rect 54250 295398 54486 295634
rect 54570 295398 54806 295634
rect 73930 295718 74166 295954
rect 74250 295718 74486 295954
rect 74570 295718 74806 295954
rect 73930 295398 74166 295634
rect 74250 295398 74486 295634
rect 74570 295398 74806 295634
rect 93930 295718 94166 295954
rect 94250 295718 94486 295954
rect 94570 295718 94806 295954
rect 93930 295398 94166 295634
rect 94250 295398 94486 295634
rect 94570 295398 94806 295634
rect 113930 295718 114166 295954
rect 114250 295718 114486 295954
rect 114570 295718 114806 295954
rect 113930 295398 114166 295634
rect 114250 295398 114486 295634
rect 114570 295398 114806 295634
rect 133930 295718 134166 295954
rect 134250 295718 134486 295954
rect 134570 295718 134806 295954
rect 133930 295398 134166 295634
rect 134250 295398 134486 295634
rect 134570 295398 134806 295634
rect 153930 295718 154166 295954
rect 154250 295718 154486 295954
rect 154570 295718 154806 295954
rect 153930 295398 154166 295634
rect 154250 295398 154486 295634
rect 154570 295398 154806 295634
rect 173930 295718 174166 295954
rect 174250 295718 174486 295954
rect 174570 295718 174806 295954
rect 173930 295398 174166 295634
rect 174250 295398 174486 295634
rect 174570 295398 174806 295634
rect 193930 295718 194166 295954
rect 194250 295718 194486 295954
rect 194570 295718 194806 295954
rect 193930 295398 194166 295634
rect 194250 295398 194486 295634
rect 194570 295398 194806 295634
rect 213930 295718 214166 295954
rect 214250 295718 214486 295954
rect 214570 295718 214806 295954
rect 213930 295398 214166 295634
rect 214250 295398 214486 295634
rect 214570 295398 214806 295634
rect 233930 295718 234166 295954
rect 234250 295718 234486 295954
rect 234570 295718 234806 295954
rect 233930 295398 234166 295634
rect 234250 295398 234486 295634
rect 234570 295398 234806 295634
rect 253930 295718 254166 295954
rect 254250 295718 254486 295954
rect 254570 295718 254806 295954
rect 253930 295398 254166 295634
rect 254250 295398 254486 295634
rect 254570 295398 254806 295634
rect 273930 295718 274166 295954
rect 274250 295718 274486 295954
rect 274570 295718 274806 295954
rect 273930 295398 274166 295634
rect 274250 295398 274486 295634
rect 274570 295398 274806 295634
rect 23930 291218 24166 291454
rect 24250 291218 24486 291454
rect 24570 291218 24806 291454
rect 23930 290898 24166 291134
rect 24250 290898 24486 291134
rect 24570 290898 24806 291134
rect 43930 291218 44166 291454
rect 44250 291218 44486 291454
rect 44570 291218 44806 291454
rect 43930 290898 44166 291134
rect 44250 290898 44486 291134
rect 44570 290898 44806 291134
rect 63930 291218 64166 291454
rect 64250 291218 64486 291454
rect 64570 291218 64806 291454
rect 63930 290898 64166 291134
rect 64250 290898 64486 291134
rect 64570 290898 64806 291134
rect 83930 291218 84166 291454
rect 84250 291218 84486 291454
rect 84570 291218 84806 291454
rect 83930 290898 84166 291134
rect 84250 290898 84486 291134
rect 84570 290898 84806 291134
rect 103930 291218 104166 291454
rect 104250 291218 104486 291454
rect 104570 291218 104806 291454
rect 103930 290898 104166 291134
rect 104250 290898 104486 291134
rect 104570 290898 104806 291134
rect 123930 291218 124166 291454
rect 124250 291218 124486 291454
rect 124570 291218 124806 291454
rect 123930 290898 124166 291134
rect 124250 290898 124486 291134
rect 124570 290898 124806 291134
rect 143930 291218 144166 291454
rect 144250 291218 144486 291454
rect 144570 291218 144806 291454
rect 143930 290898 144166 291134
rect 144250 290898 144486 291134
rect 144570 290898 144806 291134
rect 163930 291218 164166 291454
rect 164250 291218 164486 291454
rect 164570 291218 164806 291454
rect 163930 290898 164166 291134
rect 164250 290898 164486 291134
rect 164570 290898 164806 291134
rect 183930 291218 184166 291454
rect 184250 291218 184486 291454
rect 184570 291218 184806 291454
rect 183930 290898 184166 291134
rect 184250 290898 184486 291134
rect 184570 290898 184806 291134
rect 203930 291218 204166 291454
rect 204250 291218 204486 291454
rect 204570 291218 204806 291454
rect 203930 290898 204166 291134
rect 204250 290898 204486 291134
rect 204570 290898 204806 291134
rect 223930 291218 224166 291454
rect 224250 291218 224486 291454
rect 224570 291218 224806 291454
rect 223930 290898 224166 291134
rect 224250 290898 224486 291134
rect 224570 290898 224806 291134
rect 243930 291218 244166 291454
rect 244250 291218 244486 291454
rect 244570 291218 244806 291454
rect 243930 290898 244166 291134
rect 244250 290898 244486 291134
rect 244570 290898 244806 291134
rect 263930 291218 264166 291454
rect 264250 291218 264486 291454
rect 264570 291218 264806 291454
rect 263930 290898 264166 291134
rect 264250 290898 264486 291134
rect 264570 290898 264806 291134
rect 283930 291218 284166 291454
rect 284250 291218 284486 291454
rect 284570 291218 284806 291454
rect 283930 290898 284166 291134
rect 284250 290898 284486 291134
rect 284570 290898 284806 291134
rect 33930 259718 34166 259954
rect 34250 259718 34486 259954
rect 34570 259718 34806 259954
rect 33930 259398 34166 259634
rect 34250 259398 34486 259634
rect 34570 259398 34806 259634
rect 53930 259718 54166 259954
rect 54250 259718 54486 259954
rect 54570 259718 54806 259954
rect 53930 259398 54166 259634
rect 54250 259398 54486 259634
rect 54570 259398 54806 259634
rect 73930 259718 74166 259954
rect 74250 259718 74486 259954
rect 74570 259718 74806 259954
rect 73930 259398 74166 259634
rect 74250 259398 74486 259634
rect 74570 259398 74806 259634
rect 93930 259718 94166 259954
rect 94250 259718 94486 259954
rect 94570 259718 94806 259954
rect 93930 259398 94166 259634
rect 94250 259398 94486 259634
rect 94570 259398 94806 259634
rect 113930 259718 114166 259954
rect 114250 259718 114486 259954
rect 114570 259718 114806 259954
rect 113930 259398 114166 259634
rect 114250 259398 114486 259634
rect 114570 259398 114806 259634
rect 133930 259718 134166 259954
rect 134250 259718 134486 259954
rect 134570 259718 134806 259954
rect 133930 259398 134166 259634
rect 134250 259398 134486 259634
rect 134570 259398 134806 259634
rect 153930 259718 154166 259954
rect 154250 259718 154486 259954
rect 154570 259718 154806 259954
rect 153930 259398 154166 259634
rect 154250 259398 154486 259634
rect 154570 259398 154806 259634
rect 173930 259718 174166 259954
rect 174250 259718 174486 259954
rect 174570 259718 174806 259954
rect 173930 259398 174166 259634
rect 174250 259398 174486 259634
rect 174570 259398 174806 259634
rect 193930 259718 194166 259954
rect 194250 259718 194486 259954
rect 194570 259718 194806 259954
rect 193930 259398 194166 259634
rect 194250 259398 194486 259634
rect 194570 259398 194806 259634
rect 213930 259718 214166 259954
rect 214250 259718 214486 259954
rect 214570 259718 214806 259954
rect 213930 259398 214166 259634
rect 214250 259398 214486 259634
rect 214570 259398 214806 259634
rect 233930 259718 234166 259954
rect 234250 259718 234486 259954
rect 234570 259718 234806 259954
rect 233930 259398 234166 259634
rect 234250 259398 234486 259634
rect 234570 259398 234806 259634
rect 253930 259718 254166 259954
rect 254250 259718 254486 259954
rect 254570 259718 254806 259954
rect 253930 259398 254166 259634
rect 254250 259398 254486 259634
rect 254570 259398 254806 259634
rect 273930 259718 274166 259954
rect 274250 259718 274486 259954
rect 274570 259718 274806 259954
rect 273930 259398 274166 259634
rect 274250 259398 274486 259634
rect 274570 259398 274806 259634
rect 23930 255218 24166 255454
rect 24250 255218 24486 255454
rect 24570 255218 24806 255454
rect 23930 254898 24166 255134
rect 24250 254898 24486 255134
rect 24570 254898 24806 255134
rect 43930 255218 44166 255454
rect 44250 255218 44486 255454
rect 44570 255218 44806 255454
rect 43930 254898 44166 255134
rect 44250 254898 44486 255134
rect 44570 254898 44806 255134
rect 63930 255218 64166 255454
rect 64250 255218 64486 255454
rect 64570 255218 64806 255454
rect 63930 254898 64166 255134
rect 64250 254898 64486 255134
rect 64570 254898 64806 255134
rect 83930 255218 84166 255454
rect 84250 255218 84486 255454
rect 84570 255218 84806 255454
rect 83930 254898 84166 255134
rect 84250 254898 84486 255134
rect 84570 254898 84806 255134
rect 103930 255218 104166 255454
rect 104250 255218 104486 255454
rect 104570 255218 104806 255454
rect 103930 254898 104166 255134
rect 104250 254898 104486 255134
rect 104570 254898 104806 255134
rect 123930 255218 124166 255454
rect 124250 255218 124486 255454
rect 124570 255218 124806 255454
rect 123930 254898 124166 255134
rect 124250 254898 124486 255134
rect 124570 254898 124806 255134
rect 143930 255218 144166 255454
rect 144250 255218 144486 255454
rect 144570 255218 144806 255454
rect 143930 254898 144166 255134
rect 144250 254898 144486 255134
rect 144570 254898 144806 255134
rect 163930 255218 164166 255454
rect 164250 255218 164486 255454
rect 164570 255218 164806 255454
rect 163930 254898 164166 255134
rect 164250 254898 164486 255134
rect 164570 254898 164806 255134
rect 183930 255218 184166 255454
rect 184250 255218 184486 255454
rect 184570 255218 184806 255454
rect 183930 254898 184166 255134
rect 184250 254898 184486 255134
rect 184570 254898 184806 255134
rect 203930 255218 204166 255454
rect 204250 255218 204486 255454
rect 204570 255218 204806 255454
rect 203930 254898 204166 255134
rect 204250 254898 204486 255134
rect 204570 254898 204806 255134
rect 223930 255218 224166 255454
rect 224250 255218 224486 255454
rect 224570 255218 224806 255454
rect 223930 254898 224166 255134
rect 224250 254898 224486 255134
rect 224570 254898 224806 255134
rect 243930 255218 244166 255454
rect 244250 255218 244486 255454
rect 244570 255218 244806 255454
rect 243930 254898 244166 255134
rect 244250 254898 244486 255134
rect 244570 254898 244806 255134
rect 263930 255218 264166 255454
rect 264250 255218 264486 255454
rect 264570 255218 264806 255454
rect 263930 254898 264166 255134
rect 264250 254898 264486 255134
rect 264570 254898 264806 255134
rect 283930 255218 284166 255454
rect 284250 255218 284486 255454
rect 284570 255218 284806 255454
rect 283930 254898 284166 255134
rect 284250 254898 284486 255134
rect 284570 254898 284806 255134
rect 33930 223718 34166 223954
rect 34250 223718 34486 223954
rect 34570 223718 34806 223954
rect 33930 223398 34166 223634
rect 34250 223398 34486 223634
rect 34570 223398 34806 223634
rect 53930 223718 54166 223954
rect 54250 223718 54486 223954
rect 54570 223718 54806 223954
rect 53930 223398 54166 223634
rect 54250 223398 54486 223634
rect 54570 223398 54806 223634
rect 73930 223718 74166 223954
rect 74250 223718 74486 223954
rect 74570 223718 74806 223954
rect 73930 223398 74166 223634
rect 74250 223398 74486 223634
rect 74570 223398 74806 223634
rect 93930 223718 94166 223954
rect 94250 223718 94486 223954
rect 94570 223718 94806 223954
rect 93930 223398 94166 223634
rect 94250 223398 94486 223634
rect 94570 223398 94806 223634
rect 113930 223718 114166 223954
rect 114250 223718 114486 223954
rect 114570 223718 114806 223954
rect 113930 223398 114166 223634
rect 114250 223398 114486 223634
rect 114570 223398 114806 223634
rect 133930 223718 134166 223954
rect 134250 223718 134486 223954
rect 134570 223718 134806 223954
rect 133930 223398 134166 223634
rect 134250 223398 134486 223634
rect 134570 223398 134806 223634
rect 153930 223718 154166 223954
rect 154250 223718 154486 223954
rect 154570 223718 154806 223954
rect 153930 223398 154166 223634
rect 154250 223398 154486 223634
rect 154570 223398 154806 223634
rect 173930 223718 174166 223954
rect 174250 223718 174486 223954
rect 174570 223718 174806 223954
rect 173930 223398 174166 223634
rect 174250 223398 174486 223634
rect 174570 223398 174806 223634
rect 193930 223718 194166 223954
rect 194250 223718 194486 223954
rect 194570 223718 194806 223954
rect 193930 223398 194166 223634
rect 194250 223398 194486 223634
rect 194570 223398 194806 223634
rect 213930 223718 214166 223954
rect 214250 223718 214486 223954
rect 214570 223718 214806 223954
rect 213930 223398 214166 223634
rect 214250 223398 214486 223634
rect 214570 223398 214806 223634
rect 233930 223718 234166 223954
rect 234250 223718 234486 223954
rect 234570 223718 234806 223954
rect 233930 223398 234166 223634
rect 234250 223398 234486 223634
rect 234570 223398 234806 223634
rect 253930 223718 254166 223954
rect 254250 223718 254486 223954
rect 254570 223718 254806 223954
rect 253930 223398 254166 223634
rect 254250 223398 254486 223634
rect 254570 223398 254806 223634
rect 273930 223718 274166 223954
rect 274250 223718 274486 223954
rect 274570 223718 274806 223954
rect 273930 223398 274166 223634
rect 274250 223398 274486 223634
rect 274570 223398 274806 223634
rect 23930 219218 24166 219454
rect 24250 219218 24486 219454
rect 24570 219218 24806 219454
rect 23930 218898 24166 219134
rect 24250 218898 24486 219134
rect 24570 218898 24806 219134
rect 43930 219218 44166 219454
rect 44250 219218 44486 219454
rect 44570 219218 44806 219454
rect 43930 218898 44166 219134
rect 44250 218898 44486 219134
rect 44570 218898 44806 219134
rect 63930 219218 64166 219454
rect 64250 219218 64486 219454
rect 64570 219218 64806 219454
rect 63930 218898 64166 219134
rect 64250 218898 64486 219134
rect 64570 218898 64806 219134
rect 83930 219218 84166 219454
rect 84250 219218 84486 219454
rect 84570 219218 84806 219454
rect 83930 218898 84166 219134
rect 84250 218898 84486 219134
rect 84570 218898 84806 219134
rect 103930 219218 104166 219454
rect 104250 219218 104486 219454
rect 104570 219218 104806 219454
rect 103930 218898 104166 219134
rect 104250 218898 104486 219134
rect 104570 218898 104806 219134
rect 123930 219218 124166 219454
rect 124250 219218 124486 219454
rect 124570 219218 124806 219454
rect 123930 218898 124166 219134
rect 124250 218898 124486 219134
rect 124570 218898 124806 219134
rect 143930 219218 144166 219454
rect 144250 219218 144486 219454
rect 144570 219218 144806 219454
rect 143930 218898 144166 219134
rect 144250 218898 144486 219134
rect 144570 218898 144806 219134
rect 163930 219218 164166 219454
rect 164250 219218 164486 219454
rect 164570 219218 164806 219454
rect 163930 218898 164166 219134
rect 164250 218898 164486 219134
rect 164570 218898 164806 219134
rect 183930 219218 184166 219454
rect 184250 219218 184486 219454
rect 184570 219218 184806 219454
rect 183930 218898 184166 219134
rect 184250 218898 184486 219134
rect 184570 218898 184806 219134
rect 203930 219218 204166 219454
rect 204250 219218 204486 219454
rect 204570 219218 204806 219454
rect 203930 218898 204166 219134
rect 204250 218898 204486 219134
rect 204570 218898 204806 219134
rect 223930 219218 224166 219454
rect 224250 219218 224486 219454
rect 224570 219218 224806 219454
rect 223930 218898 224166 219134
rect 224250 218898 224486 219134
rect 224570 218898 224806 219134
rect 243930 219218 244166 219454
rect 244250 219218 244486 219454
rect 244570 219218 244806 219454
rect 243930 218898 244166 219134
rect 244250 218898 244486 219134
rect 244570 218898 244806 219134
rect 263930 219218 264166 219454
rect 264250 219218 264486 219454
rect 264570 219218 264806 219454
rect 263930 218898 264166 219134
rect 264250 218898 264486 219134
rect 264570 218898 264806 219134
rect 283930 219218 284166 219454
rect 284250 219218 284486 219454
rect 284570 219218 284806 219454
rect 283930 218898 284166 219134
rect 284250 218898 284486 219134
rect 284570 218898 284806 219134
rect 23930 183218 24166 183454
rect 24250 183218 24486 183454
rect 24570 183218 24806 183454
rect 23930 182898 24166 183134
rect 24250 182898 24486 183134
rect 24570 182898 24806 183134
rect 43930 183218 44166 183454
rect 44250 183218 44486 183454
rect 44570 183218 44806 183454
rect 43930 182898 44166 183134
rect 44250 182898 44486 183134
rect 44570 182898 44806 183134
rect 63930 183218 64166 183454
rect 64250 183218 64486 183454
rect 64570 183218 64806 183454
rect 63930 182898 64166 183134
rect 64250 182898 64486 183134
rect 64570 182898 64806 183134
rect 83930 183218 84166 183454
rect 84250 183218 84486 183454
rect 84570 183218 84806 183454
rect 83930 182898 84166 183134
rect 84250 182898 84486 183134
rect 84570 182898 84806 183134
rect 103930 183218 104166 183454
rect 104250 183218 104486 183454
rect 104570 183218 104806 183454
rect 103930 182898 104166 183134
rect 104250 182898 104486 183134
rect 104570 182898 104806 183134
rect 123930 183218 124166 183454
rect 124250 183218 124486 183454
rect 124570 183218 124806 183454
rect 123930 182898 124166 183134
rect 124250 182898 124486 183134
rect 124570 182898 124806 183134
rect 143930 183218 144166 183454
rect 144250 183218 144486 183454
rect 144570 183218 144806 183454
rect 143930 182898 144166 183134
rect 144250 182898 144486 183134
rect 144570 182898 144806 183134
rect 163930 183218 164166 183454
rect 164250 183218 164486 183454
rect 164570 183218 164806 183454
rect 163930 182898 164166 183134
rect 164250 182898 164486 183134
rect 164570 182898 164806 183134
rect 183930 183218 184166 183454
rect 184250 183218 184486 183454
rect 184570 183218 184806 183454
rect 183930 182898 184166 183134
rect 184250 182898 184486 183134
rect 184570 182898 184806 183134
rect 203930 183218 204166 183454
rect 204250 183218 204486 183454
rect 204570 183218 204806 183454
rect 203930 182898 204166 183134
rect 204250 182898 204486 183134
rect 204570 182898 204806 183134
rect 223930 183218 224166 183454
rect 224250 183218 224486 183454
rect 224570 183218 224806 183454
rect 223930 182898 224166 183134
rect 224250 182898 224486 183134
rect 224570 182898 224806 183134
rect 243930 183218 244166 183454
rect 244250 183218 244486 183454
rect 244570 183218 244806 183454
rect 243930 182898 244166 183134
rect 244250 182898 244486 183134
rect 244570 182898 244806 183134
rect 263930 183218 264166 183454
rect 264250 183218 264486 183454
rect 264570 183218 264806 183454
rect 263930 182898 264166 183134
rect 264250 182898 264486 183134
rect 264570 182898 264806 183134
rect 283930 183218 284166 183454
rect 284250 183218 284486 183454
rect 284570 183218 284806 183454
rect 283930 182898 284166 183134
rect 284250 182898 284486 183134
rect 284570 182898 284806 183134
rect 33930 151718 34166 151954
rect 34250 151718 34486 151954
rect 34570 151718 34806 151954
rect 33930 151398 34166 151634
rect 34250 151398 34486 151634
rect 34570 151398 34806 151634
rect 53930 151718 54166 151954
rect 54250 151718 54486 151954
rect 54570 151718 54806 151954
rect 53930 151398 54166 151634
rect 54250 151398 54486 151634
rect 54570 151398 54806 151634
rect 73930 151718 74166 151954
rect 74250 151718 74486 151954
rect 74570 151718 74806 151954
rect 73930 151398 74166 151634
rect 74250 151398 74486 151634
rect 74570 151398 74806 151634
rect 93930 151718 94166 151954
rect 94250 151718 94486 151954
rect 94570 151718 94806 151954
rect 93930 151398 94166 151634
rect 94250 151398 94486 151634
rect 94570 151398 94806 151634
rect 113930 151718 114166 151954
rect 114250 151718 114486 151954
rect 114570 151718 114806 151954
rect 113930 151398 114166 151634
rect 114250 151398 114486 151634
rect 114570 151398 114806 151634
rect 133930 151718 134166 151954
rect 134250 151718 134486 151954
rect 134570 151718 134806 151954
rect 133930 151398 134166 151634
rect 134250 151398 134486 151634
rect 134570 151398 134806 151634
rect 153930 151718 154166 151954
rect 154250 151718 154486 151954
rect 154570 151718 154806 151954
rect 153930 151398 154166 151634
rect 154250 151398 154486 151634
rect 154570 151398 154806 151634
rect 173930 151718 174166 151954
rect 174250 151718 174486 151954
rect 174570 151718 174806 151954
rect 173930 151398 174166 151634
rect 174250 151398 174486 151634
rect 174570 151398 174806 151634
rect 193930 151718 194166 151954
rect 194250 151718 194486 151954
rect 194570 151718 194806 151954
rect 193930 151398 194166 151634
rect 194250 151398 194486 151634
rect 194570 151398 194806 151634
rect 213930 151718 214166 151954
rect 214250 151718 214486 151954
rect 214570 151718 214806 151954
rect 213930 151398 214166 151634
rect 214250 151398 214486 151634
rect 214570 151398 214806 151634
rect 233930 151718 234166 151954
rect 234250 151718 234486 151954
rect 234570 151718 234806 151954
rect 233930 151398 234166 151634
rect 234250 151398 234486 151634
rect 234570 151398 234806 151634
rect 253930 151718 254166 151954
rect 254250 151718 254486 151954
rect 254570 151718 254806 151954
rect 253930 151398 254166 151634
rect 254250 151398 254486 151634
rect 254570 151398 254806 151634
rect 273930 151718 274166 151954
rect 274250 151718 274486 151954
rect 274570 151718 274806 151954
rect 273930 151398 274166 151634
rect 274250 151398 274486 151634
rect 274570 151398 274806 151634
rect 23930 147218 24166 147454
rect 24250 147218 24486 147454
rect 24570 147218 24806 147454
rect 23930 146898 24166 147134
rect 24250 146898 24486 147134
rect 24570 146898 24806 147134
rect 43930 147218 44166 147454
rect 44250 147218 44486 147454
rect 44570 147218 44806 147454
rect 43930 146898 44166 147134
rect 44250 146898 44486 147134
rect 44570 146898 44806 147134
rect 63930 147218 64166 147454
rect 64250 147218 64486 147454
rect 64570 147218 64806 147454
rect 63930 146898 64166 147134
rect 64250 146898 64486 147134
rect 64570 146898 64806 147134
rect 83930 147218 84166 147454
rect 84250 147218 84486 147454
rect 84570 147218 84806 147454
rect 83930 146898 84166 147134
rect 84250 146898 84486 147134
rect 84570 146898 84806 147134
rect 103930 147218 104166 147454
rect 104250 147218 104486 147454
rect 104570 147218 104806 147454
rect 103930 146898 104166 147134
rect 104250 146898 104486 147134
rect 104570 146898 104806 147134
rect 123930 147218 124166 147454
rect 124250 147218 124486 147454
rect 124570 147218 124806 147454
rect 123930 146898 124166 147134
rect 124250 146898 124486 147134
rect 124570 146898 124806 147134
rect 143930 147218 144166 147454
rect 144250 147218 144486 147454
rect 144570 147218 144806 147454
rect 143930 146898 144166 147134
rect 144250 146898 144486 147134
rect 144570 146898 144806 147134
rect 163930 147218 164166 147454
rect 164250 147218 164486 147454
rect 164570 147218 164806 147454
rect 163930 146898 164166 147134
rect 164250 146898 164486 147134
rect 164570 146898 164806 147134
rect 183930 147218 184166 147454
rect 184250 147218 184486 147454
rect 184570 147218 184806 147454
rect 183930 146898 184166 147134
rect 184250 146898 184486 147134
rect 184570 146898 184806 147134
rect 203930 147218 204166 147454
rect 204250 147218 204486 147454
rect 204570 147218 204806 147454
rect 203930 146898 204166 147134
rect 204250 146898 204486 147134
rect 204570 146898 204806 147134
rect 223930 147218 224166 147454
rect 224250 147218 224486 147454
rect 224570 147218 224806 147454
rect 223930 146898 224166 147134
rect 224250 146898 224486 147134
rect 224570 146898 224806 147134
rect 243930 147218 244166 147454
rect 244250 147218 244486 147454
rect 244570 147218 244806 147454
rect 243930 146898 244166 147134
rect 244250 146898 244486 147134
rect 244570 146898 244806 147134
rect 263930 147218 264166 147454
rect 264250 147218 264486 147454
rect 264570 147218 264806 147454
rect 263930 146898 264166 147134
rect 264250 146898 264486 147134
rect 264570 146898 264806 147134
rect 283930 147218 284166 147454
rect 284250 147218 284486 147454
rect 284570 147218 284806 147454
rect 283930 146898 284166 147134
rect 284250 146898 284486 147134
rect 284570 146898 284806 147134
rect 33930 115718 34166 115954
rect 34250 115718 34486 115954
rect 34570 115718 34806 115954
rect 33930 115398 34166 115634
rect 34250 115398 34486 115634
rect 34570 115398 34806 115634
rect 53930 115718 54166 115954
rect 54250 115718 54486 115954
rect 54570 115718 54806 115954
rect 53930 115398 54166 115634
rect 54250 115398 54486 115634
rect 54570 115398 54806 115634
rect 73930 115718 74166 115954
rect 74250 115718 74486 115954
rect 74570 115718 74806 115954
rect 73930 115398 74166 115634
rect 74250 115398 74486 115634
rect 74570 115398 74806 115634
rect 93930 115718 94166 115954
rect 94250 115718 94486 115954
rect 94570 115718 94806 115954
rect 93930 115398 94166 115634
rect 94250 115398 94486 115634
rect 94570 115398 94806 115634
rect 113930 115718 114166 115954
rect 114250 115718 114486 115954
rect 114570 115718 114806 115954
rect 113930 115398 114166 115634
rect 114250 115398 114486 115634
rect 114570 115398 114806 115634
rect 133930 115718 134166 115954
rect 134250 115718 134486 115954
rect 134570 115718 134806 115954
rect 133930 115398 134166 115634
rect 134250 115398 134486 115634
rect 134570 115398 134806 115634
rect 153930 115718 154166 115954
rect 154250 115718 154486 115954
rect 154570 115718 154806 115954
rect 153930 115398 154166 115634
rect 154250 115398 154486 115634
rect 154570 115398 154806 115634
rect 173930 115718 174166 115954
rect 174250 115718 174486 115954
rect 174570 115718 174806 115954
rect 173930 115398 174166 115634
rect 174250 115398 174486 115634
rect 174570 115398 174806 115634
rect 193930 115718 194166 115954
rect 194250 115718 194486 115954
rect 194570 115718 194806 115954
rect 193930 115398 194166 115634
rect 194250 115398 194486 115634
rect 194570 115398 194806 115634
rect 213930 115718 214166 115954
rect 214250 115718 214486 115954
rect 214570 115718 214806 115954
rect 213930 115398 214166 115634
rect 214250 115398 214486 115634
rect 214570 115398 214806 115634
rect 233930 115718 234166 115954
rect 234250 115718 234486 115954
rect 234570 115718 234806 115954
rect 233930 115398 234166 115634
rect 234250 115398 234486 115634
rect 234570 115398 234806 115634
rect 253930 115718 254166 115954
rect 254250 115718 254486 115954
rect 254570 115718 254806 115954
rect 253930 115398 254166 115634
rect 254250 115398 254486 115634
rect 254570 115398 254806 115634
rect 273930 115718 274166 115954
rect 274250 115718 274486 115954
rect 274570 115718 274806 115954
rect 273930 115398 274166 115634
rect 274250 115398 274486 115634
rect 274570 115398 274806 115634
rect 23930 111218 24166 111454
rect 24250 111218 24486 111454
rect 24570 111218 24806 111454
rect 23930 110898 24166 111134
rect 24250 110898 24486 111134
rect 24570 110898 24806 111134
rect 43930 111218 44166 111454
rect 44250 111218 44486 111454
rect 44570 111218 44806 111454
rect 43930 110898 44166 111134
rect 44250 110898 44486 111134
rect 44570 110898 44806 111134
rect 63930 111218 64166 111454
rect 64250 111218 64486 111454
rect 64570 111218 64806 111454
rect 63930 110898 64166 111134
rect 64250 110898 64486 111134
rect 64570 110898 64806 111134
rect 83930 111218 84166 111454
rect 84250 111218 84486 111454
rect 84570 111218 84806 111454
rect 83930 110898 84166 111134
rect 84250 110898 84486 111134
rect 84570 110898 84806 111134
rect 103930 111218 104166 111454
rect 104250 111218 104486 111454
rect 104570 111218 104806 111454
rect 103930 110898 104166 111134
rect 104250 110898 104486 111134
rect 104570 110898 104806 111134
rect 123930 111218 124166 111454
rect 124250 111218 124486 111454
rect 124570 111218 124806 111454
rect 123930 110898 124166 111134
rect 124250 110898 124486 111134
rect 124570 110898 124806 111134
rect 143930 111218 144166 111454
rect 144250 111218 144486 111454
rect 144570 111218 144806 111454
rect 143930 110898 144166 111134
rect 144250 110898 144486 111134
rect 144570 110898 144806 111134
rect 163930 111218 164166 111454
rect 164250 111218 164486 111454
rect 164570 111218 164806 111454
rect 163930 110898 164166 111134
rect 164250 110898 164486 111134
rect 164570 110898 164806 111134
rect 183930 111218 184166 111454
rect 184250 111218 184486 111454
rect 184570 111218 184806 111454
rect 183930 110898 184166 111134
rect 184250 110898 184486 111134
rect 184570 110898 184806 111134
rect 203930 111218 204166 111454
rect 204250 111218 204486 111454
rect 204570 111218 204806 111454
rect 203930 110898 204166 111134
rect 204250 110898 204486 111134
rect 204570 110898 204806 111134
rect 223930 111218 224166 111454
rect 224250 111218 224486 111454
rect 224570 111218 224806 111454
rect 223930 110898 224166 111134
rect 224250 110898 224486 111134
rect 224570 110898 224806 111134
rect 243930 111218 244166 111454
rect 244250 111218 244486 111454
rect 244570 111218 244806 111454
rect 243930 110898 244166 111134
rect 244250 110898 244486 111134
rect 244570 110898 244806 111134
rect 263930 111218 264166 111454
rect 264250 111218 264486 111454
rect 264570 111218 264806 111454
rect 263930 110898 264166 111134
rect 264250 110898 264486 111134
rect 264570 110898 264806 111134
rect 283930 111218 284166 111454
rect 284250 111218 284486 111454
rect 284570 111218 284806 111454
rect 283930 110898 284166 111134
rect 284250 110898 284486 111134
rect 284570 110898 284806 111134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 79610 43718 79846 43954
rect 79610 43398 79846 43634
rect 64250 39218 64486 39454
rect 64250 38898 64486 39134
rect 94970 39218 95206 39454
rect 94970 38898 95206 39134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 313930 691718 314166 691954
rect 314250 691718 314486 691954
rect 314570 691718 314806 691954
rect 313930 691398 314166 691634
rect 314250 691398 314486 691634
rect 314570 691398 314806 691634
rect 333930 691718 334166 691954
rect 334250 691718 334486 691954
rect 334570 691718 334806 691954
rect 333930 691398 334166 691634
rect 334250 691398 334486 691634
rect 334570 691398 334806 691634
rect 353930 691718 354166 691954
rect 354250 691718 354486 691954
rect 354570 691718 354806 691954
rect 353930 691398 354166 691634
rect 354250 691398 354486 691634
rect 354570 691398 354806 691634
rect 373930 691718 374166 691954
rect 374250 691718 374486 691954
rect 374570 691718 374806 691954
rect 373930 691398 374166 691634
rect 374250 691398 374486 691634
rect 374570 691398 374806 691634
rect 393930 691718 394166 691954
rect 394250 691718 394486 691954
rect 394570 691718 394806 691954
rect 393930 691398 394166 691634
rect 394250 691398 394486 691634
rect 394570 691398 394806 691634
rect 413930 691718 414166 691954
rect 414250 691718 414486 691954
rect 414570 691718 414806 691954
rect 413930 691398 414166 691634
rect 414250 691398 414486 691634
rect 414570 691398 414806 691634
rect 433930 691718 434166 691954
rect 434250 691718 434486 691954
rect 434570 691718 434806 691954
rect 433930 691398 434166 691634
rect 434250 691398 434486 691634
rect 434570 691398 434806 691634
rect 453930 691718 454166 691954
rect 454250 691718 454486 691954
rect 454570 691718 454806 691954
rect 453930 691398 454166 691634
rect 454250 691398 454486 691634
rect 454570 691398 454806 691634
rect 473930 691718 474166 691954
rect 474250 691718 474486 691954
rect 474570 691718 474806 691954
rect 473930 691398 474166 691634
rect 474250 691398 474486 691634
rect 474570 691398 474806 691634
rect 493930 691718 494166 691954
rect 494250 691718 494486 691954
rect 494570 691718 494806 691954
rect 493930 691398 494166 691634
rect 494250 691398 494486 691634
rect 494570 691398 494806 691634
rect 513930 691718 514166 691954
rect 514250 691718 514486 691954
rect 514570 691718 514806 691954
rect 513930 691398 514166 691634
rect 514250 691398 514486 691634
rect 514570 691398 514806 691634
rect 533930 691718 534166 691954
rect 534250 691718 534486 691954
rect 534570 691718 534806 691954
rect 533930 691398 534166 691634
rect 534250 691398 534486 691634
rect 534570 691398 534806 691634
rect 553930 691718 554166 691954
rect 554250 691718 554486 691954
rect 554570 691718 554806 691954
rect 553930 691398 554166 691634
rect 554250 691398 554486 691634
rect 554570 691398 554806 691634
rect 303930 687218 304166 687454
rect 304250 687218 304486 687454
rect 304570 687218 304806 687454
rect 303930 686898 304166 687134
rect 304250 686898 304486 687134
rect 304570 686898 304806 687134
rect 323930 687218 324166 687454
rect 324250 687218 324486 687454
rect 324570 687218 324806 687454
rect 323930 686898 324166 687134
rect 324250 686898 324486 687134
rect 324570 686898 324806 687134
rect 343930 687218 344166 687454
rect 344250 687218 344486 687454
rect 344570 687218 344806 687454
rect 343930 686898 344166 687134
rect 344250 686898 344486 687134
rect 344570 686898 344806 687134
rect 363930 687218 364166 687454
rect 364250 687218 364486 687454
rect 364570 687218 364806 687454
rect 363930 686898 364166 687134
rect 364250 686898 364486 687134
rect 364570 686898 364806 687134
rect 383930 687218 384166 687454
rect 384250 687218 384486 687454
rect 384570 687218 384806 687454
rect 383930 686898 384166 687134
rect 384250 686898 384486 687134
rect 384570 686898 384806 687134
rect 403930 687218 404166 687454
rect 404250 687218 404486 687454
rect 404570 687218 404806 687454
rect 403930 686898 404166 687134
rect 404250 686898 404486 687134
rect 404570 686898 404806 687134
rect 423930 687218 424166 687454
rect 424250 687218 424486 687454
rect 424570 687218 424806 687454
rect 423930 686898 424166 687134
rect 424250 686898 424486 687134
rect 424570 686898 424806 687134
rect 443930 687218 444166 687454
rect 444250 687218 444486 687454
rect 444570 687218 444806 687454
rect 443930 686898 444166 687134
rect 444250 686898 444486 687134
rect 444570 686898 444806 687134
rect 463930 687218 464166 687454
rect 464250 687218 464486 687454
rect 464570 687218 464806 687454
rect 463930 686898 464166 687134
rect 464250 686898 464486 687134
rect 464570 686898 464806 687134
rect 483930 687218 484166 687454
rect 484250 687218 484486 687454
rect 484570 687218 484806 687454
rect 483930 686898 484166 687134
rect 484250 686898 484486 687134
rect 484570 686898 484806 687134
rect 503930 687218 504166 687454
rect 504250 687218 504486 687454
rect 504570 687218 504806 687454
rect 503930 686898 504166 687134
rect 504250 686898 504486 687134
rect 504570 686898 504806 687134
rect 523930 687218 524166 687454
rect 524250 687218 524486 687454
rect 524570 687218 524806 687454
rect 523930 686898 524166 687134
rect 524250 686898 524486 687134
rect 524570 686898 524806 687134
rect 543930 687218 544166 687454
rect 544250 687218 544486 687454
rect 544570 687218 544806 687454
rect 543930 686898 544166 687134
rect 544250 686898 544486 687134
rect 544570 686898 544806 687134
rect 563930 687218 564166 687454
rect 564250 687218 564486 687454
rect 564570 687218 564806 687454
rect 563930 686898 564166 687134
rect 564250 686898 564486 687134
rect 564570 686898 564806 687134
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 313930 655718 314166 655954
rect 314250 655718 314486 655954
rect 314570 655718 314806 655954
rect 313930 655398 314166 655634
rect 314250 655398 314486 655634
rect 314570 655398 314806 655634
rect 333930 655718 334166 655954
rect 334250 655718 334486 655954
rect 334570 655718 334806 655954
rect 333930 655398 334166 655634
rect 334250 655398 334486 655634
rect 334570 655398 334806 655634
rect 353930 655718 354166 655954
rect 354250 655718 354486 655954
rect 354570 655718 354806 655954
rect 353930 655398 354166 655634
rect 354250 655398 354486 655634
rect 354570 655398 354806 655634
rect 373930 655718 374166 655954
rect 374250 655718 374486 655954
rect 374570 655718 374806 655954
rect 373930 655398 374166 655634
rect 374250 655398 374486 655634
rect 374570 655398 374806 655634
rect 393930 655718 394166 655954
rect 394250 655718 394486 655954
rect 394570 655718 394806 655954
rect 393930 655398 394166 655634
rect 394250 655398 394486 655634
rect 394570 655398 394806 655634
rect 413930 655718 414166 655954
rect 414250 655718 414486 655954
rect 414570 655718 414806 655954
rect 413930 655398 414166 655634
rect 414250 655398 414486 655634
rect 414570 655398 414806 655634
rect 433930 655718 434166 655954
rect 434250 655718 434486 655954
rect 434570 655718 434806 655954
rect 433930 655398 434166 655634
rect 434250 655398 434486 655634
rect 434570 655398 434806 655634
rect 453930 655718 454166 655954
rect 454250 655718 454486 655954
rect 454570 655718 454806 655954
rect 453930 655398 454166 655634
rect 454250 655398 454486 655634
rect 454570 655398 454806 655634
rect 473930 655718 474166 655954
rect 474250 655718 474486 655954
rect 474570 655718 474806 655954
rect 473930 655398 474166 655634
rect 474250 655398 474486 655634
rect 474570 655398 474806 655634
rect 493930 655718 494166 655954
rect 494250 655718 494486 655954
rect 494570 655718 494806 655954
rect 493930 655398 494166 655634
rect 494250 655398 494486 655634
rect 494570 655398 494806 655634
rect 513930 655718 514166 655954
rect 514250 655718 514486 655954
rect 514570 655718 514806 655954
rect 513930 655398 514166 655634
rect 514250 655398 514486 655634
rect 514570 655398 514806 655634
rect 533930 655718 534166 655954
rect 534250 655718 534486 655954
rect 534570 655718 534806 655954
rect 533930 655398 534166 655634
rect 534250 655398 534486 655634
rect 534570 655398 534806 655634
rect 553930 655718 554166 655954
rect 554250 655718 554486 655954
rect 554570 655718 554806 655954
rect 553930 655398 554166 655634
rect 554250 655398 554486 655634
rect 554570 655398 554806 655634
rect 303930 651218 304166 651454
rect 304250 651218 304486 651454
rect 304570 651218 304806 651454
rect 303930 650898 304166 651134
rect 304250 650898 304486 651134
rect 304570 650898 304806 651134
rect 323930 651218 324166 651454
rect 324250 651218 324486 651454
rect 324570 651218 324806 651454
rect 323930 650898 324166 651134
rect 324250 650898 324486 651134
rect 324570 650898 324806 651134
rect 343930 651218 344166 651454
rect 344250 651218 344486 651454
rect 344570 651218 344806 651454
rect 343930 650898 344166 651134
rect 344250 650898 344486 651134
rect 344570 650898 344806 651134
rect 363930 651218 364166 651454
rect 364250 651218 364486 651454
rect 364570 651218 364806 651454
rect 363930 650898 364166 651134
rect 364250 650898 364486 651134
rect 364570 650898 364806 651134
rect 383930 651218 384166 651454
rect 384250 651218 384486 651454
rect 384570 651218 384806 651454
rect 383930 650898 384166 651134
rect 384250 650898 384486 651134
rect 384570 650898 384806 651134
rect 403930 651218 404166 651454
rect 404250 651218 404486 651454
rect 404570 651218 404806 651454
rect 403930 650898 404166 651134
rect 404250 650898 404486 651134
rect 404570 650898 404806 651134
rect 423930 651218 424166 651454
rect 424250 651218 424486 651454
rect 424570 651218 424806 651454
rect 423930 650898 424166 651134
rect 424250 650898 424486 651134
rect 424570 650898 424806 651134
rect 443930 651218 444166 651454
rect 444250 651218 444486 651454
rect 444570 651218 444806 651454
rect 443930 650898 444166 651134
rect 444250 650898 444486 651134
rect 444570 650898 444806 651134
rect 463930 651218 464166 651454
rect 464250 651218 464486 651454
rect 464570 651218 464806 651454
rect 463930 650898 464166 651134
rect 464250 650898 464486 651134
rect 464570 650898 464806 651134
rect 483930 651218 484166 651454
rect 484250 651218 484486 651454
rect 484570 651218 484806 651454
rect 483930 650898 484166 651134
rect 484250 650898 484486 651134
rect 484570 650898 484806 651134
rect 503930 651218 504166 651454
rect 504250 651218 504486 651454
rect 504570 651218 504806 651454
rect 503930 650898 504166 651134
rect 504250 650898 504486 651134
rect 504570 650898 504806 651134
rect 523930 651218 524166 651454
rect 524250 651218 524486 651454
rect 524570 651218 524806 651454
rect 523930 650898 524166 651134
rect 524250 650898 524486 651134
rect 524570 650898 524806 651134
rect 543930 651218 544166 651454
rect 544250 651218 544486 651454
rect 544570 651218 544806 651454
rect 543930 650898 544166 651134
rect 544250 650898 544486 651134
rect 544570 650898 544806 651134
rect 563930 651218 564166 651454
rect 564250 651218 564486 651454
rect 564570 651218 564806 651454
rect 563930 650898 564166 651134
rect 564250 650898 564486 651134
rect 564570 650898 564806 651134
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 313930 619718 314166 619954
rect 314250 619718 314486 619954
rect 314570 619718 314806 619954
rect 313930 619398 314166 619634
rect 314250 619398 314486 619634
rect 314570 619398 314806 619634
rect 333930 619718 334166 619954
rect 334250 619718 334486 619954
rect 334570 619718 334806 619954
rect 333930 619398 334166 619634
rect 334250 619398 334486 619634
rect 334570 619398 334806 619634
rect 353930 619718 354166 619954
rect 354250 619718 354486 619954
rect 354570 619718 354806 619954
rect 353930 619398 354166 619634
rect 354250 619398 354486 619634
rect 354570 619398 354806 619634
rect 373930 619718 374166 619954
rect 374250 619718 374486 619954
rect 374570 619718 374806 619954
rect 373930 619398 374166 619634
rect 374250 619398 374486 619634
rect 374570 619398 374806 619634
rect 393930 619718 394166 619954
rect 394250 619718 394486 619954
rect 394570 619718 394806 619954
rect 393930 619398 394166 619634
rect 394250 619398 394486 619634
rect 394570 619398 394806 619634
rect 413930 619718 414166 619954
rect 414250 619718 414486 619954
rect 414570 619718 414806 619954
rect 413930 619398 414166 619634
rect 414250 619398 414486 619634
rect 414570 619398 414806 619634
rect 433930 619718 434166 619954
rect 434250 619718 434486 619954
rect 434570 619718 434806 619954
rect 433930 619398 434166 619634
rect 434250 619398 434486 619634
rect 434570 619398 434806 619634
rect 453930 619718 454166 619954
rect 454250 619718 454486 619954
rect 454570 619718 454806 619954
rect 453930 619398 454166 619634
rect 454250 619398 454486 619634
rect 454570 619398 454806 619634
rect 473930 619718 474166 619954
rect 474250 619718 474486 619954
rect 474570 619718 474806 619954
rect 473930 619398 474166 619634
rect 474250 619398 474486 619634
rect 474570 619398 474806 619634
rect 493930 619718 494166 619954
rect 494250 619718 494486 619954
rect 494570 619718 494806 619954
rect 493930 619398 494166 619634
rect 494250 619398 494486 619634
rect 494570 619398 494806 619634
rect 513930 619718 514166 619954
rect 514250 619718 514486 619954
rect 514570 619718 514806 619954
rect 513930 619398 514166 619634
rect 514250 619398 514486 619634
rect 514570 619398 514806 619634
rect 533930 619718 534166 619954
rect 534250 619718 534486 619954
rect 534570 619718 534806 619954
rect 533930 619398 534166 619634
rect 534250 619398 534486 619634
rect 534570 619398 534806 619634
rect 553930 619718 554166 619954
rect 554250 619718 554486 619954
rect 554570 619718 554806 619954
rect 553930 619398 554166 619634
rect 554250 619398 554486 619634
rect 554570 619398 554806 619634
rect 303930 615218 304166 615454
rect 304250 615218 304486 615454
rect 304570 615218 304806 615454
rect 303930 614898 304166 615134
rect 304250 614898 304486 615134
rect 304570 614898 304806 615134
rect 323930 615218 324166 615454
rect 324250 615218 324486 615454
rect 324570 615218 324806 615454
rect 323930 614898 324166 615134
rect 324250 614898 324486 615134
rect 324570 614898 324806 615134
rect 343930 615218 344166 615454
rect 344250 615218 344486 615454
rect 344570 615218 344806 615454
rect 343930 614898 344166 615134
rect 344250 614898 344486 615134
rect 344570 614898 344806 615134
rect 363930 615218 364166 615454
rect 364250 615218 364486 615454
rect 364570 615218 364806 615454
rect 363930 614898 364166 615134
rect 364250 614898 364486 615134
rect 364570 614898 364806 615134
rect 383930 615218 384166 615454
rect 384250 615218 384486 615454
rect 384570 615218 384806 615454
rect 383930 614898 384166 615134
rect 384250 614898 384486 615134
rect 384570 614898 384806 615134
rect 403930 615218 404166 615454
rect 404250 615218 404486 615454
rect 404570 615218 404806 615454
rect 403930 614898 404166 615134
rect 404250 614898 404486 615134
rect 404570 614898 404806 615134
rect 423930 615218 424166 615454
rect 424250 615218 424486 615454
rect 424570 615218 424806 615454
rect 423930 614898 424166 615134
rect 424250 614898 424486 615134
rect 424570 614898 424806 615134
rect 443930 615218 444166 615454
rect 444250 615218 444486 615454
rect 444570 615218 444806 615454
rect 443930 614898 444166 615134
rect 444250 614898 444486 615134
rect 444570 614898 444806 615134
rect 463930 615218 464166 615454
rect 464250 615218 464486 615454
rect 464570 615218 464806 615454
rect 463930 614898 464166 615134
rect 464250 614898 464486 615134
rect 464570 614898 464806 615134
rect 483930 615218 484166 615454
rect 484250 615218 484486 615454
rect 484570 615218 484806 615454
rect 483930 614898 484166 615134
rect 484250 614898 484486 615134
rect 484570 614898 484806 615134
rect 503930 615218 504166 615454
rect 504250 615218 504486 615454
rect 504570 615218 504806 615454
rect 503930 614898 504166 615134
rect 504250 614898 504486 615134
rect 504570 614898 504806 615134
rect 523930 615218 524166 615454
rect 524250 615218 524486 615454
rect 524570 615218 524806 615454
rect 523930 614898 524166 615134
rect 524250 614898 524486 615134
rect 524570 614898 524806 615134
rect 543930 615218 544166 615454
rect 544250 615218 544486 615454
rect 544570 615218 544806 615454
rect 543930 614898 544166 615134
rect 544250 614898 544486 615134
rect 544570 614898 544806 615134
rect 563930 615218 564166 615454
rect 564250 615218 564486 615454
rect 564570 615218 564806 615454
rect 563930 614898 564166 615134
rect 564250 614898 564486 615134
rect 564570 614898 564806 615134
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 313930 547718 314166 547954
rect 314250 547718 314486 547954
rect 314570 547718 314806 547954
rect 313930 547398 314166 547634
rect 314250 547398 314486 547634
rect 314570 547398 314806 547634
rect 333930 547718 334166 547954
rect 334250 547718 334486 547954
rect 334570 547718 334806 547954
rect 333930 547398 334166 547634
rect 334250 547398 334486 547634
rect 334570 547398 334806 547634
rect 353930 547718 354166 547954
rect 354250 547718 354486 547954
rect 354570 547718 354806 547954
rect 353930 547398 354166 547634
rect 354250 547398 354486 547634
rect 354570 547398 354806 547634
rect 373930 547718 374166 547954
rect 374250 547718 374486 547954
rect 374570 547718 374806 547954
rect 373930 547398 374166 547634
rect 374250 547398 374486 547634
rect 374570 547398 374806 547634
rect 393930 547718 394166 547954
rect 394250 547718 394486 547954
rect 394570 547718 394806 547954
rect 393930 547398 394166 547634
rect 394250 547398 394486 547634
rect 394570 547398 394806 547634
rect 413930 547718 414166 547954
rect 414250 547718 414486 547954
rect 414570 547718 414806 547954
rect 413930 547398 414166 547634
rect 414250 547398 414486 547634
rect 414570 547398 414806 547634
rect 433930 547718 434166 547954
rect 434250 547718 434486 547954
rect 434570 547718 434806 547954
rect 433930 547398 434166 547634
rect 434250 547398 434486 547634
rect 434570 547398 434806 547634
rect 453930 547718 454166 547954
rect 454250 547718 454486 547954
rect 454570 547718 454806 547954
rect 453930 547398 454166 547634
rect 454250 547398 454486 547634
rect 454570 547398 454806 547634
rect 473930 547718 474166 547954
rect 474250 547718 474486 547954
rect 474570 547718 474806 547954
rect 473930 547398 474166 547634
rect 474250 547398 474486 547634
rect 474570 547398 474806 547634
rect 493930 547718 494166 547954
rect 494250 547718 494486 547954
rect 494570 547718 494806 547954
rect 493930 547398 494166 547634
rect 494250 547398 494486 547634
rect 494570 547398 494806 547634
rect 513930 547718 514166 547954
rect 514250 547718 514486 547954
rect 514570 547718 514806 547954
rect 513930 547398 514166 547634
rect 514250 547398 514486 547634
rect 514570 547398 514806 547634
rect 533930 547718 534166 547954
rect 534250 547718 534486 547954
rect 534570 547718 534806 547954
rect 533930 547398 534166 547634
rect 534250 547398 534486 547634
rect 534570 547398 534806 547634
rect 553930 547718 554166 547954
rect 554250 547718 554486 547954
rect 554570 547718 554806 547954
rect 553930 547398 554166 547634
rect 554250 547398 554486 547634
rect 554570 547398 554806 547634
rect 303930 543218 304166 543454
rect 304250 543218 304486 543454
rect 304570 543218 304806 543454
rect 303930 542898 304166 543134
rect 304250 542898 304486 543134
rect 304570 542898 304806 543134
rect 323930 543218 324166 543454
rect 324250 543218 324486 543454
rect 324570 543218 324806 543454
rect 323930 542898 324166 543134
rect 324250 542898 324486 543134
rect 324570 542898 324806 543134
rect 343930 543218 344166 543454
rect 344250 543218 344486 543454
rect 344570 543218 344806 543454
rect 343930 542898 344166 543134
rect 344250 542898 344486 543134
rect 344570 542898 344806 543134
rect 363930 543218 364166 543454
rect 364250 543218 364486 543454
rect 364570 543218 364806 543454
rect 363930 542898 364166 543134
rect 364250 542898 364486 543134
rect 364570 542898 364806 543134
rect 383930 543218 384166 543454
rect 384250 543218 384486 543454
rect 384570 543218 384806 543454
rect 383930 542898 384166 543134
rect 384250 542898 384486 543134
rect 384570 542898 384806 543134
rect 403930 543218 404166 543454
rect 404250 543218 404486 543454
rect 404570 543218 404806 543454
rect 403930 542898 404166 543134
rect 404250 542898 404486 543134
rect 404570 542898 404806 543134
rect 423930 543218 424166 543454
rect 424250 543218 424486 543454
rect 424570 543218 424806 543454
rect 423930 542898 424166 543134
rect 424250 542898 424486 543134
rect 424570 542898 424806 543134
rect 443930 543218 444166 543454
rect 444250 543218 444486 543454
rect 444570 543218 444806 543454
rect 443930 542898 444166 543134
rect 444250 542898 444486 543134
rect 444570 542898 444806 543134
rect 463930 543218 464166 543454
rect 464250 543218 464486 543454
rect 464570 543218 464806 543454
rect 463930 542898 464166 543134
rect 464250 542898 464486 543134
rect 464570 542898 464806 543134
rect 483930 543218 484166 543454
rect 484250 543218 484486 543454
rect 484570 543218 484806 543454
rect 483930 542898 484166 543134
rect 484250 542898 484486 543134
rect 484570 542898 484806 543134
rect 503930 543218 504166 543454
rect 504250 543218 504486 543454
rect 504570 543218 504806 543454
rect 503930 542898 504166 543134
rect 504250 542898 504486 543134
rect 504570 542898 504806 543134
rect 523930 543218 524166 543454
rect 524250 543218 524486 543454
rect 524570 543218 524806 543454
rect 523930 542898 524166 543134
rect 524250 542898 524486 543134
rect 524570 542898 524806 543134
rect 543930 543218 544166 543454
rect 544250 543218 544486 543454
rect 544570 543218 544806 543454
rect 543930 542898 544166 543134
rect 544250 542898 544486 543134
rect 544570 542898 544806 543134
rect 563930 543218 564166 543454
rect 564250 543218 564486 543454
rect 564570 543218 564806 543454
rect 563930 542898 564166 543134
rect 564250 542898 564486 543134
rect 564570 542898 564806 543134
rect 313930 511718 314166 511954
rect 314250 511718 314486 511954
rect 314570 511718 314806 511954
rect 313930 511398 314166 511634
rect 314250 511398 314486 511634
rect 314570 511398 314806 511634
rect 333930 511718 334166 511954
rect 334250 511718 334486 511954
rect 334570 511718 334806 511954
rect 333930 511398 334166 511634
rect 334250 511398 334486 511634
rect 334570 511398 334806 511634
rect 353930 511718 354166 511954
rect 354250 511718 354486 511954
rect 354570 511718 354806 511954
rect 353930 511398 354166 511634
rect 354250 511398 354486 511634
rect 354570 511398 354806 511634
rect 373930 511718 374166 511954
rect 374250 511718 374486 511954
rect 374570 511718 374806 511954
rect 373930 511398 374166 511634
rect 374250 511398 374486 511634
rect 374570 511398 374806 511634
rect 393930 511718 394166 511954
rect 394250 511718 394486 511954
rect 394570 511718 394806 511954
rect 393930 511398 394166 511634
rect 394250 511398 394486 511634
rect 394570 511398 394806 511634
rect 413930 511718 414166 511954
rect 414250 511718 414486 511954
rect 414570 511718 414806 511954
rect 413930 511398 414166 511634
rect 414250 511398 414486 511634
rect 414570 511398 414806 511634
rect 433930 511718 434166 511954
rect 434250 511718 434486 511954
rect 434570 511718 434806 511954
rect 433930 511398 434166 511634
rect 434250 511398 434486 511634
rect 434570 511398 434806 511634
rect 453930 511718 454166 511954
rect 454250 511718 454486 511954
rect 454570 511718 454806 511954
rect 453930 511398 454166 511634
rect 454250 511398 454486 511634
rect 454570 511398 454806 511634
rect 473930 511718 474166 511954
rect 474250 511718 474486 511954
rect 474570 511718 474806 511954
rect 473930 511398 474166 511634
rect 474250 511398 474486 511634
rect 474570 511398 474806 511634
rect 493930 511718 494166 511954
rect 494250 511718 494486 511954
rect 494570 511718 494806 511954
rect 493930 511398 494166 511634
rect 494250 511398 494486 511634
rect 494570 511398 494806 511634
rect 513930 511718 514166 511954
rect 514250 511718 514486 511954
rect 514570 511718 514806 511954
rect 513930 511398 514166 511634
rect 514250 511398 514486 511634
rect 514570 511398 514806 511634
rect 533930 511718 534166 511954
rect 534250 511718 534486 511954
rect 534570 511718 534806 511954
rect 533930 511398 534166 511634
rect 534250 511398 534486 511634
rect 534570 511398 534806 511634
rect 553930 511718 554166 511954
rect 554250 511718 554486 511954
rect 554570 511718 554806 511954
rect 553930 511398 554166 511634
rect 554250 511398 554486 511634
rect 554570 511398 554806 511634
rect 303930 507218 304166 507454
rect 304250 507218 304486 507454
rect 304570 507218 304806 507454
rect 303930 506898 304166 507134
rect 304250 506898 304486 507134
rect 304570 506898 304806 507134
rect 323930 507218 324166 507454
rect 324250 507218 324486 507454
rect 324570 507218 324806 507454
rect 323930 506898 324166 507134
rect 324250 506898 324486 507134
rect 324570 506898 324806 507134
rect 343930 507218 344166 507454
rect 344250 507218 344486 507454
rect 344570 507218 344806 507454
rect 343930 506898 344166 507134
rect 344250 506898 344486 507134
rect 344570 506898 344806 507134
rect 363930 507218 364166 507454
rect 364250 507218 364486 507454
rect 364570 507218 364806 507454
rect 363930 506898 364166 507134
rect 364250 506898 364486 507134
rect 364570 506898 364806 507134
rect 383930 507218 384166 507454
rect 384250 507218 384486 507454
rect 384570 507218 384806 507454
rect 383930 506898 384166 507134
rect 384250 506898 384486 507134
rect 384570 506898 384806 507134
rect 403930 507218 404166 507454
rect 404250 507218 404486 507454
rect 404570 507218 404806 507454
rect 403930 506898 404166 507134
rect 404250 506898 404486 507134
rect 404570 506898 404806 507134
rect 423930 507218 424166 507454
rect 424250 507218 424486 507454
rect 424570 507218 424806 507454
rect 423930 506898 424166 507134
rect 424250 506898 424486 507134
rect 424570 506898 424806 507134
rect 443930 507218 444166 507454
rect 444250 507218 444486 507454
rect 444570 507218 444806 507454
rect 443930 506898 444166 507134
rect 444250 506898 444486 507134
rect 444570 506898 444806 507134
rect 463930 507218 464166 507454
rect 464250 507218 464486 507454
rect 464570 507218 464806 507454
rect 463930 506898 464166 507134
rect 464250 506898 464486 507134
rect 464570 506898 464806 507134
rect 483930 507218 484166 507454
rect 484250 507218 484486 507454
rect 484570 507218 484806 507454
rect 483930 506898 484166 507134
rect 484250 506898 484486 507134
rect 484570 506898 484806 507134
rect 503930 507218 504166 507454
rect 504250 507218 504486 507454
rect 504570 507218 504806 507454
rect 503930 506898 504166 507134
rect 504250 506898 504486 507134
rect 504570 506898 504806 507134
rect 523930 507218 524166 507454
rect 524250 507218 524486 507454
rect 524570 507218 524806 507454
rect 523930 506898 524166 507134
rect 524250 506898 524486 507134
rect 524570 506898 524806 507134
rect 543930 507218 544166 507454
rect 544250 507218 544486 507454
rect 544570 507218 544806 507454
rect 543930 506898 544166 507134
rect 544250 506898 544486 507134
rect 544570 506898 544806 507134
rect 563930 507218 564166 507454
rect 564250 507218 564486 507454
rect 564570 507218 564806 507454
rect 563930 506898 564166 507134
rect 564250 506898 564486 507134
rect 564570 506898 564806 507134
rect 313930 475718 314166 475954
rect 314250 475718 314486 475954
rect 314570 475718 314806 475954
rect 313930 475398 314166 475634
rect 314250 475398 314486 475634
rect 314570 475398 314806 475634
rect 333930 475718 334166 475954
rect 334250 475718 334486 475954
rect 334570 475718 334806 475954
rect 333930 475398 334166 475634
rect 334250 475398 334486 475634
rect 334570 475398 334806 475634
rect 353930 475718 354166 475954
rect 354250 475718 354486 475954
rect 354570 475718 354806 475954
rect 353930 475398 354166 475634
rect 354250 475398 354486 475634
rect 354570 475398 354806 475634
rect 373930 475718 374166 475954
rect 374250 475718 374486 475954
rect 374570 475718 374806 475954
rect 373930 475398 374166 475634
rect 374250 475398 374486 475634
rect 374570 475398 374806 475634
rect 393930 475718 394166 475954
rect 394250 475718 394486 475954
rect 394570 475718 394806 475954
rect 393930 475398 394166 475634
rect 394250 475398 394486 475634
rect 394570 475398 394806 475634
rect 413930 475718 414166 475954
rect 414250 475718 414486 475954
rect 414570 475718 414806 475954
rect 413930 475398 414166 475634
rect 414250 475398 414486 475634
rect 414570 475398 414806 475634
rect 433930 475718 434166 475954
rect 434250 475718 434486 475954
rect 434570 475718 434806 475954
rect 433930 475398 434166 475634
rect 434250 475398 434486 475634
rect 434570 475398 434806 475634
rect 453930 475718 454166 475954
rect 454250 475718 454486 475954
rect 454570 475718 454806 475954
rect 453930 475398 454166 475634
rect 454250 475398 454486 475634
rect 454570 475398 454806 475634
rect 473930 475718 474166 475954
rect 474250 475718 474486 475954
rect 474570 475718 474806 475954
rect 473930 475398 474166 475634
rect 474250 475398 474486 475634
rect 474570 475398 474806 475634
rect 493930 475718 494166 475954
rect 494250 475718 494486 475954
rect 494570 475718 494806 475954
rect 493930 475398 494166 475634
rect 494250 475398 494486 475634
rect 494570 475398 494806 475634
rect 513930 475718 514166 475954
rect 514250 475718 514486 475954
rect 514570 475718 514806 475954
rect 513930 475398 514166 475634
rect 514250 475398 514486 475634
rect 514570 475398 514806 475634
rect 533930 475718 534166 475954
rect 534250 475718 534486 475954
rect 534570 475718 534806 475954
rect 533930 475398 534166 475634
rect 534250 475398 534486 475634
rect 534570 475398 534806 475634
rect 553930 475718 554166 475954
rect 554250 475718 554486 475954
rect 554570 475718 554806 475954
rect 553930 475398 554166 475634
rect 554250 475398 554486 475634
rect 554570 475398 554806 475634
rect 303930 471218 304166 471454
rect 304250 471218 304486 471454
rect 304570 471218 304806 471454
rect 303930 470898 304166 471134
rect 304250 470898 304486 471134
rect 304570 470898 304806 471134
rect 323930 471218 324166 471454
rect 324250 471218 324486 471454
rect 324570 471218 324806 471454
rect 323930 470898 324166 471134
rect 324250 470898 324486 471134
rect 324570 470898 324806 471134
rect 343930 471218 344166 471454
rect 344250 471218 344486 471454
rect 344570 471218 344806 471454
rect 343930 470898 344166 471134
rect 344250 470898 344486 471134
rect 344570 470898 344806 471134
rect 363930 471218 364166 471454
rect 364250 471218 364486 471454
rect 364570 471218 364806 471454
rect 363930 470898 364166 471134
rect 364250 470898 364486 471134
rect 364570 470898 364806 471134
rect 383930 471218 384166 471454
rect 384250 471218 384486 471454
rect 384570 471218 384806 471454
rect 383930 470898 384166 471134
rect 384250 470898 384486 471134
rect 384570 470898 384806 471134
rect 403930 471218 404166 471454
rect 404250 471218 404486 471454
rect 404570 471218 404806 471454
rect 403930 470898 404166 471134
rect 404250 470898 404486 471134
rect 404570 470898 404806 471134
rect 423930 471218 424166 471454
rect 424250 471218 424486 471454
rect 424570 471218 424806 471454
rect 423930 470898 424166 471134
rect 424250 470898 424486 471134
rect 424570 470898 424806 471134
rect 443930 471218 444166 471454
rect 444250 471218 444486 471454
rect 444570 471218 444806 471454
rect 443930 470898 444166 471134
rect 444250 470898 444486 471134
rect 444570 470898 444806 471134
rect 463930 471218 464166 471454
rect 464250 471218 464486 471454
rect 464570 471218 464806 471454
rect 463930 470898 464166 471134
rect 464250 470898 464486 471134
rect 464570 470898 464806 471134
rect 483930 471218 484166 471454
rect 484250 471218 484486 471454
rect 484570 471218 484806 471454
rect 483930 470898 484166 471134
rect 484250 470898 484486 471134
rect 484570 470898 484806 471134
rect 503930 471218 504166 471454
rect 504250 471218 504486 471454
rect 504570 471218 504806 471454
rect 503930 470898 504166 471134
rect 504250 470898 504486 471134
rect 504570 470898 504806 471134
rect 523930 471218 524166 471454
rect 524250 471218 524486 471454
rect 524570 471218 524806 471454
rect 523930 470898 524166 471134
rect 524250 470898 524486 471134
rect 524570 470898 524806 471134
rect 543930 471218 544166 471454
rect 544250 471218 544486 471454
rect 544570 471218 544806 471454
rect 543930 470898 544166 471134
rect 544250 470898 544486 471134
rect 544570 470898 544806 471134
rect 563930 471218 564166 471454
rect 564250 471218 564486 471454
rect 564570 471218 564806 471454
rect 563930 470898 564166 471134
rect 564250 470898 564486 471134
rect 564570 470898 564806 471134
rect 313930 439718 314166 439954
rect 314250 439718 314486 439954
rect 314570 439718 314806 439954
rect 313930 439398 314166 439634
rect 314250 439398 314486 439634
rect 314570 439398 314806 439634
rect 333930 439718 334166 439954
rect 334250 439718 334486 439954
rect 334570 439718 334806 439954
rect 333930 439398 334166 439634
rect 334250 439398 334486 439634
rect 334570 439398 334806 439634
rect 353930 439718 354166 439954
rect 354250 439718 354486 439954
rect 354570 439718 354806 439954
rect 353930 439398 354166 439634
rect 354250 439398 354486 439634
rect 354570 439398 354806 439634
rect 373930 439718 374166 439954
rect 374250 439718 374486 439954
rect 374570 439718 374806 439954
rect 373930 439398 374166 439634
rect 374250 439398 374486 439634
rect 374570 439398 374806 439634
rect 393930 439718 394166 439954
rect 394250 439718 394486 439954
rect 394570 439718 394806 439954
rect 393930 439398 394166 439634
rect 394250 439398 394486 439634
rect 394570 439398 394806 439634
rect 413930 439718 414166 439954
rect 414250 439718 414486 439954
rect 414570 439718 414806 439954
rect 413930 439398 414166 439634
rect 414250 439398 414486 439634
rect 414570 439398 414806 439634
rect 433930 439718 434166 439954
rect 434250 439718 434486 439954
rect 434570 439718 434806 439954
rect 433930 439398 434166 439634
rect 434250 439398 434486 439634
rect 434570 439398 434806 439634
rect 453930 439718 454166 439954
rect 454250 439718 454486 439954
rect 454570 439718 454806 439954
rect 453930 439398 454166 439634
rect 454250 439398 454486 439634
rect 454570 439398 454806 439634
rect 473930 439718 474166 439954
rect 474250 439718 474486 439954
rect 474570 439718 474806 439954
rect 473930 439398 474166 439634
rect 474250 439398 474486 439634
rect 474570 439398 474806 439634
rect 493930 439718 494166 439954
rect 494250 439718 494486 439954
rect 494570 439718 494806 439954
rect 493930 439398 494166 439634
rect 494250 439398 494486 439634
rect 494570 439398 494806 439634
rect 513930 439718 514166 439954
rect 514250 439718 514486 439954
rect 514570 439718 514806 439954
rect 513930 439398 514166 439634
rect 514250 439398 514486 439634
rect 514570 439398 514806 439634
rect 533930 439718 534166 439954
rect 534250 439718 534486 439954
rect 534570 439718 534806 439954
rect 533930 439398 534166 439634
rect 534250 439398 534486 439634
rect 534570 439398 534806 439634
rect 553930 439718 554166 439954
rect 554250 439718 554486 439954
rect 554570 439718 554806 439954
rect 553930 439398 554166 439634
rect 554250 439398 554486 439634
rect 554570 439398 554806 439634
rect 303930 435218 304166 435454
rect 304250 435218 304486 435454
rect 304570 435218 304806 435454
rect 303930 434898 304166 435134
rect 304250 434898 304486 435134
rect 304570 434898 304806 435134
rect 323930 435218 324166 435454
rect 324250 435218 324486 435454
rect 324570 435218 324806 435454
rect 323930 434898 324166 435134
rect 324250 434898 324486 435134
rect 324570 434898 324806 435134
rect 343930 435218 344166 435454
rect 344250 435218 344486 435454
rect 344570 435218 344806 435454
rect 343930 434898 344166 435134
rect 344250 434898 344486 435134
rect 344570 434898 344806 435134
rect 363930 435218 364166 435454
rect 364250 435218 364486 435454
rect 364570 435218 364806 435454
rect 363930 434898 364166 435134
rect 364250 434898 364486 435134
rect 364570 434898 364806 435134
rect 383930 435218 384166 435454
rect 384250 435218 384486 435454
rect 384570 435218 384806 435454
rect 383930 434898 384166 435134
rect 384250 434898 384486 435134
rect 384570 434898 384806 435134
rect 403930 435218 404166 435454
rect 404250 435218 404486 435454
rect 404570 435218 404806 435454
rect 403930 434898 404166 435134
rect 404250 434898 404486 435134
rect 404570 434898 404806 435134
rect 423930 435218 424166 435454
rect 424250 435218 424486 435454
rect 424570 435218 424806 435454
rect 423930 434898 424166 435134
rect 424250 434898 424486 435134
rect 424570 434898 424806 435134
rect 443930 435218 444166 435454
rect 444250 435218 444486 435454
rect 444570 435218 444806 435454
rect 443930 434898 444166 435134
rect 444250 434898 444486 435134
rect 444570 434898 444806 435134
rect 463930 435218 464166 435454
rect 464250 435218 464486 435454
rect 464570 435218 464806 435454
rect 463930 434898 464166 435134
rect 464250 434898 464486 435134
rect 464570 434898 464806 435134
rect 483930 435218 484166 435454
rect 484250 435218 484486 435454
rect 484570 435218 484806 435454
rect 483930 434898 484166 435134
rect 484250 434898 484486 435134
rect 484570 434898 484806 435134
rect 503930 435218 504166 435454
rect 504250 435218 504486 435454
rect 504570 435218 504806 435454
rect 503930 434898 504166 435134
rect 504250 434898 504486 435134
rect 504570 434898 504806 435134
rect 523930 435218 524166 435454
rect 524250 435218 524486 435454
rect 524570 435218 524806 435454
rect 523930 434898 524166 435134
rect 524250 434898 524486 435134
rect 524570 434898 524806 435134
rect 543930 435218 544166 435454
rect 544250 435218 544486 435454
rect 544570 435218 544806 435454
rect 543930 434898 544166 435134
rect 544250 434898 544486 435134
rect 544570 434898 544806 435134
rect 563930 435218 564166 435454
rect 564250 435218 564486 435454
rect 564570 435218 564806 435454
rect 563930 434898 564166 435134
rect 564250 434898 564486 435134
rect 564570 434898 564806 435134
rect 313930 403718 314166 403954
rect 314250 403718 314486 403954
rect 314570 403718 314806 403954
rect 313930 403398 314166 403634
rect 314250 403398 314486 403634
rect 314570 403398 314806 403634
rect 333930 403718 334166 403954
rect 334250 403718 334486 403954
rect 334570 403718 334806 403954
rect 333930 403398 334166 403634
rect 334250 403398 334486 403634
rect 334570 403398 334806 403634
rect 353930 403718 354166 403954
rect 354250 403718 354486 403954
rect 354570 403718 354806 403954
rect 353930 403398 354166 403634
rect 354250 403398 354486 403634
rect 354570 403398 354806 403634
rect 373930 403718 374166 403954
rect 374250 403718 374486 403954
rect 374570 403718 374806 403954
rect 373930 403398 374166 403634
rect 374250 403398 374486 403634
rect 374570 403398 374806 403634
rect 393930 403718 394166 403954
rect 394250 403718 394486 403954
rect 394570 403718 394806 403954
rect 393930 403398 394166 403634
rect 394250 403398 394486 403634
rect 394570 403398 394806 403634
rect 413930 403718 414166 403954
rect 414250 403718 414486 403954
rect 414570 403718 414806 403954
rect 413930 403398 414166 403634
rect 414250 403398 414486 403634
rect 414570 403398 414806 403634
rect 433930 403718 434166 403954
rect 434250 403718 434486 403954
rect 434570 403718 434806 403954
rect 433930 403398 434166 403634
rect 434250 403398 434486 403634
rect 434570 403398 434806 403634
rect 453930 403718 454166 403954
rect 454250 403718 454486 403954
rect 454570 403718 454806 403954
rect 453930 403398 454166 403634
rect 454250 403398 454486 403634
rect 454570 403398 454806 403634
rect 473930 403718 474166 403954
rect 474250 403718 474486 403954
rect 474570 403718 474806 403954
rect 473930 403398 474166 403634
rect 474250 403398 474486 403634
rect 474570 403398 474806 403634
rect 493930 403718 494166 403954
rect 494250 403718 494486 403954
rect 494570 403718 494806 403954
rect 493930 403398 494166 403634
rect 494250 403398 494486 403634
rect 494570 403398 494806 403634
rect 513930 403718 514166 403954
rect 514250 403718 514486 403954
rect 514570 403718 514806 403954
rect 513930 403398 514166 403634
rect 514250 403398 514486 403634
rect 514570 403398 514806 403634
rect 533930 403718 534166 403954
rect 534250 403718 534486 403954
rect 534570 403718 534806 403954
rect 533930 403398 534166 403634
rect 534250 403398 534486 403634
rect 534570 403398 534806 403634
rect 553930 403718 554166 403954
rect 554250 403718 554486 403954
rect 554570 403718 554806 403954
rect 553930 403398 554166 403634
rect 554250 403398 554486 403634
rect 554570 403398 554806 403634
rect 303930 399218 304166 399454
rect 304250 399218 304486 399454
rect 304570 399218 304806 399454
rect 303930 398898 304166 399134
rect 304250 398898 304486 399134
rect 304570 398898 304806 399134
rect 323930 399218 324166 399454
rect 324250 399218 324486 399454
rect 324570 399218 324806 399454
rect 323930 398898 324166 399134
rect 324250 398898 324486 399134
rect 324570 398898 324806 399134
rect 343930 399218 344166 399454
rect 344250 399218 344486 399454
rect 344570 399218 344806 399454
rect 343930 398898 344166 399134
rect 344250 398898 344486 399134
rect 344570 398898 344806 399134
rect 363930 399218 364166 399454
rect 364250 399218 364486 399454
rect 364570 399218 364806 399454
rect 363930 398898 364166 399134
rect 364250 398898 364486 399134
rect 364570 398898 364806 399134
rect 383930 399218 384166 399454
rect 384250 399218 384486 399454
rect 384570 399218 384806 399454
rect 383930 398898 384166 399134
rect 384250 398898 384486 399134
rect 384570 398898 384806 399134
rect 403930 399218 404166 399454
rect 404250 399218 404486 399454
rect 404570 399218 404806 399454
rect 403930 398898 404166 399134
rect 404250 398898 404486 399134
rect 404570 398898 404806 399134
rect 423930 399218 424166 399454
rect 424250 399218 424486 399454
rect 424570 399218 424806 399454
rect 423930 398898 424166 399134
rect 424250 398898 424486 399134
rect 424570 398898 424806 399134
rect 443930 399218 444166 399454
rect 444250 399218 444486 399454
rect 444570 399218 444806 399454
rect 443930 398898 444166 399134
rect 444250 398898 444486 399134
rect 444570 398898 444806 399134
rect 463930 399218 464166 399454
rect 464250 399218 464486 399454
rect 464570 399218 464806 399454
rect 463930 398898 464166 399134
rect 464250 398898 464486 399134
rect 464570 398898 464806 399134
rect 483930 399218 484166 399454
rect 484250 399218 484486 399454
rect 484570 399218 484806 399454
rect 483930 398898 484166 399134
rect 484250 398898 484486 399134
rect 484570 398898 484806 399134
rect 503930 399218 504166 399454
rect 504250 399218 504486 399454
rect 504570 399218 504806 399454
rect 503930 398898 504166 399134
rect 504250 398898 504486 399134
rect 504570 398898 504806 399134
rect 523930 399218 524166 399454
rect 524250 399218 524486 399454
rect 524570 399218 524806 399454
rect 523930 398898 524166 399134
rect 524250 398898 524486 399134
rect 524570 398898 524806 399134
rect 543930 399218 544166 399454
rect 544250 399218 544486 399454
rect 544570 399218 544806 399454
rect 543930 398898 544166 399134
rect 544250 398898 544486 399134
rect 544570 398898 544806 399134
rect 563930 399218 564166 399454
rect 564250 399218 564486 399454
rect 564570 399218 564806 399454
rect 563930 398898 564166 399134
rect 564250 398898 564486 399134
rect 564570 398898 564806 399134
rect 313930 367718 314166 367954
rect 314250 367718 314486 367954
rect 314570 367718 314806 367954
rect 313930 367398 314166 367634
rect 314250 367398 314486 367634
rect 314570 367398 314806 367634
rect 333930 367718 334166 367954
rect 334250 367718 334486 367954
rect 334570 367718 334806 367954
rect 333930 367398 334166 367634
rect 334250 367398 334486 367634
rect 334570 367398 334806 367634
rect 353930 367718 354166 367954
rect 354250 367718 354486 367954
rect 354570 367718 354806 367954
rect 353930 367398 354166 367634
rect 354250 367398 354486 367634
rect 354570 367398 354806 367634
rect 373930 367718 374166 367954
rect 374250 367718 374486 367954
rect 374570 367718 374806 367954
rect 373930 367398 374166 367634
rect 374250 367398 374486 367634
rect 374570 367398 374806 367634
rect 393930 367718 394166 367954
rect 394250 367718 394486 367954
rect 394570 367718 394806 367954
rect 393930 367398 394166 367634
rect 394250 367398 394486 367634
rect 394570 367398 394806 367634
rect 413930 367718 414166 367954
rect 414250 367718 414486 367954
rect 414570 367718 414806 367954
rect 413930 367398 414166 367634
rect 414250 367398 414486 367634
rect 414570 367398 414806 367634
rect 433930 367718 434166 367954
rect 434250 367718 434486 367954
rect 434570 367718 434806 367954
rect 433930 367398 434166 367634
rect 434250 367398 434486 367634
rect 434570 367398 434806 367634
rect 453930 367718 454166 367954
rect 454250 367718 454486 367954
rect 454570 367718 454806 367954
rect 453930 367398 454166 367634
rect 454250 367398 454486 367634
rect 454570 367398 454806 367634
rect 473930 367718 474166 367954
rect 474250 367718 474486 367954
rect 474570 367718 474806 367954
rect 473930 367398 474166 367634
rect 474250 367398 474486 367634
rect 474570 367398 474806 367634
rect 493930 367718 494166 367954
rect 494250 367718 494486 367954
rect 494570 367718 494806 367954
rect 493930 367398 494166 367634
rect 494250 367398 494486 367634
rect 494570 367398 494806 367634
rect 513930 367718 514166 367954
rect 514250 367718 514486 367954
rect 514570 367718 514806 367954
rect 513930 367398 514166 367634
rect 514250 367398 514486 367634
rect 514570 367398 514806 367634
rect 533930 367718 534166 367954
rect 534250 367718 534486 367954
rect 534570 367718 534806 367954
rect 533930 367398 534166 367634
rect 534250 367398 534486 367634
rect 534570 367398 534806 367634
rect 553930 367718 554166 367954
rect 554250 367718 554486 367954
rect 554570 367718 554806 367954
rect 553930 367398 554166 367634
rect 554250 367398 554486 367634
rect 554570 367398 554806 367634
rect 303930 363218 304166 363454
rect 304250 363218 304486 363454
rect 304570 363218 304806 363454
rect 303930 362898 304166 363134
rect 304250 362898 304486 363134
rect 304570 362898 304806 363134
rect 323930 363218 324166 363454
rect 324250 363218 324486 363454
rect 324570 363218 324806 363454
rect 323930 362898 324166 363134
rect 324250 362898 324486 363134
rect 324570 362898 324806 363134
rect 343930 363218 344166 363454
rect 344250 363218 344486 363454
rect 344570 363218 344806 363454
rect 343930 362898 344166 363134
rect 344250 362898 344486 363134
rect 344570 362898 344806 363134
rect 363930 363218 364166 363454
rect 364250 363218 364486 363454
rect 364570 363218 364806 363454
rect 363930 362898 364166 363134
rect 364250 362898 364486 363134
rect 364570 362898 364806 363134
rect 383930 363218 384166 363454
rect 384250 363218 384486 363454
rect 384570 363218 384806 363454
rect 383930 362898 384166 363134
rect 384250 362898 384486 363134
rect 384570 362898 384806 363134
rect 403930 363218 404166 363454
rect 404250 363218 404486 363454
rect 404570 363218 404806 363454
rect 403930 362898 404166 363134
rect 404250 362898 404486 363134
rect 404570 362898 404806 363134
rect 423930 363218 424166 363454
rect 424250 363218 424486 363454
rect 424570 363218 424806 363454
rect 423930 362898 424166 363134
rect 424250 362898 424486 363134
rect 424570 362898 424806 363134
rect 443930 363218 444166 363454
rect 444250 363218 444486 363454
rect 444570 363218 444806 363454
rect 443930 362898 444166 363134
rect 444250 362898 444486 363134
rect 444570 362898 444806 363134
rect 463930 363218 464166 363454
rect 464250 363218 464486 363454
rect 464570 363218 464806 363454
rect 463930 362898 464166 363134
rect 464250 362898 464486 363134
rect 464570 362898 464806 363134
rect 483930 363218 484166 363454
rect 484250 363218 484486 363454
rect 484570 363218 484806 363454
rect 483930 362898 484166 363134
rect 484250 362898 484486 363134
rect 484570 362898 484806 363134
rect 503930 363218 504166 363454
rect 504250 363218 504486 363454
rect 504570 363218 504806 363454
rect 503930 362898 504166 363134
rect 504250 362898 504486 363134
rect 504570 362898 504806 363134
rect 523930 363218 524166 363454
rect 524250 363218 524486 363454
rect 524570 363218 524806 363454
rect 523930 362898 524166 363134
rect 524250 362898 524486 363134
rect 524570 362898 524806 363134
rect 543930 363218 544166 363454
rect 544250 363218 544486 363454
rect 544570 363218 544806 363454
rect 543930 362898 544166 363134
rect 544250 362898 544486 363134
rect 544570 362898 544806 363134
rect 563930 363218 564166 363454
rect 564250 363218 564486 363454
rect 564570 363218 564806 363454
rect 563930 362898 564166 363134
rect 564250 362898 564486 363134
rect 564570 362898 564806 363134
rect 313930 295718 314166 295954
rect 314250 295718 314486 295954
rect 314570 295718 314806 295954
rect 313930 295398 314166 295634
rect 314250 295398 314486 295634
rect 314570 295398 314806 295634
rect 333930 295718 334166 295954
rect 334250 295718 334486 295954
rect 334570 295718 334806 295954
rect 333930 295398 334166 295634
rect 334250 295398 334486 295634
rect 334570 295398 334806 295634
rect 353930 295718 354166 295954
rect 354250 295718 354486 295954
rect 354570 295718 354806 295954
rect 353930 295398 354166 295634
rect 354250 295398 354486 295634
rect 354570 295398 354806 295634
rect 373930 295718 374166 295954
rect 374250 295718 374486 295954
rect 374570 295718 374806 295954
rect 373930 295398 374166 295634
rect 374250 295398 374486 295634
rect 374570 295398 374806 295634
rect 393930 295718 394166 295954
rect 394250 295718 394486 295954
rect 394570 295718 394806 295954
rect 393930 295398 394166 295634
rect 394250 295398 394486 295634
rect 394570 295398 394806 295634
rect 413930 295718 414166 295954
rect 414250 295718 414486 295954
rect 414570 295718 414806 295954
rect 413930 295398 414166 295634
rect 414250 295398 414486 295634
rect 414570 295398 414806 295634
rect 433930 295718 434166 295954
rect 434250 295718 434486 295954
rect 434570 295718 434806 295954
rect 433930 295398 434166 295634
rect 434250 295398 434486 295634
rect 434570 295398 434806 295634
rect 453930 295718 454166 295954
rect 454250 295718 454486 295954
rect 454570 295718 454806 295954
rect 453930 295398 454166 295634
rect 454250 295398 454486 295634
rect 454570 295398 454806 295634
rect 473930 295718 474166 295954
rect 474250 295718 474486 295954
rect 474570 295718 474806 295954
rect 473930 295398 474166 295634
rect 474250 295398 474486 295634
rect 474570 295398 474806 295634
rect 493930 295718 494166 295954
rect 494250 295718 494486 295954
rect 494570 295718 494806 295954
rect 493930 295398 494166 295634
rect 494250 295398 494486 295634
rect 494570 295398 494806 295634
rect 513930 295718 514166 295954
rect 514250 295718 514486 295954
rect 514570 295718 514806 295954
rect 513930 295398 514166 295634
rect 514250 295398 514486 295634
rect 514570 295398 514806 295634
rect 533930 295718 534166 295954
rect 534250 295718 534486 295954
rect 534570 295718 534806 295954
rect 533930 295398 534166 295634
rect 534250 295398 534486 295634
rect 534570 295398 534806 295634
rect 553930 295718 554166 295954
rect 554250 295718 554486 295954
rect 554570 295718 554806 295954
rect 553930 295398 554166 295634
rect 554250 295398 554486 295634
rect 554570 295398 554806 295634
rect 303930 291218 304166 291454
rect 304250 291218 304486 291454
rect 304570 291218 304806 291454
rect 303930 290898 304166 291134
rect 304250 290898 304486 291134
rect 304570 290898 304806 291134
rect 323930 291218 324166 291454
rect 324250 291218 324486 291454
rect 324570 291218 324806 291454
rect 323930 290898 324166 291134
rect 324250 290898 324486 291134
rect 324570 290898 324806 291134
rect 343930 291218 344166 291454
rect 344250 291218 344486 291454
rect 344570 291218 344806 291454
rect 343930 290898 344166 291134
rect 344250 290898 344486 291134
rect 344570 290898 344806 291134
rect 363930 291218 364166 291454
rect 364250 291218 364486 291454
rect 364570 291218 364806 291454
rect 363930 290898 364166 291134
rect 364250 290898 364486 291134
rect 364570 290898 364806 291134
rect 383930 291218 384166 291454
rect 384250 291218 384486 291454
rect 384570 291218 384806 291454
rect 383930 290898 384166 291134
rect 384250 290898 384486 291134
rect 384570 290898 384806 291134
rect 403930 291218 404166 291454
rect 404250 291218 404486 291454
rect 404570 291218 404806 291454
rect 403930 290898 404166 291134
rect 404250 290898 404486 291134
rect 404570 290898 404806 291134
rect 423930 291218 424166 291454
rect 424250 291218 424486 291454
rect 424570 291218 424806 291454
rect 423930 290898 424166 291134
rect 424250 290898 424486 291134
rect 424570 290898 424806 291134
rect 443930 291218 444166 291454
rect 444250 291218 444486 291454
rect 444570 291218 444806 291454
rect 443930 290898 444166 291134
rect 444250 290898 444486 291134
rect 444570 290898 444806 291134
rect 463930 291218 464166 291454
rect 464250 291218 464486 291454
rect 464570 291218 464806 291454
rect 463930 290898 464166 291134
rect 464250 290898 464486 291134
rect 464570 290898 464806 291134
rect 483930 291218 484166 291454
rect 484250 291218 484486 291454
rect 484570 291218 484806 291454
rect 483930 290898 484166 291134
rect 484250 290898 484486 291134
rect 484570 290898 484806 291134
rect 503930 291218 504166 291454
rect 504250 291218 504486 291454
rect 504570 291218 504806 291454
rect 503930 290898 504166 291134
rect 504250 290898 504486 291134
rect 504570 290898 504806 291134
rect 523930 291218 524166 291454
rect 524250 291218 524486 291454
rect 524570 291218 524806 291454
rect 523930 290898 524166 291134
rect 524250 290898 524486 291134
rect 524570 290898 524806 291134
rect 543930 291218 544166 291454
rect 544250 291218 544486 291454
rect 544570 291218 544806 291454
rect 543930 290898 544166 291134
rect 544250 290898 544486 291134
rect 544570 290898 544806 291134
rect 563930 291218 564166 291454
rect 564250 291218 564486 291454
rect 564570 291218 564806 291454
rect 563930 290898 564166 291134
rect 564250 290898 564486 291134
rect 564570 290898 564806 291134
rect 313930 259718 314166 259954
rect 314250 259718 314486 259954
rect 314570 259718 314806 259954
rect 313930 259398 314166 259634
rect 314250 259398 314486 259634
rect 314570 259398 314806 259634
rect 333930 259718 334166 259954
rect 334250 259718 334486 259954
rect 334570 259718 334806 259954
rect 333930 259398 334166 259634
rect 334250 259398 334486 259634
rect 334570 259398 334806 259634
rect 353930 259718 354166 259954
rect 354250 259718 354486 259954
rect 354570 259718 354806 259954
rect 353930 259398 354166 259634
rect 354250 259398 354486 259634
rect 354570 259398 354806 259634
rect 373930 259718 374166 259954
rect 374250 259718 374486 259954
rect 374570 259718 374806 259954
rect 373930 259398 374166 259634
rect 374250 259398 374486 259634
rect 374570 259398 374806 259634
rect 393930 259718 394166 259954
rect 394250 259718 394486 259954
rect 394570 259718 394806 259954
rect 393930 259398 394166 259634
rect 394250 259398 394486 259634
rect 394570 259398 394806 259634
rect 413930 259718 414166 259954
rect 414250 259718 414486 259954
rect 414570 259718 414806 259954
rect 413930 259398 414166 259634
rect 414250 259398 414486 259634
rect 414570 259398 414806 259634
rect 433930 259718 434166 259954
rect 434250 259718 434486 259954
rect 434570 259718 434806 259954
rect 433930 259398 434166 259634
rect 434250 259398 434486 259634
rect 434570 259398 434806 259634
rect 453930 259718 454166 259954
rect 454250 259718 454486 259954
rect 454570 259718 454806 259954
rect 453930 259398 454166 259634
rect 454250 259398 454486 259634
rect 454570 259398 454806 259634
rect 473930 259718 474166 259954
rect 474250 259718 474486 259954
rect 474570 259718 474806 259954
rect 473930 259398 474166 259634
rect 474250 259398 474486 259634
rect 474570 259398 474806 259634
rect 493930 259718 494166 259954
rect 494250 259718 494486 259954
rect 494570 259718 494806 259954
rect 493930 259398 494166 259634
rect 494250 259398 494486 259634
rect 494570 259398 494806 259634
rect 513930 259718 514166 259954
rect 514250 259718 514486 259954
rect 514570 259718 514806 259954
rect 513930 259398 514166 259634
rect 514250 259398 514486 259634
rect 514570 259398 514806 259634
rect 533930 259718 534166 259954
rect 534250 259718 534486 259954
rect 534570 259718 534806 259954
rect 533930 259398 534166 259634
rect 534250 259398 534486 259634
rect 534570 259398 534806 259634
rect 553930 259718 554166 259954
rect 554250 259718 554486 259954
rect 554570 259718 554806 259954
rect 553930 259398 554166 259634
rect 554250 259398 554486 259634
rect 554570 259398 554806 259634
rect 303930 255218 304166 255454
rect 304250 255218 304486 255454
rect 304570 255218 304806 255454
rect 303930 254898 304166 255134
rect 304250 254898 304486 255134
rect 304570 254898 304806 255134
rect 323930 255218 324166 255454
rect 324250 255218 324486 255454
rect 324570 255218 324806 255454
rect 323930 254898 324166 255134
rect 324250 254898 324486 255134
rect 324570 254898 324806 255134
rect 343930 255218 344166 255454
rect 344250 255218 344486 255454
rect 344570 255218 344806 255454
rect 343930 254898 344166 255134
rect 344250 254898 344486 255134
rect 344570 254898 344806 255134
rect 363930 255218 364166 255454
rect 364250 255218 364486 255454
rect 364570 255218 364806 255454
rect 363930 254898 364166 255134
rect 364250 254898 364486 255134
rect 364570 254898 364806 255134
rect 383930 255218 384166 255454
rect 384250 255218 384486 255454
rect 384570 255218 384806 255454
rect 383930 254898 384166 255134
rect 384250 254898 384486 255134
rect 384570 254898 384806 255134
rect 403930 255218 404166 255454
rect 404250 255218 404486 255454
rect 404570 255218 404806 255454
rect 403930 254898 404166 255134
rect 404250 254898 404486 255134
rect 404570 254898 404806 255134
rect 423930 255218 424166 255454
rect 424250 255218 424486 255454
rect 424570 255218 424806 255454
rect 423930 254898 424166 255134
rect 424250 254898 424486 255134
rect 424570 254898 424806 255134
rect 443930 255218 444166 255454
rect 444250 255218 444486 255454
rect 444570 255218 444806 255454
rect 443930 254898 444166 255134
rect 444250 254898 444486 255134
rect 444570 254898 444806 255134
rect 463930 255218 464166 255454
rect 464250 255218 464486 255454
rect 464570 255218 464806 255454
rect 463930 254898 464166 255134
rect 464250 254898 464486 255134
rect 464570 254898 464806 255134
rect 483930 255218 484166 255454
rect 484250 255218 484486 255454
rect 484570 255218 484806 255454
rect 483930 254898 484166 255134
rect 484250 254898 484486 255134
rect 484570 254898 484806 255134
rect 503930 255218 504166 255454
rect 504250 255218 504486 255454
rect 504570 255218 504806 255454
rect 503930 254898 504166 255134
rect 504250 254898 504486 255134
rect 504570 254898 504806 255134
rect 523930 255218 524166 255454
rect 524250 255218 524486 255454
rect 524570 255218 524806 255454
rect 523930 254898 524166 255134
rect 524250 254898 524486 255134
rect 524570 254898 524806 255134
rect 543930 255218 544166 255454
rect 544250 255218 544486 255454
rect 544570 255218 544806 255454
rect 543930 254898 544166 255134
rect 544250 254898 544486 255134
rect 544570 254898 544806 255134
rect 563930 255218 564166 255454
rect 564250 255218 564486 255454
rect 564570 255218 564806 255454
rect 563930 254898 564166 255134
rect 564250 254898 564486 255134
rect 564570 254898 564806 255134
rect 313930 223718 314166 223954
rect 314250 223718 314486 223954
rect 314570 223718 314806 223954
rect 313930 223398 314166 223634
rect 314250 223398 314486 223634
rect 314570 223398 314806 223634
rect 333930 223718 334166 223954
rect 334250 223718 334486 223954
rect 334570 223718 334806 223954
rect 333930 223398 334166 223634
rect 334250 223398 334486 223634
rect 334570 223398 334806 223634
rect 353930 223718 354166 223954
rect 354250 223718 354486 223954
rect 354570 223718 354806 223954
rect 353930 223398 354166 223634
rect 354250 223398 354486 223634
rect 354570 223398 354806 223634
rect 373930 223718 374166 223954
rect 374250 223718 374486 223954
rect 374570 223718 374806 223954
rect 373930 223398 374166 223634
rect 374250 223398 374486 223634
rect 374570 223398 374806 223634
rect 393930 223718 394166 223954
rect 394250 223718 394486 223954
rect 394570 223718 394806 223954
rect 393930 223398 394166 223634
rect 394250 223398 394486 223634
rect 394570 223398 394806 223634
rect 413930 223718 414166 223954
rect 414250 223718 414486 223954
rect 414570 223718 414806 223954
rect 413930 223398 414166 223634
rect 414250 223398 414486 223634
rect 414570 223398 414806 223634
rect 433930 223718 434166 223954
rect 434250 223718 434486 223954
rect 434570 223718 434806 223954
rect 433930 223398 434166 223634
rect 434250 223398 434486 223634
rect 434570 223398 434806 223634
rect 453930 223718 454166 223954
rect 454250 223718 454486 223954
rect 454570 223718 454806 223954
rect 453930 223398 454166 223634
rect 454250 223398 454486 223634
rect 454570 223398 454806 223634
rect 473930 223718 474166 223954
rect 474250 223718 474486 223954
rect 474570 223718 474806 223954
rect 473930 223398 474166 223634
rect 474250 223398 474486 223634
rect 474570 223398 474806 223634
rect 493930 223718 494166 223954
rect 494250 223718 494486 223954
rect 494570 223718 494806 223954
rect 493930 223398 494166 223634
rect 494250 223398 494486 223634
rect 494570 223398 494806 223634
rect 513930 223718 514166 223954
rect 514250 223718 514486 223954
rect 514570 223718 514806 223954
rect 513930 223398 514166 223634
rect 514250 223398 514486 223634
rect 514570 223398 514806 223634
rect 533930 223718 534166 223954
rect 534250 223718 534486 223954
rect 534570 223718 534806 223954
rect 533930 223398 534166 223634
rect 534250 223398 534486 223634
rect 534570 223398 534806 223634
rect 553930 223718 554166 223954
rect 554250 223718 554486 223954
rect 554570 223718 554806 223954
rect 553930 223398 554166 223634
rect 554250 223398 554486 223634
rect 554570 223398 554806 223634
rect 303930 219218 304166 219454
rect 304250 219218 304486 219454
rect 304570 219218 304806 219454
rect 303930 218898 304166 219134
rect 304250 218898 304486 219134
rect 304570 218898 304806 219134
rect 323930 219218 324166 219454
rect 324250 219218 324486 219454
rect 324570 219218 324806 219454
rect 323930 218898 324166 219134
rect 324250 218898 324486 219134
rect 324570 218898 324806 219134
rect 343930 219218 344166 219454
rect 344250 219218 344486 219454
rect 344570 219218 344806 219454
rect 343930 218898 344166 219134
rect 344250 218898 344486 219134
rect 344570 218898 344806 219134
rect 363930 219218 364166 219454
rect 364250 219218 364486 219454
rect 364570 219218 364806 219454
rect 363930 218898 364166 219134
rect 364250 218898 364486 219134
rect 364570 218898 364806 219134
rect 383930 219218 384166 219454
rect 384250 219218 384486 219454
rect 384570 219218 384806 219454
rect 383930 218898 384166 219134
rect 384250 218898 384486 219134
rect 384570 218898 384806 219134
rect 403930 219218 404166 219454
rect 404250 219218 404486 219454
rect 404570 219218 404806 219454
rect 403930 218898 404166 219134
rect 404250 218898 404486 219134
rect 404570 218898 404806 219134
rect 423930 219218 424166 219454
rect 424250 219218 424486 219454
rect 424570 219218 424806 219454
rect 423930 218898 424166 219134
rect 424250 218898 424486 219134
rect 424570 218898 424806 219134
rect 443930 219218 444166 219454
rect 444250 219218 444486 219454
rect 444570 219218 444806 219454
rect 443930 218898 444166 219134
rect 444250 218898 444486 219134
rect 444570 218898 444806 219134
rect 463930 219218 464166 219454
rect 464250 219218 464486 219454
rect 464570 219218 464806 219454
rect 463930 218898 464166 219134
rect 464250 218898 464486 219134
rect 464570 218898 464806 219134
rect 483930 219218 484166 219454
rect 484250 219218 484486 219454
rect 484570 219218 484806 219454
rect 483930 218898 484166 219134
rect 484250 218898 484486 219134
rect 484570 218898 484806 219134
rect 503930 219218 504166 219454
rect 504250 219218 504486 219454
rect 504570 219218 504806 219454
rect 503930 218898 504166 219134
rect 504250 218898 504486 219134
rect 504570 218898 504806 219134
rect 523930 219218 524166 219454
rect 524250 219218 524486 219454
rect 524570 219218 524806 219454
rect 523930 218898 524166 219134
rect 524250 218898 524486 219134
rect 524570 218898 524806 219134
rect 543930 219218 544166 219454
rect 544250 219218 544486 219454
rect 544570 219218 544806 219454
rect 543930 218898 544166 219134
rect 544250 218898 544486 219134
rect 544570 218898 544806 219134
rect 563930 219218 564166 219454
rect 564250 219218 564486 219454
rect 564570 219218 564806 219454
rect 563930 218898 564166 219134
rect 564250 218898 564486 219134
rect 564570 218898 564806 219134
rect 303930 183218 304166 183454
rect 304250 183218 304486 183454
rect 304570 183218 304806 183454
rect 303930 182898 304166 183134
rect 304250 182898 304486 183134
rect 304570 182898 304806 183134
rect 323930 183218 324166 183454
rect 324250 183218 324486 183454
rect 324570 183218 324806 183454
rect 323930 182898 324166 183134
rect 324250 182898 324486 183134
rect 324570 182898 324806 183134
rect 343930 183218 344166 183454
rect 344250 183218 344486 183454
rect 344570 183218 344806 183454
rect 343930 182898 344166 183134
rect 344250 182898 344486 183134
rect 344570 182898 344806 183134
rect 363930 183218 364166 183454
rect 364250 183218 364486 183454
rect 364570 183218 364806 183454
rect 363930 182898 364166 183134
rect 364250 182898 364486 183134
rect 364570 182898 364806 183134
rect 383930 183218 384166 183454
rect 384250 183218 384486 183454
rect 384570 183218 384806 183454
rect 383930 182898 384166 183134
rect 384250 182898 384486 183134
rect 384570 182898 384806 183134
rect 403930 183218 404166 183454
rect 404250 183218 404486 183454
rect 404570 183218 404806 183454
rect 403930 182898 404166 183134
rect 404250 182898 404486 183134
rect 404570 182898 404806 183134
rect 423930 183218 424166 183454
rect 424250 183218 424486 183454
rect 424570 183218 424806 183454
rect 423930 182898 424166 183134
rect 424250 182898 424486 183134
rect 424570 182898 424806 183134
rect 443930 183218 444166 183454
rect 444250 183218 444486 183454
rect 444570 183218 444806 183454
rect 443930 182898 444166 183134
rect 444250 182898 444486 183134
rect 444570 182898 444806 183134
rect 463930 183218 464166 183454
rect 464250 183218 464486 183454
rect 464570 183218 464806 183454
rect 463930 182898 464166 183134
rect 464250 182898 464486 183134
rect 464570 182898 464806 183134
rect 483930 183218 484166 183454
rect 484250 183218 484486 183454
rect 484570 183218 484806 183454
rect 483930 182898 484166 183134
rect 484250 182898 484486 183134
rect 484570 182898 484806 183134
rect 503930 183218 504166 183454
rect 504250 183218 504486 183454
rect 504570 183218 504806 183454
rect 503930 182898 504166 183134
rect 504250 182898 504486 183134
rect 504570 182898 504806 183134
rect 523930 183218 524166 183454
rect 524250 183218 524486 183454
rect 524570 183218 524806 183454
rect 523930 182898 524166 183134
rect 524250 182898 524486 183134
rect 524570 182898 524806 183134
rect 543930 183218 544166 183454
rect 544250 183218 544486 183454
rect 544570 183218 544806 183454
rect 543930 182898 544166 183134
rect 544250 182898 544486 183134
rect 544570 182898 544806 183134
rect 563930 183218 564166 183454
rect 564250 183218 564486 183454
rect 564570 183218 564806 183454
rect 563930 182898 564166 183134
rect 564250 182898 564486 183134
rect 564570 182898 564806 183134
rect 313930 151718 314166 151954
rect 314250 151718 314486 151954
rect 314570 151718 314806 151954
rect 313930 151398 314166 151634
rect 314250 151398 314486 151634
rect 314570 151398 314806 151634
rect 333930 151718 334166 151954
rect 334250 151718 334486 151954
rect 334570 151718 334806 151954
rect 333930 151398 334166 151634
rect 334250 151398 334486 151634
rect 334570 151398 334806 151634
rect 353930 151718 354166 151954
rect 354250 151718 354486 151954
rect 354570 151718 354806 151954
rect 353930 151398 354166 151634
rect 354250 151398 354486 151634
rect 354570 151398 354806 151634
rect 373930 151718 374166 151954
rect 374250 151718 374486 151954
rect 374570 151718 374806 151954
rect 373930 151398 374166 151634
rect 374250 151398 374486 151634
rect 374570 151398 374806 151634
rect 393930 151718 394166 151954
rect 394250 151718 394486 151954
rect 394570 151718 394806 151954
rect 393930 151398 394166 151634
rect 394250 151398 394486 151634
rect 394570 151398 394806 151634
rect 413930 151718 414166 151954
rect 414250 151718 414486 151954
rect 414570 151718 414806 151954
rect 413930 151398 414166 151634
rect 414250 151398 414486 151634
rect 414570 151398 414806 151634
rect 433930 151718 434166 151954
rect 434250 151718 434486 151954
rect 434570 151718 434806 151954
rect 433930 151398 434166 151634
rect 434250 151398 434486 151634
rect 434570 151398 434806 151634
rect 453930 151718 454166 151954
rect 454250 151718 454486 151954
rect 454570 151718 454806 151954
rect 453930 151398 454166 151634
rect 454250 151398 454486 151634
rect 454570 151398 454806 151634
rect 473930 151718 474166 151954
rect 474250 151718 474486 151954
rect 474570 151718 474806 151954
rect 473930 151398 474166 151634
rect 474250 151398 474486 151634
rect 474570 151398 474806 151634
rect 493930 151718 494166 151954
rect 494250 151718 494486 151954
rect 494570 151718 494806 151954
rect 493930 151398 494166 151634
rect 494250 151398 494486 151634
rect 494570 151398 494806 151634
rect 513930 151718 514166 151954
rect 514250 151718 514486 151954
rect 514570 151718 514806 151954
rect 513930 151398 514166 151634
rect 514250 151398 514486 151634
rect 514570 151398 514806 151634
rect 533930 151718 534166 151954
rect 534250 151718 534486 151954
rect 534570 151718 534806 151954
rect 533930 151398 534166 151634
rect 534250 151398 534486 151634
rect 534570 151398 534806 151634
rect 553930 151718 554166 151954
rect 554250 151718 554486 151954
rect 554570 151718 554806 151954
rect 553930 151398 554166 151634
rect 554250 151398 554486 151634
rect 554570 151398 554806 151634
rect 303930 147218 304166 147454
rect 304250 147218 304486 147454
rect 304570 147218 304806 147454
rect 303930 146898 304166 147134
rect 304250 146898 304486 147134
rect 304570 146898 304806 147134
rect 323930 147218 324166 147454
rect 324250 147218 324486 147454
rect 324570 147218 324806 147454
rect 323930 146898 324166 147134
rect 324250 146898 324486 147134
rect 324570 146898 324806 147134
rect 343930 147218 344166 147454
rect 344250 147218 344486 147454
rect 344570 147218 344806 147454
rect 343930 146898 344166 147134
rect 344250 146898 344486 147134
rect 344570 146898 344806 147134
rect 363930 147218 364166 147454
rect 364250 147218 364486 147454
rect 364570 147218 364806 147454
rect 363930 146898 364166 147134
rect 364250 146898 364486 147134
rect 364570 146898 364806 147134
rect 383930 147218 384166 147454
rect 384250 147218 384486 147454
rect 384570 147218 384806 147454
rect 383930 146898 384166 147134
rect 384250 146898 384486 147134
rect 384570 146898 384806 147134
rect 403930 147218 404166 147454
rect 404250 147218 404486 147454
rect 404570 147218 404806 147454
rect 403930 146898 404166 147134
rect 404250 146898 404486 147134
rect 404570 146898 404806 147134
rect 423930 147218 424166 147454
rect 424250 147218 424486 147454
rect 424570 147218 424806 147454
rect 423930 146898 424166 147134
rect 424250 146898 424486 147134
rect 424570 146898 424806 147134
rect 443930 147218 444166 147454
rect 444250 147218 444486 147454
rect 444570 147218 444806 147454
rect 443930 146898 444166 147134
rect 444250 146898 444486 147134
rect 444570 146898 444806 147134
rect 463930 147218 464166 147454
rect 464250 147218 464486 147454
rect 464570 147218 464806 147454
rect 463930 146898 464166 147134
rect 464250 146898 464486 147134
rect 464570 146898 464806 147134
rect 483930 147218 484166 147454
rect 484250 147218 484486 147454
rect 484570 147218 484806 147454
rect 483930 146898 484166 147134
rect 484250 146898 484486 147134
rect 484570 146898 484806 147134
rect 503930 147218 504166 147454
rect 504250 147218 504486 147454
rect 504570 147218 504806 147454
rect 503930 146898 504166 147134
rect 504250 146898 504486 147134
rect 504570 146898 504806 147134
rect 523930 147218 524166 147454
rect 524250 147218 524486 147454
rect 524570 147218 524806 147454
rect 523930 146898 524166 147134
rect 524250 146898 524486 147134
rect 524570 146898 524806 147134
rect 543930 147218 544166 147454
rect 544250 147218 544486 147454
rect 544570 147218 544806 147454
rect 543930 146898 544166 147134
rect 544250 146898 544486 147134
rect 544570 146898 544806 147134
rect 563930 147218 564166 147454
rect 564250 147218 564486 147454
rect 564570 147218 564806 147454
rect 563930 146898 564166 147134
rect 564250 146898 564486 147134
rect 564570 146898 564806 147134
rect 313930 115718 314166 115954
rect 314250 115718 314486 115954
rect 314570 115718 314806 115954
rect 313930 115398 314166 115634
rect 314250 115398 314486 115634
rect 314570 115398 314806 115634
rect 333930 115718 334166 115954
rect 334250 115718 334486 115954
rect 334570 115718 334806 115954
rect 333930 115398 334166 115634
rect 334250 115398 334486 115634
rect 334570 115398 334806 115634
rect 353930 115718 354166 115954
rect 354250 115718 354486 115954
rect 354570 115718 354806 115954
rect 353930 115398 354166 115634
rect 354250 115398 354486 115634
rect 354570 115398 354806 115634
rect 373930 115718 374166 115954
rect 374250 115718 374486 115954
rect 374570 115718 374806 115954
rect 373930 115398 374166 115634
rect 374250 115398 374486 115634
rect 374570 115398 374806 115634
rect 393930 115718 394166 115954
rect 394250 115718 394486 115954
rect 394570 115718 394806 115954
rect 393930 115398 394166 115634
rect 394250 115398 394486 115634
rect 394570 115398 394806 115634
rect 413930 115718 414166 115954
rect 414250 115718 414486 115954
rect 414570 115718 414806 115954
rect 413930 115398 414166 115634
rect 414250 115398 414486 115634
rect 414570 115398 414806 115634
rect 433930 115718 434166 115954
rect 434250 115718 434486 115954
rect 434570 115718 434806 115954
rect 433930 115398 434166 115634
rect 434250 115398 434486 115634
rect 434570 115398 434806 115634
rect 453930 115718 454166 115954
rect 454250 115718 454486 115954
rect 454570 115718 454806 115954
rect 453930 115398 454166 115634
rect 454250 115398 454486 115634
rect 454570 115398 454806 115634
rect 473930 115718 474166 115954
rect 474250 115718 474486 115954
rect 474570 115718 474806 115954
rect 473930 115398 474166 115634
rect 474250 115398 474486 115634
rect 474570 115398 474806 115634
rect 493930 115718 494166 115954
rect 494250 115718 494486 115954
rect 494570 115718 494806 115954
rect 493930 115398 494166 115634
rect 494250 115398 494486 115634
rect 494570 115398 494806 115634
rect 513930 115718 514166 115954
rect 514250 115718 514486 115954
rect 514570 115718 514806 115954
rect 513930 115398 514166 115634
rect 514250 115398 514486 115634
rect 514570 115398 514806 115634
rect 533930 115718 534166 115954
rect 534250 115718 534486 115954
rect 534570 115718 534806 115954
rect 533930 115398 534166 115634
rect 534250 115398 534486 115634
rect 534570 115398 534806 115634
rect 553930 115718 554166 115954
rect 554250 115718 554486 115954
rect 554570 115718 554806 115954
rect 553930 115398 554166 115634
rect 554250 115398 554486 115634
rect 554570 115398 554806 115634
rect 303930 111218 304166 111454
rect 304250 111218 304486 111454
rect 304570 111218 304806 111454
rect 303930 110898 304166 111134
rect 304250 110898 304486 111134
rect 304570 110898 304806 111134
rect 323930 111218 324166 111454
rect 324250 111218 324486 111454
rect 324570 111218 324806 111454
rect 323930 110898 324166 111134
rect 324250 110898 324486 111134
rect 324570 110898 324806 111134
rect 343930 111218 344166 111454
rect 344250 111218 344486 111454
rect 344570 111218 344806 111454
rect 343930 110898 344166 111134
rect 344250 110898 344486 111134
rect 344570 110898 344806 111134
rect 363930 111218 364166 111454
rect 364250 111218 364486 111454
rect 364570 111218 364806 111454
rect 363930 110898 364166 111134
rect 364250 110898 364486 111134
rect 364570 110898 364806 111134
rect 383930 111218 384166 111454
rect 384250 111218 384486 111454
rect 384570 111218 384806 111454
rect 383930 110898 384166 111134
rect 384250 110898 384486 111134
rect 384570 110898 384806 111134
rect 403930 111218 404166 111454
rect 404250 111218 404486 111454
rect 404570 111218 404806 111454
rect 403930 110898 404166 111134
rect 404250 110898 404486 111134
rect 404570 110898 404806 111134
rect 423930 111218 424166 111454
rect 424250 111218 424486 111454
rect 424570 111218 424806 111454
rect 423930 110898 424166 111134
rect 424250 110898 424486 111134
rect 424570 110898 424806 111134
rect 443930 111218 444166 111454
rect 444250 111218 444486 111454
rect 444570 111218 444806 111454
rect 443930 110898 444166 111134
rect 444250 110898 444486 111134
rect 444570 110898 444806 111134
rect 463930 111218 464166 111454
rect 464250 111218 464486 111454
rect 464570 111218 464806 111454
rect 463930 110898 464166 111134
rect 464250 110898 464486 111134
rect 464570 110898 464806 111134
rect 483930 111218 484166 111454
rect 484250 111218 484486 111454
rect 484570 111218 484806 111454
rect 483930 110898 484166 111134
rect 484250 110898 484486 111134
rect 484570 110898 484806 111134
rect 503930 111218 504166 111454
rect 504250 111218 504486 111454
rect 504570 111218 504806 111454
rect 503930 110898 504166 111134
rect 504250 110898 504486 111134
rect 504570 110898 504806 111134
rect 523930 111218 524166 111454
rect 524250 111218 524486 111454
rect 524570 111218 524806 111454
rect 523930 110898 524166 111134
rect 524250 110898 524486 111134
rect 524570 110898 524806 111134
rect 543930 111218 544166 111454
rect 544250 111218 544486 111454
rect 544570 111218 544806 111454
rect 543930 110898 544166 111134
rect 544250 110898 544486 111134
rect 544570 110898 544806 111134
rect 563930 111218 564166 111454
rect 564250 111218 564486 111454
rect 564570 111218 564806 111454
rect 563930 110898 564166 111134
rect 564250 110898 564486 111134
rect 564570 110898 564806 111134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 213930 43718 214166 43954
rect 214250 43718 214486 43954
rect 214570 43718 214806 43954
rect 213930 43398 214166 43634
rect 214250 43398 214486 43634
rect 214570 43398 214806 43634
rect 233930 43718 234166 43954
rect 234250 43718 234486 43954
rect 234570 43718 234806 43954
rect 233930 43398 234166 43634
rect 234250 43398 234486 43634
rect 234570 43398 234806 43634
rect 253930 43718 254166 43954
rect 254250 43718 254486 43954
rect 254570 43718 254806 43954
rect 253930 43398 254166 43634
rect 254250 43398 254486 43634
rect 254570 43398 254806 43634
rect 273930 43718 274166 43954
rect 274250 43718 274486 43954
rect 274570 43718 274806 43954
rect 273930 43398 274166 43634
rect 274250 43398 274486 43634
rect 274570 43398 274806 43634
rect 293930 43718 294166 43954
rect 294250 43718 294486 43954
rect 294570 43718 294806 43954
rect 293930 43398 294166 43634
rect 294250 43398 294486 43634
rect 294570 43398 294806 43634
rect 313930 43718 314166 43954
rect 314250 43718 314486 43954
rect 314570 43718 314806 43954
rect 313930 43398 314166 43634
rect 314250 43398 314486 43634
rect 314570 43398 314806 43634
rect 333930 43718 334166 43954
rect 334250 43718 334486 43954
rect 334570 43718 334806 43954
rect 333930 43398 334166 43634
rect 334250 43398 334486 43634
rect 334570 43398 334806 43634
rect 353930 43718 354166 43954
rect 354250 43718 354486 43954
rect 354570 43718 354806 43954
rect 353930 43398 354166 43634
rect 354250 43398 354486 43634
rect 354570 43398 354806 43634
rect 373930 43718 374166 43954
rect 374250 43718 374486 43954
rect 374570 43718 374806 43954
rect 373930 43398 374166 43634
rect 374250 43398 374486 43634
rect 374570 43398 374806 43634
rect 393930 43718 394166 43954
rect 394250 43718 394486 43954
rect 394570 43718 394806 43954
rect 393930 43398 394166 43634
rect 394250 43398 394486 43634
rect 394570 43398 394806 43634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 203930 39218 204166 39454
rect 204250 39218 204486 39454
rect 204570 39218 204806 39454
rect 203930 38898 204166 39134
rect 204250 38898 204486 39134
rect 204570 38898 204806 39134
rect 223930 39218 224166 39454
rect 224250 39218 224486 39454
rect 224570 39218 224806 39454
rect 223930 38898 224166 39134
rect 224250 38898 224486 39134
rect 224570 38898 224806 39134
rect 243930 39218 244166 39454
rect 244250 39218 244486 39454
rect 244570 39218 244806 39454
rect 243930 38898 244166 39134
rect 244250 38898 244486 39134
rect 244570 38898 244806 39134
rect 263930 39218 264166 39454
rect 264250 39218 264486 39454
rect 264570 39218 264806 39454
rect 263930 38898 264166 39134
rect 264250 38898 264486 39134
rect 264570 38898 264806 39134
rect 283930 39218 284166 39454
rect 284250 39218 284486 39454
rect 284570 39218 284806 39454
rect 283930 38898 284166 39134
rect 284250 38898 284486 39134
rect 284570 38898 284806 39134
rect 303930 39218 304166 39454
rect 304250 39218 304486 39454
rect 304570 39218 304806 39454
rect 303930 38898 304166 39134
rect 304250 38898 304486 39134
rect 304570 38898 304806 39134
rect 323930 39218 324166 39454
rect 324250 39218 324486 39454
rect 324570 39218 324806 39454
rect 323930 38898 324166 39134
rect 324250 38898 324486 39134
rect 324570 38898 324806 39134
rect 343930 39218 344166 39454
rect 344250 39218 344486 39454
rect 344570 39218 344806 39454
rect 343930 38898 344166 39134
rect 344250 38898 344486 39134
rect 344570 38898 344806 39134
rect 363930 39218 364166 39454
rect 364250 39218 364486 39454
rect 364570 39218 364806 39454
rect 363930 38898 364166 39134
rect 364250 38898 364486 39134
rect 364570 38898 364806 39134
rect 383930 39218 384166 39454
rect 384250 39218 384486 39454
rect 384570 39218 384806 39454
rect 383930 38898 384166 39134
rect 384250 38898 384486 39134
rect 384570 38898 384806 39134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 33930 691954
rect 34166 691718 34250 691954
rect 34486 691718 34570 691954
rect 34806 691718 53930 691954
rect 54166 691718 54250 691954
rect 54486 691718 54570 691954
rect 54806 691718 73930 691954
rect 74166 691718 74250 691954
rect 74486 691718 74570 691954
rect 74806 691718 93930 691954
rect 94166 691718 94250 691954
rect 94486 691718 94570 691954
rect 94806 691718 113930 691954
rect 114166 691718 114250 691954
rect 114486 691718 114570 691954
rect 114806 691718 133930 691954
rect 134166 691718 134250 691954
rect 134486 691718 134570 691954
rect 134806 691718 153930 691954
rect 154166 691718 154250 691954
rect 154486 691718 154570 691954
rect 154806 691718 173930 691954
rect 174166 691718 174250 691954
rect 174486 691718 174570 691954
rect 174806 691718 193930 691954
rect 194166 691718 194250 691954
rect 194486 691718 194570 691954
rect 194806 691718 213930 691954
rect 214166 691718 214250 691954
rect 214486 691718 214570 691954
rect 214806 691718 233930 691954
rect 234166 691718 234250 691954
rect 234486 691718 234570 691954
rect 234806 691718 253930 691954
rect 254166 691718 254250 691954
rect 254486 691718 254570 691954
rect 254806 691718 273930 691954
rect 274166 691718 274250 691954
rect 274486 691718 274570 691954
rect 274806 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 313930 691954
rect 314166 691718 314250 691954
rect 314486 691718 314570 691954
rect 314806 691718 333930 691954
rect 334166 691718 334250 691954
rect 334486 691718 334570 691954
rect 334806 691718 353930 691954
rect 354166 691718 354250 691954
rect 354486 691718 354570 691954
rect 354806 691718 373930 691954
rect 374166 691718 374250 691954
rect 374486 691718 374570 691954
rect 374806 691718 393930 691954
rect 394166 691718 394250 691954
rect 394486 691718 394570 691954
rect 394806 691718 413930 691954
rect 414166 691718 414250 691954
rect 414486 691718 414570 691954
rect 414806 691718 433930 691954
rect 434166 691718 434250 691954
rect 434486 691718 434570 691954
rect 434806 691718 453930 691954
rect 454166 691718 454250 691954
rect 454486 691718 454570 691954
rect 454806 691718 473930 691954
rect 474166 691718 474250 691954
rect 474486 691718 474570 691954
rect 474806 691718 493930 691954
rect 494166 691718 494250 691954
rect 494486 691718 494570 691954
rect 494806 691718 513930 691954
rect 514166 691718 514250 691954
rect 514486 691718 514570 691954
rect 514806 691718 533930 691954
rect 534166 691718 534250 691954
rect 534486 691718 534570 691954
rect 534806 691718 553930 691954
rect 554166 691718 554250 691954
rect 554486 691718 554570 691954
rect 554806 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 33930 691634
rect 34166 691398 34250 691634
rect 34486 691398 34570 691634
rect 34806 691398 53930 691634
rect 54166 691398 54250 691634
rect 54486 691398 54570 691634
rect 54806 691398 73930 691634
rect 74166 691398 74250 691634
rect 74486 691398 74570 691634
rect 74806 691398 93930 691634
rect 94166 691398 94250 691634
rect 94486 691398 94570 691634
rect 94806 691398 113930 691634
rect 114166 691398 114250 691634
rect 114486 691398 114570 691634
rect 114806 691398 133930 691634
rect 134166 691398 134250 691634
rect 134486 691398 134570 691634
rect 134806 691398 153930 691634
rect 154166 691398 154250 691634
rect 154486 691398 154570 691634
rect 154806 691398 173930 691634
rect 174166 691398 174250 691634
rect 174486 691398 174570 691634
rect 174806 691398 193930 691634
rect 194166 691398 194250 691634
rect 194486 691398 194570 691634
rect 194806 691398 213930 691634
rect 214166 691398 214250 691634
rect 214486 691398 214570 691634
rect 214806 691398 233930 691634
rect 234166 691398 234250 691634
rect 234486 691398 234570 691634
rect 234806 691398 253930 691634
rect 254166 691398 254250 691634
rect 254486 691398 254570 691634
rect 254806 691398 273930 691634
rect 274166 691398 274250 691634
rect 274486 691398 274570 691634
rect 274806 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 313930 691634
rect 314166 691398 314250 691634
rect 314486 691398 314570 691634
rect 314806 691398 333930 691634
rect 334166 691398 334250 691634
rect 334486 691398 334570 691634
rect 334806 691398 353930 691634
rect 354166 691398 354250 691634
rect 354486 691398 354570 691634
rect 354806 691398 373930 691634
rect 374166 691398 374250 691634
rect 374486 691398 374570 691634
rect 374806 691398 393930 691634
rect 394166 691398 394250 691634
rect 394486 691398 394570 691634
rect 394806 691398 413930 691634
rect 414166 691398 414250 691634
rect 414486 691398 414570 691634
rect 414806 691398 433930 691634
rect 434166 691398 434250 691634
rect 434486 691398 434570 691634
rect 434806 691398 453930 691634
rect 454166 691398 454250 691634
rect 454486 691398 454570 691634
rect 454806 691398 473930 691634
rect 474166 691398 474250 691634
rect 474486 691398 474570 691634
rect 474806 691398 493930 691634
rect 494166 691398 494250 691634
rect 494486 691398 494570 691634
rect 494806 691398 513930 691634
rect 514166 691398 514250 691634
rect 514486 691398 514570 691634
rect 514806 691398 533930 691634
rect 534166 691398 534250 691634
rect 534486 691398 534570 691634
rect 534806 691398 553930 691634
rect 554166 691398 554250 691634
rect 554486 691398 554570 691634
rect 554806 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 23930 687454
rect 24166 687218 24250 687454
rect 24486 687218 24570 687454
rect 24806 687218 43930 687454
rect 44166 687218 44250 687454
rect 44486 687218 44570 687454
rect 44806 687218 63930 687454
rect 64166 687218 64250 687454
rect 64486 687218 64570 687454
rect 64806 687218 83930 687454
rect 84166 687218 84250 687454
rect 84486 687218 84570 687454
rect 84806 687218 103930 687454
rect 104166 687218 104250 687454
rect 104486 687218 104570 687454
rect 104806 687218 123930 687454
rect 124166 687218 124250 687454
rect 124486 687218 124570 687454
rect 124806 687218 143930 687454
rect 144166 687218 144250 687454
rect 144486 687218 144570 687454
rect 144806 687218 163930 687454
rect 164166 687218 164250 687454
rect 164486 687218 164570 687454
rect 164806 687218 183930 687454
rect 184166 687218 184250 687454
rect 184486 687218 184570 687454
rect 184806 687218 203930 687454
rect 204166 687218 204250 687454
rect 204486 687218 204570 687454
rect 204806 687218 223930 687454
rect 224166 687218 224250 687454
rect 224486 687218 224570 687454
rect 224806 687218 243930 687454
rect 244166 687218 244250 687454
rect 244486 687218 244570 687454
rect 244806 687218 263930 687454
rect 264166 687218 264250 687454
rect 264486 687218 264570 687454
rect 264806 687218 283930 687454
rect 284166 687218 284250 687454
rect 284486 687218 284570 687454
rect 284806 687218 303930 687454
rect 304166 687218 304250 687454
rect 304486 687218 304570 687454
rect 304806 687218 323930 687454
rect 324166 687218 324250 687454
rect 324486 687218 324570 687454
rect 324806 687218 343930 687454
rect 344166 687218 344250 687454
rect 344486 687218 344570 687454
rect 344806 687218 363930 687454
rect 364166 687218 364250 687454
rect 364486 687218 364570 687454
rect 364806 687218 383930 687454
rect 384166 687218 384250 687454
rect 384486 687218 384570 687454
rect 384806 687218 403930 687454
rect 404166 687218 404250 687454
rect 404486 687218 404570 687454
rect 404806 687218 423930 687454
rect 424166 687218 424250 687454
rect 424486 687218 424570 687454
rect 424806 687218 443930 687454
rect 444166 687218 444250 687454
rect 444486 687218 444570 687454
rect 444806 687218 463930 687454
rect 464166 687218 464250 687454
rect 464486 687218 464570 687454
rect 464806 687218 483930 687454
rect 484166 687218 484250 687454
rect 484486 687218 484570 687454
rect 484806 687218 503930 687454
rect 504166 687218 504250 687454
rect 504486 687218 504570 687454
rect 504806 687218 523930 687454
rect 524166 687218 524250 687454
rect 524486 687218 524570 687454
rect 524806 687218 543930 687454
rect 544166 687218 544250 687454
rect 544486 687218 544570 687454
rect 544806 687218 563930 687454
rect 564166 687218 564250 687454
rect 564486 687218 564570 687454
rect 564806 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 23930 687134
rect 24166 686898 24250 687134
rect 24486 686898 24570 687134
rect 24806 686898 43930 687134
rect 44166 686898 44250 687134
rect 44486 686898 44570 687134
rect 44806 686898 63930 687134
rect 64166 686898 64250 687134
rect 64486 686898 64570 687134
rect 64806 686898 83930 687134
rect 84166 686898 84250 687134
rect 84486 686898 84570 687134
rect 84806 686898 103930 687134
rect 104166 686898 104250 687134
rect 104486 686898 104570 687134
rect 104806 686898 123930 687134
rect 124166 686898 124250 687134
rect 124486 686898 124570 687134
rect 124806 686898 143930 687134
rect 144166 686898 144250 687134
rect 144486 686898 144570 687134
rect 144806 686898 163930 687134
rect 164166 686898 164250 687134
rect 164486 686898 164570 687134
rect 164806 686898 183930 687134
rect 184166 686898 184250 687134
rect 184486 686898 184570 687134
rect 184806 686898 203930 687134
rect 204166 686898 204250 687134
rect 204486 686898 204570 687134
rect 204806 686898 223930 687134
rect 224166 686898 224250 687134
rect 224486 686898 224570 687134
rect 224806 686898 243930 687134
rect 244166 686898 244250 687134
rect 244486 686898 244570 687134
rect 244806 686898 263930 687134
rect 264166 686898 264250 687134
rect 264486 686898 264570 687134
rect 264806 686898 283930 687134
rect 284166 686898 284250 687134
rect 284486 686898 284570 687134
rect 284806 686898 303930 687134
rect 304166 686898 304250 687134
rect 304486 686898 304570 687134
rect 304806 686898 323930 687134
rect 324166 686898 324250 687134
rect 324486 686898 324570 687134
rect 324806 686898 343930 687134
rect 344166 686898 344250 687134
rect 344486 686898 344570 687134
rect 344806 686898 363930 687134
rect 364166 686898 364250 687134
rect 364486 686898 364570 687134
rect 364806 686898 383930 687134
rect 384166 686898 384250 687134
rect 384486 686898 384570 687134
rect 384806 686898 403930 687134
rect 404166 686898 404250 687134
rect 404486 686898 404570 687134
rect 404806 686898 423930 687134
rect 424166 686898 424250 687134
rect 424486 686898 424570 687134
rect 424806 686898 443930 687134
rect 444166 686898 444250 687134
rect 444486 686898 444570 687134
rect 444806 686898 463930 687134
rect 464166 686898 464250 687134
rect 464486 686898 464570 687134
rect 464806 686898 483930 687134
rect 484166 686898 484250 687134
rect 484486 686898 484570 687134
rect 484806 686898 503930 687134
rect 504166 686898 504250 687134
rect 504486 686898 504570 687134
rect 504806 686898 523930 687134
rect 524166 686898 524250 687134
rect 524486 686898 524570 687134
rect 524806 686898 543930 687134
rect 544166 686898 544250 687134
rect 544486 686898 544570 687134
rect 544806 686898 563930 687134
rect 564166 686898 564250 687134
rect 564486 686898 564570 687134
rect 564806 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 33930 655954
rect 34166 655718 34250 655954
rect 34486 655718 34570 655954
rect 34806 655718 53930 655954
rect 54166 655718 54250 655954
rect 54486 655718 54570 655954
rect 54806 655718 73930 655954
rect 74166 655718 74250 655954
rect 74486 655718 74570 655954
rect 74806 655718 93930 655954
rect 94166 655718 94250 655954
rect 94486 655718 94570 655954
rect 94806 655718 113930 655954
rect 114166 655718 114250 655954
rect 114486 655718 114570 655954
rect 114806 655718 133930 655954
rect 134166 655718 134250 655954
rect 134486 655718 134570 655954
rect 134806 655718 153930 655954
rect 154166 655718 154250 655954
rect 154486 655718 154570 655954
rect 154806 655718 173930 655954
rect 174166 655718 174250 655954
rect 174486 655718 174570 655954
rect 174806 655718 193930 655954
rect 194166 655718 194250 655954
rect 194486 655718 194570 655954
rect 194806 655718 213930 655954
rect 214166 655718 214250 655954
rect 214486 655718 214570 655954
rect 214806 655718 233930 655954
rect 234166 655718 234250 655954
rect 234486 655718 234570 655954
rect 234806 655718 253930 655954
rect 254166 655718 254250 655954
rect 254486 655718 254570 655954
rect 254806 655718 273930 655954
rect 274166 655718 274250 655954
rect 274486 655718 274570 655954
rect 274806 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 313930 655954
rect 314166 655718 314250 655954
rect 314486 655718 314570 655954
rect 314806 655718 333930 655954
rect 334166 655718 334250 655954
rect 334486 655718 334570 655954
rect 334806 655718 353930 655954
rect 354166 655718 354250 655954
rect 354486 655718 354570 655954
rect 354806 655718 373930 655954
rect 374166 655718 374250 655954
rect 374486 655718 374570 655954
rect 374806 655718 393930 655954
rect 394166 655718 394250 655954
rect 394486 655718 394570 655954
rect 394806 655718 413930 655954
rect 414166 655718 414250 655954
rect 414486 655718 414570 655954
rect 414806 655718 433930 655954
rect 434166 655718 434250 655954
rect 434486 655718 434570 655954
rect 434806 655718 453930 655954
rect 454166 655718 454250 655954
rect 454486 655718 454570 655954
rect 454806 655718 473930 655954
rect 474166 655718 474250 655954
rect 474486 655718 474570 655954
rect 474806 655718 493930 655954
rect 494166 655718 494250 655954
rect 494486 655718 494570 655954
rect 494806 655718 513930 655954
rect 514166 655718 514250 655954
rect 514486 655718 514570 655954
rect 514806 655718 533930 655954
rect 534166 655718 534250 655954
rect 534486 655718 534570 655954
rect 534806 655718 553930 655954
rect 554166 655718 554250 655954
rect 554486 655718 554570 655954
rect 554806 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 33930 655634
rect 34166 655398 34250 655634
rect 34486 655398 34570 655634
rect 34806 655398 53930 655634
rect 54166 655398 54250 655634
rect 54486 655398 54570 655634
rect 54806 655398 73930 655634
rect 74166 655398 74250 655634
rect 74486 655398 74570 655634
rect 74806 655398 93930 655634
rect 94166 655398 94250 655634
rect 94486 655398 94570 655634
rect 94806 655398 113930 655634
rect 114166 655398 114250 655634
rect 114486 655398 114570 655634
rect 114806 655398 133930 655634
rect 134166 655398 134250 655634
rect 134486 655398 134570 655634
rect 134806 655398 153930 655634
rect 154166 655398 154250 655634
rect 154486 655398 154570 655634
rect 154806 655398 173930 655634
rect 174166 655398 174250 655634
rect 174486 655398 174570 655634
rect 174806 655398 193930 655634
rect 194166 655398 194250 655634
rect 194486 655398 194570 655634
rect 194806 655398 213930 655634
rect 214166 655398 214250 655634
rect 214486 655398 214570 655634
rect 214806 655398 233930 655634
rect 234166 655398 234250 655634
rect 234486 655398 234570 655634
rect 234806 655398 253930 655634
rect 254166 655398 254250 655634
rect 254486 655398 254570 655634
rect 254806 655398 273930 655634
rect 274166 655398 274250 655634
rect 274486 655398 274570 655634
rect 274806 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 313930 655634
rect 314166 655398 314250 655634
rect 314486 655398 314570 655634
rect 314806 655398 333930 655634
rect 334166 655398 334250 655634
rect 334486 655398 334570 655634
rect 334806 655398 353930 655634
rect 354166 655398 354250 655634
rect 354486 655398 354570 655634
rect 354806 655398 373930 655634
rect 374166 655398 374250 655634
rect 374486 655398 374570 655634
rect 374806 655398 393930 655634
rect 394166 655398 394250 655634
rect 394486 655398 394570 655634
rect 394806 655398 413930 655634
rect 414166 655398 414250 655634
rect 414486 655398 414570 655634
rect 414806 655398 433930 655634
rect 434166 655398 434250 655634
rect 434486 655398 434570 655634
rect 434806 655398 453930 655634
rect 454166 655398 454250 655634
rect 454486 655398 454570 655634
rect 454806 655398 473930 655634
rect 474166 655398 474250 655634
rect 474486 655398 474570 655634
rect 474806 655398 493930 655634
rect 494166 655398 494250 655634
rect 494486 655398 494570 655634
rect 494806 655398 513930 655634
rect 514166 655398 514250 655634
rect 514486 655398 514570 655634
rect 514806 655398 533930 655634
rect 534166 655398 534250 655634
rect 534486 655398 534570 655634
rect 534806 655398 553930 655634
rect 554166 655398 554250 655634
rect 554486 655398 554570 655634
rect 554806 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 23930 651454
rect 24166 651218 24250 651454
rect 24486 651218 24570 651454
rect 24806 651218 43930 651454
rect 44166 651218 44250 651454
rect 44486 651218 44570 651454
rect 44806 651218 63930 651454
rect 64166 651218 64250 651454
rect 64486 651218 64570 651454
rect 64806 651218 83930 651454
rect 84166 651218 84250 651454
rect 84486 651218 84570 651454
rect 84806 651218 103930 651454
rect 104166 651218 104250 651454
rect 104486 651218 104570 651454
rect 104806 651218 123930 651454
rect 124166 651218 124250 651454
rect 124486 651218 124570 651454
rect 124806 651218 143930 651454
rect 144166 651218 144250 651454
rect 144486 651218 144570 651454
rect 144806 651218 163930 651454
rect 164166 651218 164250 651454
rect 164486 651218 164570 651454
rect 164806 651218 183930 651454
rect 184166 651218 184250 651454
rect 184486 651218 184570 651454
rect 184806 651218 203930 651454
rect 204166 651218 204250 651454
rect 204486 651218 204570 651454
rect 204806 651218 223930 651454
rect 224166 651218 224250 651454
rect 224486 651218 224570 651454
rect 224806 651218 243930 651454
rect 244166 651218 244250 651454
rect 244486 651218 244570 651454
rect 244806 651218 263930 651454
rect 264166 651218 264250 651454
rect 264486 651218 264570 651454
rect 264806 651218 283930 651454
rect 284166 651218 284250 651454
rect 284486 651218 284570 651454
rect 284806 651218 303930 651454
rect 304166 651218 304250 651454
rect 304486 651218 304570 651454
rect 304806 651218 323930 651454
rect 324166 651218 324250 651454
rect 324486 651218 324570 651454
rect 324806 651218 343930 651454
rect 344166 651218 344250 651454
rect 344486 651218 344570 651454
rect 344806 651218 363930 651454
rect 364166 651218 364250 651454
rect 364486 651218 364570 651454
rect 364806 651218 383930 651454
rect 384166 651218 384250 651454
rect 384486 651218 384570 651454
rect 384806 651218 403930 651454
rect 404166 651218 404250 651454
rect 404486 651218 404570 651454
rect 404806 651218 423930 651454
rect 424166 651218 424250 651454
rect 424486 651218 424570 651454
rect 424806 651218 443930 651454
rect 444166 651218 444250 651454
rect 444486 651218 444570 651454
rect 444806 651218 463930 651454
rect 464166 651218 464250 651454
rect 464486 651218 464570 651454
rect 464806 651218 483930 651454
rect 484166 651218 484250 651454
rect 484486 651218 484570 651454
rect 484806 651218 503930 651454
rect 504166 651218 504250 651454
rect 504486 651218 504570 651454
rect 504806 651218 523930 651454
rect 524166 651218 524250 651454
rect 524486 651218 524570 651454
rect 524806 651218 543930 651454
rect 544166 651218 544250 651454
rect 544486 651218 544570 651454
rect 544806 651218 563930 651454
rect 564166 651218 564250 651454
rect 564486 651218 564570 651454
rect 564806 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 23930 651134
rect 24166 650898 24250 651134
rect 24486 650898 24570 651134
rect 24806 650898 43930 651134
rect 44166 650898 44250 651134
rect 44486 650898 44570 651134
rect 44806 650898 63930 651134
rect 64166 650898 64250 651134
rect 64486 650898 64570 651134
rect 64806 650898 83930 651134
rect 84166 650898 84250 651134
rect 84486 650898 84570 651134
rect 84806 650898 103930 651134
rect 104166 650898 104250 651134
rect 104486 650898 104570 651134
rect 104806 650898 123930 651134
rect 124166 650898 124250 651134
rect 124486 650898 124570 651134
rect 124806 650898 143930 651134
rect 144166 650898 144250 651134
rect 144486 650898 144570 651134
rect 144806 650898 163930 651134
rect 164166 650898 164250 651134
rect 164486 650898 164570 651134
rect 164806 650898 183930 651134
rect 184166 650898 184250 651134
rect 184486 650898 184570 651134
rect 184806 650898 203930 651134
rect 204166 650898 204250 651134
rect 204486 650898 204570 651134
rect 204806 650898 223930 651134
rect 224166 650898 224250 651134
rect 224486 650898 224570 651134
rect 224806 650898 243930 651134
rect 244166 650898 244250 651134
rect 244486 650898 244570 651134
rect 244806 650898 263930 651134
rect 264166 650898 264250 651134
rect 264486 650898 264570 651134
rect 264806 650898 283930 651134
rect 284166 650898 284250 651134
rect 284486 650898 284570 651134
rect 284806 650898 303930 651134
rect 304166 650898 304250 651134
rect 304486 650898 304570 651134
rect 304806 650898 323930 651134
rect 324166 650898 324250 651134
rect 324486 650898 324570 651134
rect 324806 650898 343930 651134
rect 344166 650898 344250 651134
rect 344486 650898 344570 651134
rect 344806 650898 363930 651134
rect 364166 650898 364250 651134
rect 364486 650898 364570 651134
rect 364806 650898 383930 651134
rect 384166 650898 384250 651134
rect 384486 650898 384570 651134
rect 384806 650898 403930 651134
rect 404166 650898 404250 651134
rect 404486 650898 404570 651134
rect 404806 650898 423930 651134
rect 424166 650898 424250 651134
rect 424486 650898 424570 651134
rect 424806 650898 443930 651134
rect 444166 650898 444250 651134
rect 444486 650898 444570 651134
rect 444806 650898 463930 651134
rect 464166 650898 464250 651134
rect 464486 650898 464570 651134
rect 464806 650898 483930 651134
rect 484166 650898 484250 651134
rect 484486 650898 484570 651134
rect 484806 650898 503930 651134
rect 504166 650898 504250 651134
rect 504486 650898 504570 651134
rect 504806 650898 523930 651134
rect 524166 650898 524250 651134
rect 524486 650898 524570 651134
rect 524806 650898 543930 651134
rect 544166 650898 544250 651134
rect 544486 650898 544570 651134
rect 544806 650898 563930 651134
rect 564166 650898 564250 651134
rect 564486 650898 564570 651134
rect 564806 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 33930 619954
rect 34166 619718 34250 619954
rect 34486 619718 34570 619954
rect 34806 619718 53930 619954
rect 54166 619718 54250 619954
rect 54486 619718 54570 619954
rect 54806 619718 73930 619954
rect 74166 619718 74250 619954
rect 74486 619718 74570 619954
rect 74806 619718 93930 619954
rect 94166 619718 94250 619954
rect 94486 619718 94570 619954
rect 94806 619718 113930 619954
rect 114166 619718 114250 619954
rect 114486 619718 114570 619954
rect 114806 619718 133930 619954
rect 134166 619718 134250 619954
rect 134486 619718 134570 619954
rect 134806 619718 153930 619954
rect 154166 619718 154250 619954
rect 154486 619718 154570 619954
rect 154806 619718 173930 619954
rect 174166 619718 174250 619954
rect 174486 619718 174570 619954
rect 174806 619718 193930 619954
rect 194166 619718 194250 619954
rect 194486 619718 194570 619954
rect 194806 619718 213930 619954
rect 214166 619718 214250 619954
rect 214486 619718 214570 619954
rect 214806 619718 233930 619954
rect 234166 619718 234250 619954
rect 234486 619718 234570 619954
rect 234806 619718 253930 619954
rect 254166 619718 254250 619954
rect 254486 619718 254570 619954
rect 254806 619718 273930 619954
rect 274166 619718 274250 619954
rect 274486 619718 274570 619954
rect 274806 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 313930 619954
rect 314166 619718 314250 619954
rect 314486 619718 314570 619954
rect 314806 619718 333930 619954
rect 334166 619718 334250 619954
rect 334486 619718 334570 619954
rect 334806 619718 353930 619954
rect 354166 619718 354250 619954
rect 354486 619718 354570 619954
rect 354806 619718 373930 619954
rect 374166 619718 374250 619954
rect 374486 619718 374570 619954
rect 374806 619718 393930 619954
rect 394166 619718 394250 619954
rect 394486 619718 394570 619954
rect 394806 619718 413930 619954
rect 414166 619718 414250 619954
rect 414486 619718 414570 619954
rect 414806 619718 433930 619954
rect 434166 619718 434250 619954
rect 434486 619718 434570 619954
rect 434806 619718 453930 619954
rect 454166 619718 454250 619954
rect 454486 619718 454570 619954
rect 454806 619718 473930 619954
rect 474166 619718 474250 619954
rect 474486 619718 474570 619954
rect 474806 619718 493930 619954
rect 494166 619718 494250 619954
rect 494486 619718 494570 619954
rect 494806 619718 513930 619954
rect 514166 619718 514250 619954
rect 514486 619718 514570 619954
rect 514806 619718 533930 619954
rect 534166 619718 534250 619954
rect 534486 619718 534570 619954
rect 534806 619718 553930 619954
rect 554166 619718 554250 619954
rect 554486 619718 554570 619954
rect 554806 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 33930 619634
rect 34166 619398 34250 619634
rect 34486 619398 34570 619634
rect 34806 619398 53930 619634
rect 54166 619398 54250 619634
rect 54486 619398 54570 619634
rect 54806 619398 73930 619634
rect 74166 619398 74250 619634
rect 74486 619398 74570 619634
rect 74806 619398 93930 619634
rect 94166 619398 94250 619634
rect 94486 619398 94570 619634
rect 94806 619398 113930 619634
rect 114166 619398 114250 619634
rect 114486 619398 114570 619634
rect 114806 619398 133930 619634
rect 134166 619398 134250 619634
rect 134486 619398 134570 619634
rect 134806 619398 153930 619634
rect 154166 619398 154250 619634
rect 154486 619398 154570 619634
rect 154806 619398 173930 619634
rect 174166 619398 174250 619634
rect 174486 619398 174570 619634
rect 174806 619398 193930 619634
rect 194166 619398 194250 619634
rect 194486 619398 194570 619634
rect 194806 619398 213930 619634
rect 214166 619398 214250 619634
rect 214486 619398 214570 619634
rect 214806 619398 233930 619634
rect 234166 619398 234250 619634
rect 234486 619398 234570 619634
rect 234806 619398 253930 619634
rect 254166 619398 254250 619634
rect 254486 619398 254570 619634
rect 254806 619398 273930 619634
rect 274166 619398 274250 619634
rect 274486 619398 274570 619634
rect 274806 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 313930 619634
rect 314166 619398 314250 619634
rect 314486 619398 314570 619634
rect 314806 619398 333930 619634
rect 334166 619398 334250 619634
rect 334486 619398 334570 619634
rect 334806 619398 353930 619634
rect 354166 619398 354250 619634
rect 354486 619398 354570 619634
rect 354806 619398 373930 619634
rect 374166 619398 374250 619634
rect 374486 619398 374570 619634
rect 374806 619398 393930 619634
rect 394166 619398 394250 619634
rect 394486 619398 394570 619634
rect 394806 619398 413930 619634
rect 414166 619398 414250 619634
rect 414486 619398 414570 619634
rect 414806 619398 433930 619634
rect 434166 619398 434250 619634
rect 434486 619398 434570 619634
rect 434806 619398 453930 619634
rect 454166 619398 454250 619634
rect 454486 619398 454570 619634
rect 454806 619398 473930 619634
rect 474166 619398 474250 619634
rect 474486 619398 474570 619634
rect 474806 619398 493930 619634
rect 494166 619398 494250 619634
rect 494486 619398 494570 619634
rect 494806 619398 513930 619634
rect 514166 619398 514250 619634
rect 514486 619398 514570 619634
rect 514806 619398 533930 619634
rect 534166 619398 534250 619634
rect 534486 619398 534570 619634
rect 534806 619398 553930 619634
rect 554166 619398 554250 619634
rect 554486 619398 554570 619634
rect 554806 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 23930 615454
rect 24166 615218 24250 615454
rect 24486 615218 24570 615454
rect 24806 615218 43930 615454
rect 44166 615218 44250 615454
rect 44486 615218 44570 615454
rect 44806 615218 63930 615454
rect 64166 615218 64250 615454
rect 64486 615218 64570 615454
rect 64806 615218 83930 615454
rect 84166 615218 84250 615454
rect 84486 615218 84570 615454
rect 84806 615218 103930 615454
rect 104166 615218 104250 615454
rect 104486 615218 104570 615454
rect 104806 615218 123930 615454
rect 124166 615218 124250 615454
rect 124486 615218 124570 615454
rect 124806 615218 143930 615454
rect 144166 615218 144250 615454
rect 144486 615218 144570 615454
rect 144806 615218 163930 615454
rect 164166 615218 164250 615454
rect 164486 615218 164570 615454
rect 164806 615218 183930 615454
rect 184166 615218 184250 615454
rect 184486 615218 184570 615454
rect 184806 615218 203930 615454
rect 204166 615218 204250 615454
rect 204486 615218 204570 615454
rect 204806 615218 223930 615454
rect 224166 615218 224250 615454
rect 224486 615218 224570 615454
rect 224806 615218 243930 615454
rect 244166 615218 244250 615454
rect 244486 615218 244570 615454
rect 244806 615218 263930 615454
rect 264166 615218 264250 615454
rect 264486 615218 264570 615454
rect 264806 615218 283930 615454
rect 284166 615218 284250 615454
rect 284486 615218 284570 615454
rect 284806 615218 303930 615454
rect 304166 615218 304250 615454
rect 304486 615218 304570 615454
rect 304806 615218 323930 615454
rect 324166 615218 324250 615454
rect 324486 615218 324570 615454
rect 324806 615218 343930 615454
rect 344166 615218 344250 615454
rect 344486 615218 344570 615454
rect 344806 615218 363930 615454
rect 364166 615218 364250 615454
rect 364486 615218 364570 615454
rect 364806 615218 383930 615454
rect 384166 615218 384250 615454
rect 384486 615218 384570 615454
rect 384806 615218 403930 615454
rect 404166 615218 404250 615454
rect 404486 615218 404570 615454
rect 404806 615218 423930 615454
rect 424166 615218 424250 615454
rect 424486 615218 424570 615454
rect 424806 615218 443930 615454
rect 444166 615218 444250 615454
rect 444486 615218 444570 615454
rect 444806 615218 463930 615454
rect 464166 615218 464250 615454
rect 464486 615218 464570 615454
rect 464806 615218 483930 615454
rect 484166 615218 484250 615454
rect 484486 615218 484570 615454
rect 484806 615218 503930 615454
rect 504166 615218 504250 615454
rect 504486 615218 504570 615454
rect 504806 615218 523930 615454
rect 524166 615218 524250 615454
rect 524486 615218 524570 615454
rect 524806 615218 543930 615454
rect 544166 615218 544250 615454
rect 544486 615218 544570 615454
rect 544806 615218 563930 615454
rect 564166 615218 564250 615454
rect 564486 615218 564570 615454
rect 564806 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 23930 615134
rect 24166 614898 24250 615134
rect 24486 614898 24570 615134
rect 24806 614898 43930 615134
rect 44166 614898 44250 615134
rect 44486 614898 44570 615134
rect 44806 614898 63930 615134
rect 64166 614898 64250 615134
rect 64486 614898 64570 615134
rect 64806 614898 83930 615134
rect 84166 614898 84250 615134
rect 84486 614898 84570 615134
rect 84806 614898 103930 615134
rect 104166 614898 104250 615134
rect 104486 614898 104570 615134
rect 104806 614898 123930 615134
rect 124166 614898 124250 615134
rect 124486 614898 124570 615134
rect 124806 614898 143930 615134
rect 144166 614898 144250 615134
rect 144486 614898 144570 615134
rect 144806 614898 163930 615134
rect 164166 614898 164250 615134
rect 164486 614898 164570 615134
rect 164806 614898 183930 615134
rect 184166 614898 184250 615134
rect 184486 614898 184570 615134
rect 184806 614898 203930 615134
rect 204166 614898 204250 615134
rect 204486 614898 204570 615134
rect 204806 614898 223930 615134
rect 224166 614898 224250 615134
rect 224486 614898 224570 615134
rect 224806 614898 243930 615134
rect 244166 614898 244250 615134
rect 244486 614898 244570 615134
rect 244806 614898 263930 615134
rect 264166 614898 264250 615134
rect 264486 614898 264570 615134
rect 264806 614898 283930 615134
rect 284166 614898 284250 615134
rect 284486 614898 284570 615134
rect 284806 614898 303930 615134
rect 304166 614898 304250 615134
rect 304486 614898 304570 615134
rect 304806 614898 323930 615134
rect 324166 614898 324250 615134
rect 324486 614898 324570 615134
rect 324806 614898 343930 615134
rect 344166 614898 344250 615134
rect 344486 614898 344570 615134
rect 344806 614898 363930 615134
rect 364166 614898 364250 615134
rect 364486 614898 364570 615134
rect 364806 614898 383930 615134
rect 384166 614898 384250 615134
rect 384486 614898 384570 615134
rect 384806 614898 403930 615134
rect 404166 614898 404250 615134
rect 404486 614898 404570 615134
rect 404806 614898 423930 615134
rect 424166 614898 424250 615134
rect 424486 614898 424570 615134
rect 424806 614898 443930 615134
rect 444166 614898 444250 615134
rect 444486 614898 444570 615134
rect 444806 614898 463930 615134
rect 464166 614898 464250 615134
rect 464486 614898 464570 615134
rect 464806 614898 483930 615134
rect 484166 614898 484250 615134
rect 484486 614898 484570 615134
rect 484806 614898 503930 615134
rect 504166 614898 504250 615134
rect 504486 614898 504570 615134
rect 504806 614898 523930 615134
rect 524166 614898 524250 615134
rect 524486 614898 524570 615134
rect 524806 614898 543930 615134
rect 544166 614898 544250 615134
rect 544486 614898 544570 615134
rect 544806 614898 563930 615134
rect 564166 614898 564250 615134
rect 564486 614898 564570 615134
rect 564806 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 33930 547954
rect 34166 547718 34250 547954
rect 34486 547718 34570 547954
rect 34806 547718 53930 547954
rect 54166 547718 54250 547954
rect 54486 547718 54570 547954
rect 54806 547718 73930 547954
rect 74166 547718 74250 547954
rect 74486 547718 74570 547954
rect 74806 547718 93930 547954
rect 94166 547718 94250 547954
rect 94486 547718 94570 547954
rect 94806 547718 113930 547954
rect 114166 547718 114250 547954
rect 114486 547718 114570 547954
rect 114806 547718 133930 547954
rect 134166 547718 134250 547954
rect 134486 547718 134570 547954
rect 134806 547718 153930 547954
rect 154166 547718 154250 547954
rect 154486 547718 154570 547954
rect 154806 547718 173930 547954
rect 174166 547718 174250 547954
rect 174486 547718 174570 547954
rect 174806 547718 193930 547954
rect 194166 547718 194250 547954
rect 194486 547718 194570 547954
rect 194806 547718 213930 547954
rect 214166 547718 214250 547954
rect 214486 547718 214570 547954
rect 214806 547718 233930 547954
rect 234166 547718 234250 547954
rect 234486 547718 234570 547954
rect 234806 547718 253930 547954
rect 254166 547718 254250 547954
rect 254486 547718 254570 547954
rect 254806 547718 273930 547954
rect 274166 547718 274250 547954
rect 274486 547718 274570 547954
rect 274806 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 313930 547954
rect 314166 547718 314250 547954
rect 314486 547718 314570 547954
rect 314806 547718 333930 547954
rect 334166 547718 334250 547954
rect 334486 547718 334570 547954
rect 334806 547718 353930 547954
rect 354166 547718 354250 547954
rect 354486 547718 354570 547954
rect 354806 547718 373930 547954
rect 374166 547718 374250 547954
rect 374486 547718 374570 547954
rect 374806 547718 393930 547954
rect 394166 547718 394250 547954
rect 394486 547718 394570 547954
rect 394806 547718 413930 547954
rect 414166 547718 414250 547954
rect 414486 547718 414570 547954
rect 414806 547718 433930 547954
rect 434166 547718 434250 547954
rect 434486 547718 434570 547954
rect 434806 547718 453930 547954
rect 454166 547718 454250 547954
rect 454486 547718 454570 547954
rect 454806 547718 473930 547954
rect 474166 547718 474250 547954
rect 474486 547718 474570 547954
rect 474806 547718 493930 547954
rect 494166 547718 494250 547954
rect 494486 547718 494570 547954
rect 494806 547718 513930 547954
rect 514166 547718 514250 547954
rect 514486 547718 514570 547954
rect 514806 547718 533930 547954
rect 534166 547718 534250 547954
rect 534486 547718 534570 547954
rect 534806 547718 553930 547954
rect 554166 547718 554250 547954
rect 554486 547718 554570 547954
rect 554806 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 33930 547634
rect 34166 547398 34250 547634
rect 34486 547398 34570 547634
rect 34806 547398 53930 547634
rect 54166 547398 54250 547634
rect 54486 547398 54570 547634
rect 54806 547398 73930 547634
rect 74166 547398 74250 547634
rect 74486 547398 74570 547634
rect 74806 547398 93930 547634
rect 94166 547398 94250 547634
rect 94486 547398 94570 547634
rect 94806 547398 113930 547634
rect 114166 547398 114250 547634
rect 114486 547398 114570 547634
rect 114806 547398 133930 547634
rect 134166 547398 134250 547634
rect 134486 547398 134570 547634
rect 134806 547398 153930 547634
rect 154166 547398 154250 547634
rect 154486 547398 154570 547634
rect 154806 547398 173930 547634
rect 174166 547398 174250 547634
rect 174486 547398 174570 547634
rect 174806 547398 193930 547634
rect 194166 547398 194250 547634
rect 194486 547398 194570 547634
rect 194806 547398 213930 547634
rect 214166 547398 214250 547634
rect 214486 547398 214570 547634
rect 214806 547398 233930 547634
rect 234166 547398 234250 547634
rect 234486 547398 234570 547634
rect 234806 547398 253930 547634
rect 254166 547398 254250 547634
rect 254486 547398 254570 547634
rect 254806 547398 273930 547634
rect 274166 547398 274250 547634
rect 274486 547398 274570 547634
rect 274806 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 313930 547634
rect 314166 547398 314250 547634
rect 314486 547398 314570 547634
rect 314806 547398 333930 547634
rect 334166 547398 334250 547634
rect 334486 547398 334570 547634
rect 334806 547398 353930 547634
rect 354166 547398 354250 547634
rect 354486 547398 354570 547634
rect 354806 547398 373930 547634
rect 374166 547398 374250 547634
rect 374486 547398 374570 547634
rect 374806 547398 393930 547634
rect 394166 547398 394250 547634
rect 394486 547398 394570 547634
rect 394806 547398 413930 547634
rect 414166 547398 414250 547634
rect 414486 547398 414570 547634
rect 414806 547398 433930 547634
rect 434166 547398 434250 547634
rect 434486 547398 434570 547634
rect 434806 547398 453930 547634
rect 454166 547398 454250 547634
rect 454486 547398 454570 547634
rect 454806 547398 473930 547634
rect 474166 547398 474250 547634
rect 474486 547398 474570 547634
rect 474806 547398 493930 547634
rect 494166 547398 494250 547634
rect 494486 547398 494570 547634
rect 494806 547398 513930 547634
rect 514166 547398 514250 547634
rect 514486 547398 514570 547634
rect 514806 547398 533930 547634
rect 534166 547398 534250 547634
rect 534486 547398 534570 547634
rect 534806 547398 553930 547634
rect 554166 547398 554250 547634
rect 554486 547398 554570 547634
rect 554806 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 23930 543454
rect 24166 543218 24250 543454
rect 24486 543218 24570 543454
rect 24806 543218 43930 543454
rect 44166 543218 44250 543454
rect 44486 543218 44570 543454
rect 44806 543218 63930 543454
rect 64166 543218 64250 543454
rect 64486 543218 64570 543454
rect 64806 543218 83930 543454
rect 84166 543218 84250 543454
rect 84486 543218 84570 543454
rect 84806 543218 103930 543454
rect 104166 543218 104250 543454
rect 104486 543218 104570 543454
rect 104806 543218 123930 543454
rect 124166 543218 124250 543454
rect 124486 543218 124570 543454
rect 124806 543218 143930 543454
rect 144166 543218 144250 543454
rect 144486 543218 144570 543454
rect 144806 543218 163930 543454
rect 164166 543218 164250 543454
rect 164486 543218 164570 543454
rect 164806 543218 183930 543454
rect 184166 543218 184250 543454
rect 184486 543218 184570 543454
rect 184806 543218 203930 543454
rect 204166 543218 204250 543454
rect 204486 543218 204570 543454
rect 204806 543218 223930 543454
rect 224166 543218 224250 543454
rect 224486 543218 224570 543454
rect 224806 543218 243930 543454
rect 244166 543218 244250 543454
rect 244486 543218 244570 543454
rect 244806 543218 263930 543454
rect 264166 543218 264250 543454
rect 264486 543218 264570 543454
rect 264806 543218 283930 543454
rect 284166 543218 284250 543454
rect 284486 543218 284570 543454
rect 284806 543218 303930 543454
rect 304166 543218 304250 543454
rect 304486 543218 304570 543454
rect 304806 543218 323930 543454
rect 324166 543218 324250 543454
rect 324486 543218 324570 543454
rect 324806 543218 343930 543454
rect 344166 543218 344250 543454
rect 344486 543218 344570 543454
rect 344806 543218 363930 543454
rect 364166 543218 364250 543454
rect 364486 543218 364570 543454
rect 364806 543218 383930 543454
rect 384166 543218 384250 543454
rect 384486 543218 384570 543454
rect 384806 543218 403930 543454
rect 404166 543218 404250 543454
rect 404486 543218 404570 543454
rect 404806 543218 423930 543454
rect 424166 543218 424250 543454
rect 424486 543218 424570 543454
rect 424806 543218 443930 543454
rect 444166 543218 444250 543454
rect 444486 543218 444570 543454
rect 444806 543218 463930 543454
rect 464166 543218 464250 543454
rect 464486 543218 464570 543454
rect 464806 543218 483930 543454
rect 484166 543218 484250 543454
rect 484486 543218 484570 543454
rect 484806 543218 503930 543454
rect 504166 543218 504250 543454
rect 504486 543218 504570 543454
rect 504806 543218 523930 543454
rect 524166 543218 524250 543454
rect 524486 543218 524570 543454
rect 524806 543218 543930 543454
rect 544166 543218 544250 543454
rect 544486 543218 544570 543454
rect 544806 543218 563930 543454
rect 564166 543218 564250 543454
rect 564486 543218 564570 543454
rect 564806 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 23930 543134
rect 24166 542898 24250 543134
rect 24486 542898 24570 543134
rect 24806 542898 43930 543134
rect 44166 542898 44250 543134
rect 44486 542898 44570 543134
rect 44806 542898 63930 543134
rect 64166 542898 64250 543134
rect 64486 542898 64570 543134
rect 64806 542898 83930 543134
rect 84166 542898 84250 543134
rect 84486 542898 84570 543134
rect 84806 542898 103930 543134
rect 104166 542898 104250 543134
rect 104486 542898 104570 543134
rect 104806 542898 123930 543134
rect 124166 542898 124250 543134
rect 124486 542898 124570 543134
rect 124806 542898 143930 543134
rect 144166 542898 144250 543134
rect 144486 542898 144570 543134
rect 144806 542898 163930 543134
rect 164166 542898 164250 543134
rect 164486 542898 164570 543134
rect 164806 542898 183930 543134
rect 184166 542898 184250 543134
rect 184486 542898 184570 543134
rect 184806 542898 203930 543134
rect 204166 542898 204250 543134
rect 204486 542898 204570 543134
rect 204806 542898 223930 543134
rect 224166 542898 224250 543134
rect 224486 542898 224570 543134
rect 224806 542898 243930 543134
rect 244166 542898 244250 543134
rect 244486 542898 244570 543134
rect 244806 542898 263930 543134
rect 264166 542898 264250 543134
rect 264486 542898 264570 543134
rect 264806 542898 283930 543134
rect 284166 542898 284250 543134
rect 284486 542898 284570 543134
rect 284806 542898 303930 543134
rect 304166 542898 304250 543134
rect 304486 542898 304570 543134
rect 304806 542898 323930 543134
rect 324166 542898 324250 543134
rect 324486 542898 324570 543134
rect 324806 542898 343930 543134
rect 344166 542898 344250 543134
rect 344486 542898 344570 543134
rect 344806 542898 363930 543134
rect 364166 542898 364250 543134
rect 364486 542898 364570 543134
rect 364806 542898 383930 543134
rect 384166 542898 384250 543134
rect 384486 542898 384570 543134
rect 384806 542898 403930 543134
rect 404166 542898 404250 543134
rect 404486 542898 404570 543134
rect 404806 542898 423930 543134
rect 424166 542898 424250 543134
rect 424486 542898 424570 543134
rect 424806 542898 443930 543134
rect 444166 542898 444250 543134
rect 444486 542898 444570 543134
rect 444806 542898 463930 543134
rect 464166 542898 464250 543134
rect 464486 542898 464570 543134
rect 464806 542898 483930 543134
rect 484166 542898 484250 543134
rect 484486 542898 484570 543134
rect 484806 542898 503930 543134
rect 504166 542898 504250 543134
rect 504486 542898 504570 543134
rect 504806 542898 523930 543134
rect 524166 542898 524250 543134
rect 524486 542898 524570 543134
rect 524806 542898 543930 543134
rect 544166 542898 544250 543134
rect 544486 542898 544570 543134
rect 544806 542898 563930 543134
rect 564166 542898 564250 543134
rect 564486 542898 564570 543134
rect 564806 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 33930 511954
rect 34166 511718 34250 511954
rect 34486 511718 34570 511954
rect 34806 511718 53930 511954
rect 54166 511718 54250 511954
rect 54486 511718 54570 511954
rect 54806 511718 73930 511954
rect 74166 511718 74250 511954
rect 74486 511718 74570 511954
rect 74806 511718 93930 511954
rect 94166 511718 94250 511954
rect 94486 511718 94570 511954
rect 94806 511718 113930 511954
rect 114166 511718 114250 511954
rect 114486 511718 114570 511954
rect 114806 511718 133930 511954
rect 134166 511718 134250 511954
rect 134486 511718 134570 511954
rect 134806 511718 153930 511954
rect 154166 511718 154250 511954
rect 154486 511718 154570 511954
rect 154806 511718 173930 511954
rect 174166 511718 174250 511954
rect 174486 511718 174570 511954
rect 174806 511718 193930 511954
rect 194166 511718 194250 511954
rect 194486 511718 194570 511954
rect 194806 511718 213930 511954
rect 214166 511718 214250 511954
rect 214486 511718 214570 511954
rect 214806 511718 233930 511954
rect 234166 511718 234250 511954
rect 234486 511718 234570 511954
rect 234806 511718 253930 511954
rect 254166 511718 254250 511954
rect 254486 511718 254570 511954
rect 254806 511718 273930 511954
rect 274166 511718 274250 511954
rect 274486 511718 274570 511954
rect 274806 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 313930 511954
rect 314166 511718 314250 511954
rect 314486 511718 314570 511954
rect 314806 511718 333930 511954
rect 334166 511718 334250 511954
rect 334486 511718 334570 511954
rect 334806 511718 353930 511954
rect 354166 511718 354250 511954
rect 354486 511718 354570 511954
rect 354806 511718 373930 511954
rect 374166 511718 374250 511954
rect 374486 511718 374570 511954
rect 374806 511718 393930 511954
rect 394166 511718 394250 511954
rect 394486 511718 394570 511954
rect 394806 511718 413930 511954
rect 414166 511718 414250 511954
rect 414486 511718 414570 511954
rect 414806 511718 433930 511954
rect 434166 511718 434250 511954
rect 434486 511718 434570 511954
rect 434806 511718 453930 511954
rect 454166 511718 454250 511954
rect 454486 511718 454570 511954
rect 454806 511718 473930 511954
rect 474166 511718 474250 511954
rect 474486 511718 474570 511954
rect 474806 511718 493930 511954
rect 494166 511718 494250 511954
rect 494486 511718 494570 511954
rect 494806 511718 513930 511954
rect 514166 511718 514250 511954
rect 514486 511718 514570 511954
rect 514806 511718 533930 511954
rect 534166 511718 534250 511954
rect 534486 511718 534570 511954
rect 534806 511718 553930 511954
rect 554166 511718 554250 511954
rect 554486 511718 554570 511954
rect 554806 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 33930 511634
rect 34166 511398 34250 511634
rect 34486 511398 34570 511634
rect 34806 511398 53930 511634
rect 54166 511398 54250 511634
rect 54486 511398 54570 511634
rect 54806 511398 73930 511634
rect 74166 511398 74250 511634
rect 74486 511398 74570 511634
rect 74806 511398 93930 511634
rect 94166 511398 94250 511634
rect 94486 511398 94570 511634
rect 94806 511398 113930 511634
rect 114166 511398 114250 511634
rect 114486 511398 114570 511634
rect 114806 511398 133930 511634
rect 134166 511398 134250 511634
rect 134486 511398 134570 511634
rect 134806 511398 153930 511634
rect 154166 511398 154250 511634
rect 154486 511398 154570 511634
rect 154806 511398 173930 511634
rect 174166 511398 174250 511634
rect 174486 511398 174570 511634
rect 174806 511398 193930 511634
rect 194166 511398 194250 511634
rect 194486 511398 194570 511634
rect 194806 511398 213930 511634
rect 214166 511398 214250 511634
rect 214486 511398 214570 511634
rect 214806 511398 233930 511634
rect 234166 511398 234250 511634
rect 234486 511398 234570 511634
rect 234806 511398 253930 511634
rect 254166 511398 254250 511634
rect 254486 511398 254570 511634
rect 254806 511398 273930 511634
rect 274166 511398 274250 511634
rect 274486 511398 274570 511634
rect 274806 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 313930 511634
rect 314166 511398 314250 511634
rect 314486 511398 314570 511634
rect 314806 511398 333930 511634
rect 334166 511398 334250 511634
rect 334486 511398 334570 511634
rect 334806 511398 353930 511634
rect 354166 511398 354250 511634
rect 354486 511398 354570 511634
rect 354806 511398 373930 511634
rect 374166 511398 374250 511634
rect 374486 511398 374570 511634
rect 374806 511398 393930 511634
rect 394166 511398 394250 511634
rect 394486 511398 394570 511634
rect 394806 511398 413930 511634
rect 414166 511398 414250 511634
rect 414486 511398 414570 511634
rect 414806 511398 433930 511634
rect 434166 511398 434250 511634
rect 434486 511398 434570 511634
rect 434806 511398 453930 511634
rect 454166 511398 454250 511634
rect 454486 511398 454570 511634
rect 454806 511398 473930 511634
rect 474166 511398 474250 511634
rect 474486 511398 474570 511634
rect 474806 511398 493930 511634
rect 494166 511398 494250 511634
rect 494486 511398 494570 511634
rect 494806 511398 513930 511634
rect 514166 511398 514250 511634
rect 514486 511398 514570 511634
rect 514806 511398 533930 511634
rect 534166 511398 534250 511634
rect 534486 511398 534570 511634
rect 534806 511398 553930 511634
rect 554166 511398 554250 511634
rect 554486 511398 554570 511634
rect 554806 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 23930 507454
rect 24166 507218 24250 507454
rect 24486 507218 24570 507454
rect 24806 507218 43930 507454
rect 44166 507218 44250 507454
rect 44486 507218 44570 507454
rect 44806 507218 63930 507454
rect 64166 507218 64250 507454
rect 64486 507218 64570 507454
rect 64806 507218 83930 507454
rect 84166 507218 84250 507454
rect 84486 507218 84570 507454
rect 84806 507218 103930 507454
rect 104166 507218 104250 507454
rect 104486 507218 104570 507454
rect 104806 507218 123930 507454
rect 124166 507218 124250 507454
rect 124486 507218 124570 507454
rect 124806 507218 143930 507454
rect 144166 507218 144250 507454
rect 144486 507218 144570 507454
rect 144806 507218 163930 507454
rect 164166 507218 164250 507454
rect 164486 507218 164570 507454
rect 164806 507218 183930 507454
rect 184166 507218 184250 507454
rect 184486 507218 184570 507454
rect 184806 507218 203930 507454
rect 204166 507218 204250 507454
rect 204486 507218 204570 507454
rect 204806 507218 223930 507454
rect 224166 507218 224250 507454
rect 224486 507218 224570 507454
rect 224806 507218 243930 507454
rect 244166 507218 244250 507454
rect 244486 507218 244570 507454
rect 244806 507218 263930 507454
rect 264166 507218 264250 507454
rect 264486 507218 264570 507454
rect 264806 507218 283930 507454
rect 284166 507218 284250 507454
rect 284486 507218 284570 507454
rect 284806 507218 303930 507454
rect 304166 507218 304250 507454
rect 304486 507218 304570 507454
rect 304806 507218 323930 507454
rect 324166 507218 324250 507454
rect 324486 507218 324570 507454
rect 324806 507218 343930 507454
rect 344166 507218 344250 507454
rect 344486 507218 344570 507454
rect 344806 507218 363930 507454
rect 364166 507218 364250 507454
rect 364486 507218 364570 507454
rect 364806 507218 383930 507454
rect 384166 507218 384250 507454
rect 384486 507218 384570 507454
rect 384806 507218 403930 507454
rect 404166 507218 404250 507454
rect 404486 507218 404570 507454
rect 404806 507218 423930 507454
rect 424166 507218 424250 507454
rect 424486 507218 424570 507454
rect 424806 507218 443930 507454
rect 444166 507218 444250 507454
rect 444486 507218 444570 507454
rect 444806 507218 463930 507454
rect 464166 507218 464250 507454
rect 464486 507218 464570 507454
rect 464806 507218 483930 507454
rect 484166 507218 484250 507454
rect 484486 507218 484570 507454
rect 484806 507218 503930 507454
rect 504166 507218 504250 507454
rect 504486 507218 504570 507454
rect 504806 507218 523930 507454
rect 524166 507218 524250 507454
rect 524486 507218 524570 507454
rect 524806 507218 543930 507454
rect 544166 507218 544250 507454
rect 544486 507218 544570 507454
rect 544806 507218 563930 507454
rect 564166 507218 564250 507454
rect 564486 507218 564570 507454
rect 564806 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 23930 507134
rect 24166 506898 24250 507134
rect 24486 506898 24570 507134
rect 24806 506898 43930 507134
rect 44166 506898 44250 507134
rect 44486 506898 44570 507134
rect 44806 506898 63930 507134
rect 64166 506898 64250 507134
rect 64486 506898 64570 507134
rect 64806 506898 83930 507134
rect 84166 506898 84250 507134
rect 84486 506898 84570 507134
rect 84806 506898 103930 507134
rect 104166 506898 104250 507134
rect 104486 506898 104570 507134
rect 104806 506898 123930 507134
rect 124166 506898 124250 507134
rect 124486 506898 124570 507134
rect 124806 506898 143930 507134
rect 144166 506898 144250 507134
rect 144486 506898 144570 507134
rect 144806 506898 163930 507134
rect 164166 506898 164250 507134
rect 164486 506898 164570 507134
rect 164806 506898 183930 507134
rect 184166 506898 184250 507134
rect 184486 506898 184570 507134
rect 184806 506898 203930 507134
rect 204166 506898 204250 507134
rect 204486 506898 204570 507134
rect 204806 506898 223930 507134
rect 224166 506898 224250 507134
rect 224486 506898 224570 507134
rect 224806 506898 243930 507134
rect 244166 506898 244250 507134
rect 244486 506898 244570 507134
rect 244806 506898 263930 507134
rect 264166 506898 264250 507134
rect 264486 506898 264570 507134
rect 264806 506898 283930 507134
rect 284166 506898 284250 507134
rect 284486 506898 284570 507134
rect 284806 506898 303930 507134
rect 304166 506898 304250 507134
rect 304486 506898 304570 507134
rect 304806 506898 323930 507134
rect 324166 506898 324250 507134
rect 324486 506898 324570 507134
rect 324806 506898 343930 507134
rect 344166 506898 344250 507134
rect 344486 506898 344570 507134
rect 344806 506898 363930 507134
rect 364166 506898 364250 507134
rect 364486 506898 364570 507134
rect 364806 506898 383930 507134
rect 384166 506898 384250 507134
rect 384486 506898 384570 507134
rect 384806 506898 403930 507134
rect 404166 506898 404250 507134
rect 404486 506898 404570 507134
rect 404806 506898 423930 507134
rect 424166 506898 424250 507134
rect 424486 506898 424570 507134
rect 424806 506898 443930 507134
rect 444166 506898 444250 507134
rect 444486 506898 444570 507134
rect 444806 506898 463930 507134
rect 464166 506898 464250 507134
rect 464486 506898 464570 507134
rect 464806 506898 483930 507134
rect 484166 506898 484250 507134
rect 484486 506898 484570 507134
rect 484806 506898 503930 507134
rect 504166 506898 504250 507134
rect 504486 506898 504570 507134
rect 504806 506898 523930 507134
rect 524166 506898 524250 507134
rect 524486 506898 524570 507134
rect 524806 506898 543930 507134
rect 544166 506898 544250 507134
rect 544486 506898 544570 507134
rect 544806 506898 563930 507134
rect 564166 506898 564250 507134
rect 564486 506898 564570 507134
rect 564806 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 33930 475954
rect 34166 475718 34250 475954
rect 34486 475718 34570 475954
rect 34806 475718 53930 475954
rect 54166 475718 54250 475954
rect 54486 475718 54570 475954
rect 54806 475718 73930 475954
rect 74166 475718 74250 475954
rect 74486 475718 74570 475954
rect 74806 475718 93930 475954
rect 94166 475718 94250 475954
rect 94486 475718 94570 475954
rect 94806 475718 113930 475954
rect 114166 475718 114250 475954
rect 114486 475718 114570 475954
rect 114806 475718 133930 475954
rect 134166 475718 134250 475954
rect 134486 475718 134570 475954
rect 134806 475718 153930 475954
rect 154166 475718 154250 475954
rect 154486 475718 154570 475954
rect 154806 475718 173930 475954
rect 174166 475718 174250 475954
rect 174486 475718 174570 475954
rect 174806 475718 193930 475954
rect 194166 475718 194250 475954
rect 194486 475718 194570 475954
rect 194806 475718 213930 475954
rect 214166 475718 214250 475954
rect 214486 475718 214570 475954
rect 214806 475718 233930 475954
rect 234166 475718 234250 475954
rect 234486 475718 234570 475954
rect 234806 475718 253930 475954
rect 254166 475718 254250 475954
rect 254486 475718 254570 475954
rect 254806 475718 273930 475954
rect 274166 475718 274250 475954
rect 274486 475718 274570 475954
rect 274806 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 313930 475954
rect 314166 475718 314250 475954
rect 314486 475718 314570 475954
rect 314806 475718 333930 475954
rect 334166 475718 334250 475954
rect 334486 475718 334570 475954
rect 334806 475718 353930 475954
rect 354166 475718 354250 475954
rect 354486 475718 354570 475954
rect 354806 475718 373930 475954
rect 374166 475718 374250 475954
rect 374486 475718 374570 475954
rect 374806 475718 393930 475954
rect 394166 475718 394250 475954
rect 394486 475718 394570 475954
rect 394806 475718 413930 475954
rect 414166 475718 414250 475954
rect 414486 475718 414570 475954
rect 414806 475718 433930 475954
rect 434166 475718 434250 475954
rect 434486 475718 434570 475954
rect 434806 475718 453930 475954
rect 454166 475718 454250 475954
rect 454486 475718 454570 475954
rect 454806 475718 473930 475954
rect 474166 475718 474250 475954
rect 474486 475718 474570 475954
rect 474806 475718 493930 475954
rect 494166 475718 494250 475954
rect 494486 475718 494570 475954
rect 494806 475718 513930 475954
rect 514166 475718 514250 475954
rect 514486 475718 514570 475954
rect 514806 475718 533930 475954
rect 534166 475718 534250 475954
rect 534486 475718 534570 475954
rect 534806 475718 553930 475954
rect 554166 475718 554250 475954
rect 554486 475718 554570 475954
rect 554806 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 33930 475634
rect 34166 475398 34250 475634
rect 34486 475398 34570 475634
rect 34806 475398 53930 475634
rect 54166 475398 54250 475634
rect 54486 475398 54570 475634
rect 54806 475398 73930 475634
rect 74166 475398 74250 475634
rect 74486 475398 74570 475634
rect 74806 475398 93930 475634
rect 94166 475398 94250 475634
rect 94486 475398 94570 475634
rect 94806 475398 113930 475634
rect 114166 475398 114250 475634
rect 114486 475398 114570 475634
rect 114806 475398 133930 475634
rect 134166 475398 134250 475634
rect 134486 475398 134570 475634
rect 134806 475398 153930 475634
rect 154166 475398 154250 475634
rect 154486 475398 154570 475634
rect 154806 475398 173930 475634
rect 174166 475398 174250 475634
rect 174486 475398 174570 475634
rect 174806 475398 193930 475634
rect 194166 475398 194250 475634
rect 194486 475398 194570 475634
rect 194806 475398 213930 475634
rect 214166 475398 214250 475634
rect 214486 475398 214570 475634
rect 214806 475398 233930 475634
rect 234166 475398 234250 475634
rect 234486 475398 234570 475634
rect 234806 475398 253930 475634
rect 254166 475398 254250 475634
rect 254486 475398 254570 475634
rect 254806 475398 273930 475634
rect 274166 475398 274250 475634
rect 274486 475398 274570 475634
rect 274806 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 313930 475634
rect 314166 475398 314250 475634
rect 314486 475398 314570 475634
rect 314806 475398 333930 475634
rect 334166 475398 334250 475634
rect 334486 475398 334570 475634
rect 334806 475398 353930 475634
rect 354166 475398 354250 475634
rect 354486 475398 354570 475634
rect 354806 475398 373930 475634
rect 374166 475398 374250 475634
rect 374486 475398 374570 475634
rect 374806 475398 393930 475634
rect 394166 475398 394250 475634
rect 394486 475398 394570 475634
rect 394806 475398 413930 475634
rect 414166 475398 414250 475634
rect 414486 475398 414570 475634
rect 414806 475398 433930 475634
rect 434166 475398 434250 475634
rect 434486 475398 434570 475634
rect 434806 475398 453930 475634
rect 454166 475398 454250 475634
rect 454486 475398 454570 475634
rect 454806 475398 473930 475634
rect 474166 475398 474250 475634
rect 474486 475398 474570 475634
rect 474806 475398 493930 475634
rect 494166 475398 494250 475634
rect 494486 475398 494570 475634
rect 494806 475398 513930 475634
rect 514166 475398 514250 475634
rect 514486 475398 514570 475634
rect 514806 475398 533930 475634
rect 534166 475398 534250 475634
rect 534486 475398 534570 475634
rect 534806 475398 553930 475634
rect 554166 475398 554250 475634
rect 554486 475398 554570 475634
rect 554806 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 23930 471454
rect 24166 471218 24250 471454
rect 24486 471218 24570 471454
rect 24806 471218 43930 471454
rect 44166 471218 44250 471454
rect 44486 471218 44570 471454
rect 44806 471218 63930 471454
rect 64166 471218 64250 471454
rect 64486 471218 64570 471454
rect 64806 471218 83930 471454
rect 84166 471218 84250 471454
rect 84486 471218 84570 471454
rect 84806 471218 103930 471454
rect 104166 471218 104250 471454
rect 104486 471218 104570 471454
rect 104806 471218 123930 471454
rect 124166 471218 124250 471454
rect 124486 471218 124570 471454
rect 124806 471218 143930 471454
rect 144166 471218 144250 471454
rect 144486 471218 144570 471454
rect 144806 471218 163930 471454
rect 164166 471218 164250 471454
rect 164486 471218 164570 471454
rect 164806 471218 183930 471454
rect 184166 471218 184250 471454
rect 184486 471218 184570 471454
rect 184806 471218 203930 471454
rect 204166 471218 204250 471454
rect 204486 471218 204570 471454
rect 204806 471218 223930 471454
rect 224166 471218 224250 471454
rect 224486 471218 224570 471454
rect 224806 471218 243930 471454
rect 244166 471218 244250 471454
rect 244486 471218 244570 471454
rect 244806 471218 263930 471454
rect 264166 471218 264250 471454
rect 264486 471218 264570 471454
rect 264806 471218 283930 471454
rect 284166 471218 284250 471454
rect 284486 471218 284570 471454
rect 284806 471218 303930 471454
rect 304166 471218 304250 471454
rect 304486 471218 304570 471454
rect 304806 471218 323930 471454
rect 324166 471218 324250 471454
rect 324486 471218 324570 471454
rect 324806 471218 343930 471454
rect 344166 471218 344250 471454
rect 344486 471218 344570 471454
rect 344806 471218 363930 471454
rect 364166 471218 364250 471454
rect 364486 471218 364570 471454
rect 364806 471218 383930 471454
rect 384166 471218 384250 471454
rect 384486 471218 384570 471454
rect 384806 471218 403930 471454
rect 404166 471218 404250 471454
rect 404486 471218 404570 471454
rect 404806 471218 423930 471454
rect 424166 471218 424250 471454
rect 424486 471218 424570 471454
rect 424806 471218 443930 471454
rect 444166 471218 444250 471454
rect 444486 471218 444570 471454
rect 444806 471218 463930 471454
rect 464166 471218 464250 471454
rect 464486 471218 464570 471454
rect 464806 471218 483930 471454
rect 484166 471218 484250 471454
rect 484486 471218 484570 471454
rect 484806 471218 503930 471454
rect 504166 471218 504250 471454
rect 504486 471218 504570 471454
rect 504806 471218 523930 471454
rect 524166 471218 524250 471454
rect 524486 471218 524570 471454
rect 524806 471218 543930 471454
rect 544166 471218 544250 471454
rect 544486 471218 544570 471454
rect 544806 471218 563930 471454
rect 564166 471218 564250 471454
rect 564486 471218 564570 471454
rect 564806 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 23930 471134
rect 24166 470898 24250 471134
rect 24486 470898 24570 471134
rect 24806 470898 43930 471134
rect 44166 470898 44250 471134
rect 44486 470898 44570 471134
rect 44806 470898 63930 471134
rect 64166 470898 64250 471134
rect 64486 470898 64570 471134
rect 64806 470898 83930 471134
rect 84166 470898 84250 471134
rect 84486 470898 84570 471134
rect 84806 470898 103930 471134
rect 104166 470898 104250 471134
rect 104486 470898 104570 471134
rect 104806 470898 123930 471134
rect 124166 470898 124250 471134
rect 124486 470898 124570 471134
rect 124806 470898 143930 471134
rect 144166 470898 144250 471134
rect 144486 470898 144570 471134
rect 144806 470898 163930 471134
rect 164166 470898 164250 471134
rect 164486 470898 164570 471134
rect 164806 470898 183930 471134
rect 184166 470898 184250 471134
rect 184486 470898 184570 471134
rect 184806 470898 203930 471134
rect 204166 470898 204250 471134
rect 204486 470898 204570 471134
rect 204806 470898 223930 471134
rect 224166 470898 224250 471134
rect 224486 470898 224570 471134
rect 224806 470898 243930 471134
rect 244166 470898 244250 471134
rect 244486 470898 244570 471134
rect 244806 470898 263930 471134
rect 264166 470898 264250 471134
rect 264486 470898 264570 471134
rect 264806 470898 283930 471134
rect 284166 470898 284250 471134
rect 284486 470898 284570 471134
rect 284806 470898 303930 471134
rect 304166 470898 304250 471134
rect 304486 470898 304570 471134
rect 304806 470898 323930 471134
rect 324166 470898 324250 471134
rect 324486 470898 324570 471134
rect 324806 470898 343930 471134
rect 344166 470898 344250 471134
rect 344486 470898 344570 471134
rect 344806 470898 363930 471134
rect 364166 470898 364250 471134
rect 364486 470898 364570 471134
rect 364806 470898 383930 471134
rect 384166 470898 384250 471134
rect 384486 470898 384570 471134
rect 384806 470898 403930 471134
rect 404166 470898 404250 471134
rect 404486 470898 404570 471134
rect 404806 470898 423930 471134
rect 424166 470898 424250 471134
rect 424486 470898 424570 471134
rect 424806 470898 443930 471134
rect 444166 470898 444250 471134
rect 444486 470898 444570 471134
rect 444806 470898 463930 471134
rect 464166 470898 464250 471134
rect 464486 470898 464570 471134
rect 464806 470898 483930 471134
rect 484166 470898 484250 471134
rect 484486 470898 484570 471134
rect 484806 470898 503930 471134
rect 504166 470898 504250 471134
rect 504486 470898 504570 471134
rect 504806 470898 523930 471134
rect 524166 470898 524250 471134
rect 524486 470898 524570 471134
rect 524806 470898 543930 471134
rect 544166 470898 544250 471134
rect 544486 470898 544570 471134
rect 544806 470898 563930 471134
rect 564166 470898 564250 471134
rect 564486 470898 564570 471134
rect 564806 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 33930 439954
rect 34166 439718 34250 439954
rect 34486 439718 34570 439954
rect 34806 439718 53930 439954
rect 54166 439718 54250 439954
rect 54486 439718 54570 439954
rect 54806 439718 73930 439954
rect 74166 439718 74250 439954
rect 74486 439718 74570 439954
rect 74806 439718 93930 439954
rect 94166 439718 94250 439954
rect 94486 439718 94570 439954
rect 94806 439718 113930 439954
rect 114166 439718 114250 439954
rect 114486 439718 114570 439954
rect 114806 439718 133930 439954
rect 134166 439718 134250 439954
rect 134486 439718 134570 439954
rect 134806 439718 153930 439954
rect 154166 439718 154250 439954
rect 154486 439718 154570 439954
rect 154806 439718 173930 439954
rect 174166 439718 174250 439954
rect 174486 439718 174570 439954
rect 174806 439718 193930 439954
rect 194166 439718 194250 439954
rect 194486 439718 194570 439954
rect 194806 439718 213930 439954
rect 214166 439718 214250 439954
rect 214486 439718 214570 439954
rect 214806 439718 233930 439954
rect 234166 439718 234250 439954
rect 234486 439718 234570 439954
rect 234806 439718 253930 439954
rect 254166 439718 254250 439954
rect 254486 439718 254570 439954
rect 254806 439718 273930 439954
rect 274166 439718 274250 439954
rect 274486 439718 274570 439954
rect 274806 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 313930 439954
rect 314166 439718 314250 439954
rect 314486 439718 314570 439954
rect 314806 439718 333930 439954
rect 334166 439718 334250 439954
rect 334486 439718 334570 439954
rect 334806 439718 353930 439954
rect 354166 439718 354250 439954
rect 354486 439718 354570 439954
rect 354806 439718 373930 439954
rect 374166 439718 374250 439954
rect 374486 439718 374570 439954
rect 374806 439718 393930 439954
rect 394166 439718 394250 439954
rect 394486 439718 394570 439954
rect 394806 439718 413930 439954
rect 414166 439718 414250 439954
rect 414486 439718 414570 439954
rect 414806 439718 433930 439954
rect 434166 439718 434250 439954
rect 434486 439718 434570 439954
rect 434806 439718 453930 439954
rect 454166 439718 454250 439954
rect 454486 439718 454570 439954
rect 454806 439718 473930 439954
rect 474166 439718 474250 439954
rect 474486 439718 474570 439954
rect 474806 439718 493930 439954
rect 494166 439718 494250 439954
rect 494486 439718 494570 439954
rect 494806 439718 513930 439954
rect 514166 439718 514250 439954
rect 514486 439718 514570 439954
rect 514806 439718 533930 439954
rect 534166 439718 534250 439954
rect 534486 439718 534570 439954
rect 534806 439718 553930 439954
rect 554166 439718 554250 439954
rect 554486 439718 554570 439954
rect 554806 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 33930 439634
rect 34166 439398 34250 439634
rect 34486 439398 34570 439634
rect 34806 439398 53930 439634
rect 54166 439398 54250 439634
rect 54486 439398 54570 439634
rect 54806 439398 73930 439634
rect 74166 439398 74250 439634
rect 74486 439398 74570 439634
rect 74806 439398 93930 439634
rect 94166 439398 94250 439634
rect 94486 439398 94570 439634
rect 94806 439398 113930 439634
rect 114166 439398 114250 439634
rect 114486 439398 114570 439634
rect 114806 439398 133930 439634
rect 134166 439398 134250 439634
rect 134486 439398 134570 439634
rect 134806 439398 153930 439634
rect 154166 439398 154250 439634
rect 154486 439398 154570 439634
rect 154806 439398 173930 439634
rect 174166 439398 174250 439634
rect 174486 439398 174570 439634
rect 174806 439398 193930 439634
rect 194166 439398 194250 439634
rect 194486 439398 194570 439634
rect 194806 439398 213930 439634
rect 214166 439398 214250 439634
rect 214486 439398 214570 439634
rect 214806 439398 233930 439634
rect 234166 439398 234250 439634
rect 234486 439398 234570 439634
rect 234806 439398 253930 439634
rect 254166 439398 254250 439634
rect 254486 439398 254570 439634
rect 254806 439398 273930 439634
rect 274166 439398 274250 439634
rect 274486 439398 274570 439634
rect 274806 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 313930 439634
rect 314166 439398 314250 439634
rect 314486 439398 314570 439634
rect 314806 439398 333930 439634
rect 334166 439398 334250 439634
rect 334486 439398 334570 439634
rect 334806 439398 353930 439634
rect 354166 439398 354250 439634
rect 354486 439398 354570 439634
rect 354806 439398 373930 439634
rect 374166 439398 374250 439634
rect 374486 439398 374570 439634
rect 374806 439398 393930 439634
rect 394166 439398 394250 439634
rect 394486 439398 394570 439634
rect 394806 439398 413930 439634
rect 414166 439398 414250 439634
rect 414486 439398 414570 439634
rect 414806 439398 433930 439634
rect 434166 439398 434250 439634
rect 434486 439398 434570 439634
rect 434806 439398 453930 439634
rect 454166 439398 454250 439634
rect 454486 439398 454570 439634
rect 454806 439398 473930 439634
rect 474166 439398 474250 439634
rect 474486 439398 474570 439634
rect 474806 439398 493930 439634
rect 494166 439398 494250 439634
rect 494486 439398 494570 439634
rect 494806 439398 513930 439634
rect 514166 439398 514250 439634
rect 514486 439398 514570 439634
rect 514806 439398 533930 439634
rect 534166 439398 534250 439634
rect 534486 439398 534570 439634
rect 534806 439398 553930 439634
rect 554166 439398 554250 439634
rect 554486 439398 554570 439634
rect 554806 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 23930 435454
rect 24166 435218 24250 435454
rect 24486 435218 24570 435454
rect 24806 435218 43930 435454
rect 44166 435218 44250 435454
rect 44486 435218 44570 435454
rect 44806 435218 63930 435454
rect 64166 435218 64250 435454
rect 64486 435218 64570 435454
rect 64806 435218 83930 435454
rect 84166 435218 84250 435454
rect 84486 435218 84570 435454
rect 84806 435218 103930 435454
rect 104166 435218 104250 435454
rect 104486 435218 104570 435454
rect 104806 435218 123930 435454
rect 124166 435218 124250 435454
rect 124486 435218 124570 435454
rect 124806 435218 143930 435454
rect 144166 435218 144250 435454
rect 144486 435218 144570 435454
rect 144806 435218 163930 435454
rect 164166 435218 164250 435454
rect 164486 435218 164570 435454
rect 164806 435218 183930 435454
rect 184166 435218 184250 435454
rect 184486 435218 184570 435454
rect 184806 435218 203930 435454
rect 204166 435218 204250 435454
rect 204486 435218 204570 435454
rect 204806 435218 223930 435454
rect 224166 435218 224250 435454
rect 224486 435218 224570 435454
rect 224806 435218 243930 435454
rect 244166 435218 244250 435454
rect 244486 435218 244570 435454
rect 244806 435218 263930 435454
rect 264166 435218 264250 435454
rect 264486 435218 264570 435454
rect 264806 435218 283930 435454
rect 284166 435218 284250 435454
rect 284486 435218 284570 435454
rect 284806 435218 303930 435454
rect 304166 435218 304250 435454
rect 304486 435218 304570 435454
rect 304806 435218 323930 435454
rect 324166 435218 324250 435454
rect 324486 435218 324570 435454
rect 324806 435218 343930 435454
rect 344166 435218 344250 435454
rect 344486 435218 344570 435454
rect 344806 435218 363930 435454
rect 364166 435218 364250 435454
rect 364486 435218 364570 435454
rect 364806 435218 383930 435454
rect 384166 435218 384250 435454
rect 384486 435218 384570 435454
rect 384806 435218 403930 435454
rect 404166 435218 404250 435454
rect 404486 435218 404570 435454
rect 404806 435218 423930 435454
rect 424166 435218 424250 435454
rect 424486 435218 424570 435454
rect 424806 435218 443930 435454
rect 444166 435218 444250 435454
rect 444486 435218 444570 435454
rect 444806 435218 463930 435454
rect 464166 435218 464250 435454
rect 464486 435218 464570 435454
rect 464806 435218 483930 435454
rect 484166 435218 484250 435454
rect 484486 435218 484570 435454
rect 484806 435218 503930 435454
rect 504166 435218 504250 435454
rect 504486 435218 504570 435454
rect 504806 435218 523930 435454
rect 524166 435218 524250 435454
rect 524486 435218 524570 435454
rect 524806 435218 543930 435454
rect 544166 435218 544250 435454
rect 544486 435218 544570 435454
rect 544806 435218 563930 435454
rect 564166 435218 564250 435454
rect 564486 435218 564570 435454
rect 564806 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 23930 435134
rect 24166 434898 24250 435134
rect 24486 434898 24570 435134
rect 24806 434898 43930 435134
rect 44166 434898 44250 435134
rect 44486 434898 44570 435134
rect 44806 434898 63930 435134
rect 64166 434898 64250 435134
rect 64486 434898 64570 435134
rect 64806 434898 83930 435134
rect 84166 434898 84250 435134
rect 84486 434898 84570 435134
rect 84806 434898 103930 435134
rect 104166 434898 104250 435134
rect 104486 434898 104570 435134
rect 104806 434898 123930 435134
rect 124166 434898 124250 435134
rect 124486 434898 124570 435134
rect 124806 434898 143930 435134
rect 144166 434898 144250 435134
rect 144486 434898 144570 435134
rect 144806 434898 163930 435134
rect 164166 434898 164250 435134
rect 164486 434898 164570 435134
rect 164806 434898 183930 435134
rect 184166 434898 184250 435134
rect 184486 434898 184570 435134
rect 184806 434898 203930 435134
rect 204166 434898 204250 435134
rect 204486 434898 204570 435134
rect 204806 434898 223930 435134
rect 224166 434898 224250 435134
rect 224486 434898 224570 435134
rect 224806 434898 243930 435134
rect 244166 434898 244250 435134
rect 244486 434898 244570 435134
rect 244806 434898 263930 435134
rect 264166 434898 264250 435134
rect 264486 434898 264570 435134
rect 264806 434898 283930 435134
rect 284166 434898 284250 435134
rect 284486 434898 284570 435134
rect 284806 434898 303930 435134
rect 304166 434898 304250 435134
rect 304486 434898 304570 435134
rect 304806 434898 323930 435134
rect 324166 434898 324250 435134
rect 324486 434898 324570 435134
rect 324806 434898 343930 435134
rect 344166 434898 344250 435134
rect 344486 434898 344570 435134
rect 344806 434898 363930 435134
rect 364166 434898 364250 435134
rect 364486 434898 364570 435134
rect 364806 434898 383930 435134
rect 384166 434898 384250 435134
rect 384486 434898 384570 435134
rect 384806 434898 403930 435134
rect 404166 434898 404250 435134
rect 404486 434898 404570 435134
rect 404806 434898 423930 435134
rect 424166 434898 424250 435134
rect 424486 434898 424570 435134
rect 424806 434898 443930 435134
rect 444166 434898 444250 435134
rect 444486 434898 444570 435134
rect 444806 434898 463930 435134
rect 464166 434898 464250 435134
rect 464486 434898 464570 435134
rect 464806 434898 483930 435134
rect 484166 434898 484250 435134
rect 484486 434898 484570 435134
rect 484806 434898 503930 435134
rect 504166 434898 504250 435134
rect 504486 434898 504570 435134
rect 504806 434898 523930 435134
rect 524166 434898 524250 435134
rect 524486 434898 524570 435134
rect 524806 434898 543930 435134
rect 544166 434898 544250 435134
rect 544486 434898 544570 435134
rect 544806 434898 563930 435134
rect 564166 434898 564250 435134
rect 564486 434898 564570 435134
rect 564806 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 33930 403954
rect 34166 403718 34250 403954
rect 34486 403718 34570 403954
rect 34806 403718 53930 403954
rect 54166 403718 54250 403954
rect 54486 403718 54570 403954
rect 54806 403718 73930 403954
rect 74166 403718 74250 403954
rect 74486 403718 74570 403954
rect 74806 403718 93930 403954
rect 94166 403718 94250 403954
rect 94486 403718 94570 403954
rect 94806 403718 113930 403954
rect 114166 403718 114250 403954
rect 114486 403718 114570 403954
rect 114806 403718 133930 403954
rect 134166 403718 134250 403954
rect 134486 403718 134570 403954
rect 134806 403718 153930 403954
rect 154166 403718 154250 403954
rect 154486 403718 154570 403954
rect 154806 403718 173930 403954
rect 174166 403718 174250 403954
rect 174486 403718 174570 403954
rect 174806 403718 193930 403954
rect 194166 403718 194250 403954
rect 194486 403718 194570 403954
rect 194806 403718 213930 403954
rect 214166 403718 214250 403954
rect 214486 403718 214570 403954
rect 214806 403718 233930 403954
rect 234166 403718 234250 403954
rect 234486 403718 234570 403954
rect 234806 403718 253930 403954
rect 254166 403718 254250 403954
rect 254486 403718 254570 403954
rect 254806 403718 273930 403954
rect 274166 403718 274250 403954
rect 274486 403718 274570 403954
rect 274806 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 313930 403954
rect 314166 403718 314250 403954
rect 314486 403718 314570 403954
rect 314806 403718 333930 403954
rect 334166 403718 334250 403954
rect 334486 403718 334570 403954
rect 334806 403718 353930 403954
rect 354166 403718 354250 403954
rect 354486 403718 354570 403954
rect 354806 403718 373930 403954
rect 374166 403718 374250 403954
rect 374486 403718 374570 403954
rect 374806 403718 393930 403954
rect 394166 403718 394250 403954
rect 394486 403718 394570 403954
rect 394806 403718 413930 403954
rect 414166 403718 414250 403954
rect 414486 403718 414570 403954
rect 414806 403718 433930 403954
rect 434166 403718 434250 403954
rect 434486 403718 434570 403954
rect 434806 403718 453930 403954
rect 454166 403718 454250 403954
rect 454486 403718 454570 403954
rect 454806 403718 473930 403954
rect 474166 403718 474250 403954
rect 474486 403718 474570 403954
rect 474806 403718 493930 403954
rect 494166 403718 494250 403954
rect 494486 403718 494570 403954
rect 494806 403718 513930 403954
rect 514166 403718 514250 403954
rect 514486 403718 514570 403954
rect 514806 403718 533930 403954
rect 534166 403718 534250 403954
rect 534486 403718 534570 403954
rect 534806 403718 553930 403954
rect 554166 403718 554250 403954
rect 554486 403718 554570 403954
rect 554806 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 33930 403634
rect 34166 403398 34250 403634
rect 34486 403398 34570 403634
rect 34806 403398 53930 403634
rect 54166 403398 54250 403634
rect 54486 403398 54570 403634
rect 54806 403398 73930 403634
rect 74166 403398 74250 403634
rect 74486 403398 74570 403634
rect 74806 403398 93930 403634
rect 94166 403398 94250 403634
rect 94486 403398 94570 403634
rect 94806 403398 113930 403634
rect 114166 403398 114250 403634
rect 114486 403398 114570 403634
rect 114806 403398 133930 403634
rect 134166 403398 134250 403634
rect 134486 403398 134570 403634
rect 134806 403398 153930 403634
rect 154166 403398 154250 403634
rect 154486 403398 154570 403634
rect 154806 403398 173930 403634
rect 174166 403398 174250 403634
rect 174486 403398 174570 403634
rect 174806 403398 193930 403634
rect 194166 403398 194250 403634
rect 194486 403398 194570 403634
rect 194806 403398 213930 403634
rect 214166 403398 214250 403634
rect 214486 403398 214570 403634
rect 214806 403398 233930 403634
rect 234166 403398 234250 403634
rect 234486 403398 234570 403634
rect 234806 403398 253930 403634
rect 254166 403398 254250 403634
rect 254486 403398 254570 403634
rect 254806 403398 273930 403634
rect 274166 403398 274250 403634
rect 274486 403398 274570 403634
rect 274806 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 313930 403634
rect 314166 403398 314250 403634
rect 314486 403398 314570 403634
rect 314806 403398 333930 403634
rect 334166 403398 334250 403634
rect 334486 403398 334570 403634
rect 334806 403398 353930 403634
rect 354166 403398 354250 403634
rect 354486 403398 354570 403634
rect 354806 403398 373930 403634
rect 374166 403398 374250 403634
rect 374486 403398 374570 403634
rect 374806 403398 393930 403634
rect 394166 403398 394250 403634
rect 394486 403398 394570 403634
rect 394806 403398 413930 403634
rect 414166 403398 414250 403634
rect 414486 403398 414570 403634
rect 414806 403398 433930 403634
rect 434166 403398 434250 403634
rect 434486 403398 434570 403634
rect 434806 403398 453930 403634
rect 454166 403398 454250 403634
rect 454486 403398 454570 403634
rect 454806 403398 473930 403634
rect 474166 403398 474250 403634
rect 474486 403398 474570 403634
rect 474806 403398 493930 403634
rect 494166 403398 494250 403634
rect 494486 403398 494570 403634
rect 494806 403398 513930 403634
rect 514166 403398 514250 403634
rect 514486 403398 514570 403634
rect 514806 403398 533930 403634
rect 534166 403398 534250 403634
rect 534486 403398 534570 403634
rect 534806 403398 553930 403634
rect 554166 403398 554250 403634
rect 554486 403398 554570 403634
rect 554806 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 23930 399454
rect 24166 399218 24250 399454
rect 24486 399218 24570 399454
rect 24806 399218 43930 399454
rect 44166 399218 44250 399454
rect 44486 399218 44570 399454
rect 44806 399218 63930 399454
rect 64166 399218 64250 399454
rect 64486 399218 64570 399454
rect 64806 399218 83930 399454
rect 84166 399218 84250 399454
rect 84486 399218 84570 399454
rect 84806 399218 103930 399454
rect 104166 399218 104250 399454
rect 104486 399218 104570 399454
rect 104806 399218 123930 399454
rect 124166 399218 124250 399454
rect 124486 399218 124570 399454
rect 124806 399218 143930 399454
rect 144166 399218 144250 399454
rect 144486 399218 144570 399454
rect 144806 399218 163930 399454
rect 164166 399218 164250 399454
rect 164486 399218 164570 399454
rect 164806 399218 183930 399454
rect 184166 399218 184250 399454
rect 184486 399218 184570 399454
rect 184806 399218 203930 399454
rect 204166 399218 204250 399454
rect 204486 399218 204570 399454
rect 204806 399218 223930 399454
rect 224166 399218 224250 399454
rect 224486 399218 224570 399454
rect 224806 399218 243930 399454
rect 244166 399218 244250 399454
rect 244486 399218 244570 399454
rect 244806 399218 263930 399454
rect 264166 399218 264250 399454
rect 264486 399218 264570 399454
rect 264806 399218 283930 399454
rect 284166 399218 284250 399454
rect 284486 399218 284570 399454
rect 284806 399218 303930 399454
rect 304166 399218 304250 399454
rect 304486 399218 304570 399454
rect 304806 399218 323930 399454
rect 324166 399218 324250 399454
rect 324486 399218 324570 399454
rect 324806 399218 343930 399454
rect 344166 399218 344250 399454
rect 344486 399218 344570 399454
rect 344806 399218 363930 399454
rect 364166 399218 364250 399454
rect 364486 399218 364570 399454
rect 364806 399218 383930 399454
rect 384166 399218 384250 399454
rect 384486 399218 384570 399454
rect 384806 399218 403930 399454
rect 404166 399218 404250 399454
rect 404486 399218 404570 399454
rect 404806 399218 423930 399454
rect 424166 399218 424250 399454
rect 424486 399218 424570 399454
rect 424806 399218 443930 399454
rect 444166 399218 444250 399454
rect 444486 399218 444570 399454
rect 444806 399218 463930 399454
rect 464166 399218 464250 399454
rect 464486 399218 464570 399454
rect 464806 399218 483930 399454
rect 484166 399218 484250 399454
rect 484486 399218 484570 399454
rect 484806 399218 503930 399454
rect 504166 399218 504250 399454
rect 504486 399218 504570 399454
rect 504806 399218 523930 399454
rect 524166 399218 524250 399454
rect 524486 399218 524570 399454
rect 524806 399218 543930 399454
rect 544166 399218 544250 399454
rect 544486 399218 544570 399454
rect 544806 399218 563930 399454
rect 564166 399218 564250 399454
rect 564486 399218 564570 399454
rect 564806 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 23930 399134
rect 24166 398898 24250 399134
rect 24486 398898 24570 399134
rect 24806 398898 43930 399134
rect 44166 398898 44250 399134
rect 44486 398898 44570 399134
rect 44806 398898 63930 399134
rect 64166 398898 64250 399134
rect 64486 398898 64570 399134
rect 64806 398898 83930 399134
rect 84166 398898 84250 399134
rect 84486 398898 84570 399134
rect 84806 398898 103930 399134
rect 104166 398898 104250 399134
rect 104486 398898 104570 399134
rect 104806 398898 123930 399134
rect 124166 398898 124250 399134
rect 124486 398898 124570 399134
rect 124806 398898 143930 399134
rect 144166 398898 144250 399134
rect 144486 398898 144570 399134
rect 144806 398898 163930 399134
rect 164166 398898 164250 399134
rect 164486 398898 164570 399134
rect 164806 398898 183930 399134
rect 184166 398898 184250 399134
rect 184486 398898 184570 399134
rect 184806 398898 203930 399134
rect 204166 398898 204250 399134
rect 204486 398898 204570 399134
rect 204806 398898 223930 399134
rect 224166 398898 224250 399134
rect 224486 398898 224570 399134
rect 224806 398898 243930 399134
rect 244166 398898 244250 399134
rect 244486 398898 244570 399134
rect 244806 398898 263930 399134
rect 264166 398898 264250 399134
rect 264486 398898 264570 399134
rect 264806 398898 283930 399134
rect 284166 398898 284250 399134
rect 284486 398898 284570 399134
rect 284806 398898 303930 399134
rect 304166 398898 304250 399134
rect 304486 398898 304570 399134
rect 304806 398898 323930 399134
rect 324166 398898 324250 399134
rect 324486 398898 324570 399134
rect 324806 398898 343930 399134
rect 344166 398898 344250 399134
rect 344486 398898 344570 399134
rect 344806 398898 363930 399134
rect 364166 398898 364250 399134
rect 364486 398898 364570 399134
rect 364806 398898 383930 399134
rect 384166 398898 384250 399134
rect 384486 398898 384570 399134
rect 384806 398898 403930 399134
rect 404166 398898 404250 399134
rect 404486 398898 404570 399134
rect 404806 398898 423930 399134
rect 424166 398898 424250 399134
rect 424486 398898 424570 399134
rect 424806 398898 443930 399134
rect 444166 398898 444250 399134
rect 444486 398898 444570 399134
rect 444806 398898 463930 399134
rect 464166 398898 464250 399134
rect 464486 398898 464570 399134
rect 464806 398898 483930 399134
rect 484166 398898 484250 399134
rect 484486 398898 484570 399134
rect 484806 398898 503930 399134
rect 504166 398898 504250 399134
rect 504486 398898 504570 399134
rect 504806 398898 523930 399134
rect 524166 398898 524250 399134
rect 524486 398898 524570 399134
rect 524806 398898 543930 399134
rect 544166 398898 544250 399134
rect 544486 398898 544570 399134
rect 544806 398898 563930 399134
rect 564166 398898 564250 399134
rect 564486 398898 564570 399134
rect 564806 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 33930 367954
rect 34166 367718 34250 367954
rect 34486 367718 34570 367954
rect 34806 367718 53930 367954
rect 54166 367718 54250 367954
rect 54486 367718 54570 367954
rect 54806 367718 73930 367954
rect 74166 367718 74250 367954
rect 74486 367718 74570 367954
rect 74806 367718 93930 367954
rect 94166 367718 94250 367954
rect 94486 367718 94570 367954
rect 94806 367718 113930 367954
rect 114166 367718 114250 367954
rect 114486 367718 114570 367954
rect 114806 367718 133930 367954
rect 134166 367718 134250 367954
rect 134486 367718 134570 367954
rect 134806 367718 153930 367954
rect 154166 367718 154250 367954
rect 154486 367718 154570 367954
rect 154806 367718 173930 367954
rect 174166 367718 174250 367954
rect 174486 367718 174570 367954
rect 174806 367718 193930 367954
rect 194166 367718 194250 367954
rect 194486 367718 194570 367954
rect 194806 367718 213930 367954
rect 214166 367718 214250 367954
rect 214486 367718 214570 367954
rect 214806 367718 233930 367954
rect 234166 367718 234250 367954
rect 234486 367718 234570 367954
rect 234806 367718 253930 367954
rect 254166 367718 254250 367954
rect 254486 367718 254570 367954
rect 254806 367718 273930 367954
rect 274166 367718 274250 367954
rect 274486 367718 274570 367954
rect 274806 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 313930 367954
rect 314166 367718 314250 367954
rect 314486 367718 314570 367954
rect 314806 367718 333930 367954
rect 334166 367718 334250 367954
rect 334486 367718 334570 367954
rect 334806 367718 353930 367954
rect 354166 367718 354250 367954
rect 354486 367718 354570 367954
rect 354806 367718 373930 367954
rect 374166 367718 374250 367954
rect 374486 367718 374570 367954
rect 374806 367718 393930 367954
rect 394166 367718 394250 367954
rect 394486 367718 394570 367954
rect 394806 367718 413930 367954
rect 414166 367718 414250 367954
rect 414486 367718 414570 367954
rect 414806 367718 433930 367954
rect 434166 367718 434250 367954
rect 434486 367718 434570 367954
rect 434806 367718 453930 367954
rect 454166 367718 454250 367954
rect 454486 367718 454570 367954
rect 454806 367718 473930 367954
rect 474166 367718 474250 367954
rect 474486 367718 474570 367954
rect 474806 367718 493930 367954
rect 494166 367718 494250 367954
rect 494486 367718 494570 367954
rect 494806 367718 513930 367954
rect 514166 367718 514250 367954
rect 514486 367718 514570 367954
rect 514806 367718 533930 367954
rect 534166 367718 534250 367954
rect 534486 367718 534570 367954
rect 534806 367718 553930 367954
rect 554166 367718 554250 367954
rect 554486 367718 554570 367954
rect 554806 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 33930 367634
rect 34166 367398 34250 367634
rect 34486 367398 34570 367634
rect 34806 367398 53930 367634
rect 54166 367398 54250 367634
rect 54486 367398 54570 367634
rect 54806 367398 73930 367634
rect 74166 367398 74250 367634
rect 74486 367398 74570 367634
rect 74806 367398 93930 367634
rect 94166 367398 94250 367634
rect 94486 367398 94570 367634
rect 94806 367398 113930 367634
rect 114166 367398 114250 367634
rect 114486 367398 114570 367634
rect 114806 367398 133930 367634
rect 134166 367398 134250 367634
rect 134486 367398 134570 367634
rect 134806 367398 153930 367634
rect 154166 367398 154250 367634
rect 154486 367398 154570 367634
rect 154806 367398 173930 367634
rect 174166 367398 174250 367634
rect 174486 367398 174570 367634
rect 174806 367398 193930 367634
rect 194166 367398 194250 367634
rect 194486 367398 194570 367634
rect 194806 367398 213930 367634
rect 214166 367398 214250 367634
rect 214486 367398 214570 367634
rect 214806 367398 233930 367634
rect 234166 367398 234250 367634
rect 234486 367398 234570 367634
rect 234806 367398 253930 367634
rect 254166 367398 254250 367634
rect 254486 367398 254570 367634
rect 254806 367398 273930 367634
rect 274166 367398 274250 367634
rect 274486 367398 274570 367634
rect 274806 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 313930 367634
rect 314166 367398 314250 367634
rect 314486 367398 314570 367634
rect 314806 367398 333930 367634
rect 334166 367398 334250 367634
rect 334486 367398 334570 367634
rect 334806 367398 353930 367634
rect 354166 367398 354250 367634
rect 354486 367398 354570 367634
rect 354806 367398 373930 367634
rect 374166 367398 374250 367634
rect 374486 367398 374570 367634
rect 374806 367398 393930 367634
rect 394166 367398 394250 367634
rect 394486 367398 394570 367634
rect 394806 367398 413930 367634
rect 414166 367398 414250 367634
rect 414486 367398 414570 367634
rect 414806 367398 433930 367634
rect 434166 367398 434250 367634
rect 434486 367398 434570 367634
rect 434806 367398 453930 367634
rect 454166 367398 454250 367634
rect 454486 367398 454570 367634
rect 454806 367398 473930 367634
rect 474166 367398 474250 367634
rect 474486 367398 474570 367634
rect 474806 367398 493930 367634
rect 494166 367398 494250 367634
rect 494486 367398 494570 367634
rect 494806 367398 513930 367634
rect 514166 367398 514250 367634
rect 514486 367398 514570 367634
rect 514806 367398 533930 367634
rect 534166 367398 534250 367634
rect 534486 367398 534570 367634
rect 534806 367398 553930 367634
rect 554166 367398 554250 367634
rect 554486 367398 554570 367634
rect 554806 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 23930 363454
rect 24166 363218 24250 363454
rect 24486 363218 24570 363454
rect 24806 363218 43930 363454
rect 44166 363218 44250 363454
rect 44486 363218 44570 363454
rect 44806 363218 63930 363454
rect 64166 363218 64250 363454
rect 64486 363218 64570 363454
rect 64806 363218 83930 363454
rect 84166 363218 84250 363454
rect 84486 363218 84570 363454
rect 84806 363218 103930 363454
rect 104166 363218 104250 363454
rect 104486 363218 104570 363454
rect 104806 363218 123930 363454
rect 124166 363218 124250 363454
rect 124486 363218 124570 363454
rect 124806 363218 143930 363454
rect 144166 363218 144250 363454
rect 144486 363218 144570 363454
rect 144806 363218 163930 363454
rect 164166 363218 164250 363454
rect 164486 363218 164570 363454
rect 164806 363218 183930 363454
rect 184166 363218 184250 363454
rect 184486 363218 184570 363454
rect 184806 363218 203930 363454
rect 204166 363218 204250 363454
rect 204486 363218 204570 363454
rect 204806 363218 223930 363454
rect 224166 363218 224250 363454
rect 224486 363218 224570 363454
rect 224806 363218 243930 363454
rect 244166 363218 244250 363454
rect 244486 363218 244570 363454
rect 244806 363218 263930 363454
rect 264166 363218 264250 363454
rect 264486 363218 264570 363454
rect 264806 363218 283930 363454
rect 284166 363218 284250 363454
rect 284486 363218 284570 363454
rect 284806 363218 303930 363454
rect 304166 363218 304250 363454
rect 304486 363218 304570 363454
rect 304806 363218 323930 363454
rect 324166 363218 324250 363454
rect 324486 363218 324570 363454
rect 324806 363218 343930 363454
rect 344166 363218 344250 363454
rect 344486 363218 344570 363454
rect 344806 363218 363930 363454
rect 364166 363218 364250 363454
rect 364486 363218 364570 363454
rect 364806 363218 383930 363454
rect 384166 363218 384250 363454
rect 384486 363218 384570 363454
rect 384806 363218 403930 363454
rect 404166 363218 404250 363454
rect 404486 363218 404570 363454
rect 404806 363218 423930 363454
rect 424166 363218 424250 363454
rect 424486 363218 424570 363454
rect 424806 363218 443930 363454
rect 444166 363218 444250 363454
rect 444486 363218 444570 363454
rect 444806 363218 463930 363454
rect 464166 363218 464250 363454
rect 464486 363218 464570 363454
rect 464806 363218 483930 363454
rect 484166 363218 484250 363454
rect 484486 363218 484570 363454
rect 484806 363218 503930 363454
rect 504166 363218 504250 363454
rect 504486 363218 504570 363454
rect 504806 363218 523930 363454
rect 524166 363218 524250 363454
rect 524486 363218 524570 363454
rect 524806 363218 543930 363454
rect 544166 363218 544250 363454
rect 544486 363218 544570 363454
rect 544806 363218 563930 363454
rect 564166 363218 564250 363454
rect 564486 363218 564570 363454
rect 564806 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 23930 363134
rect 24166 362898 24250 363134
rect 24486 362898 24570 363134
rect 24806 362898 43930 363134
rect 44166 362898 44250 363134
rect 44486 362898 44570 363134
rect 44806 362898 63930 363134
rect 64166 362898 64250 363134
rect 64486 362898 64570 363134
rect 64806 362898 83930 363134
rect 84166 362898 84250 363134
rect 84486 362898 84570 363134
rect 84806 362898 103930 363134
rect 104166 362898 104250 363134
rect 104486 362898 104570 363134
rect 104806 362898 123930 363134
rect 124166 362898 124250 363134
rect 124486 362898 124570 363134
rect 124806 362898 143930 363134
rect 144166 362898 144250 363134
rect 144486 362898 144570 363134
rect 144806 362898 163930 363134
rect 164166 362898 164250 363134
rect 164486 362898 164570 363134
rect 164806 362898 183930 363134
rect 184166 362898 184250 363134
rect 184486 362898 184570 363134
rect 184806 362898 203930 363134
rect 204166 362898 204250 363134
rect 204486 362898 204570 363134
rect 204806 362898 223930 363134
rect 224166 362898 224250 363134
rect 224486 362898 224570 363134
rect 224806 362898 243930 363134
rect 244166 362898 244250 363134
rect 244486 362898 244570 363134
rect 244806 362898 263930 363134
rect 264166 362898 264250 363134
rect 264486 362898 264570 363134
rect 264806 362898 283930 363134
rect 284166 362898 284250 363134
rect 284486 362898 284570 363134
rect 284806 362898 303930 363134
rect 304166 362898 304250 363134
rect 304486 362898 304570 363134
rect 304806 362898 323930 363134
rect 324166 362898 324250 363134
rect 324486 362898 324570 363134
rect 324806 362898 343930 363134
rect 344166 362898 344250 363134
rect 344486 362898 344570 363134
rect 344806 362898 363930 363134
rect 364166 362898 364250 363134
rect 364486 362898 364570 363134
rect 364806 362898 383930 363134
rect 384166 362898 384250 363134
rect 384486 362898 384570 363134
rect 384806 362898 403930 363134
rect 404166 362898 404250 363134
rect 404486 362898 404570 363134
rect 404806 362898 423930 363134
rect 424166 362898 424250 363134
rect 424486 362898 424570 363134
rect 424806 362898 443930 363134
rect 444166 362898 444250 363134
rect 444486 362898 444570 363134
rect 444806 362898 463930 363134
rect 464166 362898 464250 363134
rect 464486 362898 464570 363134
rect 464806 362898 483930 363134
rect 484166 362898 484250 363134
rect 484486 362898 484570 363134
rect 484806 362898 503930 363134
rect 504166 362898 504250 363134
rect 504486 362898 504570 363134
rect 504806 362898 523930 363134
rect 524166 362898 524250 363134
rect 524486 362898 524570 363134
rect 524806 362898 543930 363134
rect 544166 362898 544250 363134
rect 544486 362898 544570 363134
rect 544806 362898 563930 363134
rect 564166 362898 564250 363134
rect 564486 362898 564570 363134
rect 564806 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 33930 295954
rect 34166 295718 34250 295954
rect 34486 295718 34570 295954
rect 34806 295718 53930 295954
rect 54166 295718 54250 295954
rect 54486 295718 54570 295954
rect 54806 295718 73930 295954
rect 74166 295718 74250 295954
rect 74486 295718 74570 295954
rect 74806 295718 93930 295954
rect 94166 295718 94250 295954
rect 94486 295718 94570 295954
rect 94806 295718 113930 295954
rect 114166 295718 114250 295954
rect 114486 295718 114570 295954
rect 114806 295718 133930 295954
rect 134166 295718 134250 295954
rect 134486 295718 134570 295954
rect 134806 295718 153930 295954
rect 154166 295718 154250 295954
rect 154486 295718 154570 295954
rect 154806 295718 173930 295954
rect 174166 295718 174250 295954
rect 174486 295718 174570 295954
rect 174806 295718 193930 295954
rect 194166 295718 194250 295954
rect 194486 295718 194570 295954
rect 194806 295718 213930 295954
rect 214166 295718 214250 295954
rect 214486 295718 214570 295954
rect 214806 295718 233930 295954
rect 234166 295718 234250 295954
rect 234486 295718 234570 295954
rect 234806 295718 253930 295954
rect 254166 295718 254250 295954
rect 254486 295718 254570 295954
rect 254806 295718 273930 295954
rect 274166 295718 274250 295954
rect 274486 295718 274570 295954
rect 274806 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 313930 295954
rect 314166 295718 314250 295954
rect 314486 295718 314570 295954
rect 314806 295718 333930 295954
rect 334166 295718 334250 295954
rect 334486 295718 334570 295954
rect 334806 295718 353930 295954
rect 354166 295718 354250 295954
rect 354486 295718 354570 295954
rect 354806 295718 373930 295954
rect 374166 295718 374250 295954
rect 374486 295718 374570 295954
rect 374806 295718 393930 295954
rect 394166 295718 394250 295954
rect 394486 295718 394570 295954
rect 394806 295718 413930 295954
rect 414166 295718 414250 295954
rect 414486 295718 414570 295954
rect 414806 295718 433930 295954
rect 434166 295718 434250 295954
rect 434486 295718 434570 295954
rect 434806 295718 453930 295954
rect 454166 295718 454250 295954
rect 454486 295718 454570 295954
rect 454806 295718 473930 295954
rect 474166 295718 474250 295954
rect 474486 295718 474570 295954
rect 474806 295718 493930 295954
rect 494166 295718 494250 295954
rect 494486 295718 494570 295954
rect 494806 295718 513930 295954
rect 514166 295718 514250 295954
rect 514486 295718 514570 295954
rect 514806 295718 533930 295954
rect 534166 295718 534250 295954
rect 534486 295718 534570 295954
rect 534806 295718 553930 295954
rect 554166 295718 554250 295954
rect 554486 295718 554570 295954
rect 554806 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 33930 295634
rect 34166 295398 34250 295634
rect 34486 295398 34570 295634
rect 34806 295398 53930 295634
rect 54166 295398 54250 295634
rect 54486 295398 54570 295634
rect 54806 295398 73930 295634
rect 74166 295398 74250 295634
rect 74486 295398 74570 295634
rect 74806 295398 93930 295634
rect 94166 295398 94250 295634
rect 94486 295398 94570 295634
rect 94806 295398 113930 295634
rect 114166 295398 114250 295634
rect 114486 295398 114570 295634
rect 114806 295398 133930 295634
rect 134166 295398 134250 295634
rect 134486 295398 134570 295634
rect 134806 295398 153930 295634
rect 154166 295398 154250 295634
rect 154486 295398 154570 295634
rect 154806 295398 173930 295634
rect 174166 295398 174250 295634
rect 174486 295398 174570 295634
rect 174806 295398 193930 295634
rect 194166 295398 194250 295634
rect 194486 295398 194570 295634
rect 194806 295398 213930 295634
rect 214166 295398 214250 295634
rect 214486 295398 214570 295634
rect 214806 295398 233930 295634
rect 234166 295398 234250 295634
rect 234486 295398 234570 295634
rect 234806 295398 253930 295634
rect 254166 295398 254250 295634
rect 254486 295398 254570 295634
rect 254806 295398 273930 295634
rect 274166 295398 274250 295634
rect 274486 295398 274570 295634
rect 274806 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 313930 295634
rect 314166 295398 314250 295634
rect 314486 295398 314570 295634
rect 314806 295398 333930 295634
rect 334166 295398 334250 295634
rect 334486 295398 334570 295634
rect 334806 295398 353930 295634
rect 354166 295398 354250 295634
rect 354486 295398 354570 295634
rect 354806 295398 373930 295634
rect 374166 295398 374250 295634
rect 374486 295398 374570 295634
rect 374806 295398 393930 295634
rect 394166 295398 394250 295634
rect 394486 295398 394570 295634
rect 394806 295398 413930 295634
rect 414166 295398 414250 295634
rect 414486 295398 414570 295634
rect 414806 295398 433930 295634
rect 434166 295398 434250 295634
rect 434486 295398 434570 295634
rect 434806 295398 453930 295634
rect 454166 295398 454250 295634
rect 454486 295398 454570 295634
rect 454806 295398 473930 295634
rect 474166 295398 474250 295634
rect 474486 295398 474570 295634
rect 474806 295398 493930 295634
rect 494166 295398 494250 295634
rect 494486 295398 494570 295634
rect 494806 295398 513930 295634
rect 514166 295398 514250 295634
rect 514486 295398 514570 295634
rect 514806 295398 533930 295634
rect 534166 295398 534250 295634
rect 534486 295398 534570 295634
rect 534806 295398 553930 295634
rect 554166 295398 554250 295634
rect 554486 295398 554570 295634
rect 554806 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 23930 291454
rect 24166 291218 24250 291454
rect 24486 291218 24570 291454
rect 24806 291218 43930 291454
rect 44166 291218 44250 291454
rect 44486 291218 44570 291454
rect 44806 291218 63930 291454
rect 64166 291218 64250 291454
rect 64486 291218 64570 291454
rect 64806 291218 83930 291454
rect 84166 291218 84250 291454
rect 84486 291218 84570 291454
rect 84806 291218 103930 291454
rect 104166 291218 104250 291454
rect 104486 291218 104570 291454
rect 104806 291218 123930 291454
rect 124166 291218 124250 291454
rect 124486 291218 124570 291454
rect 124806 291218 143930 291454
rect 144166 291218 144250 291454
rect 144486 291218 144570 291454
rect 144806 291218 163930 291454
rect 164166 291218 164250 291454
rect 164486 291218 164570 291454
rect 164806 291218 183930 291454
rect 184166 291218 184250 291454
rect 184486 291218 184570 291454
rect 184806 291218 203930 291454
rect 204166 291218 204250 291454
rect 204486 291218 204570 291454
rect 204806 291218 223930 291454
rect 224166 291218 224250 291454
rect 224486 291218 224570 291454
rect 224806 291218 243930 291454
rect 244166 291218 244250 291454
rect 244486 291218 244570 291454
rect 244806 291218 263930 291454
rect 264166 291218 264250 291454
rect 264486 291218 264570 291454
rect 264806 291218 283930 291454
rect 284166 291218 284250 291454
rect 284486 291218 284570 291454
rect 284806 291218 303930 291454
rect 304166 291218 304250 291454
rect 304486 291218 304570 291454
rect 304806 291218 323930 291454
rect 324166 291218 324250 291454
rect 324486 291218 324570 291454
rect 324806 291218 343930 291454
rect 344166 291218 344250 291454
rect 344486 291218 344570 291454
rect 344806 291218 363930 291454
rect 364166 291218 364250 291454
rect 364486 291218 364570 291454
rect 364806 291218 383930 291454
rect 384166 291218 384250 291454
rect 384486 291218 384570 291454
rect 384806 291218 403930 291454
rect 404166 291218 404250 291454
rect 404486 291218 404570 291454
rect 404806 291218 423930 291454
rect 424166 291218 424250 291454
rect 424486 291218 424570 291454
rect 424806 291218 443930 291454
rect 444166 291218 444250 291454
rect 444486 291218 444570 291454
rect 444806 291218 463930 291454
rect 464166 291218 464250 291454
rect 464486 291218 464570 291454
rect 464806 291218 483930 291454
rect 484166 291218 484250 291454
rect 484486 291218 484570 291454
rect 484806 291218 503930 291454
rect 504166 291218 504250 291454
rect 504486 291218 504570 291454
rect 504806 291218 523930 291454
rect 524166 291218 524250 291454
rect 524486 291218 524570 291454
rect 524806 291218 543930 291454
rect 544166 291218 544250 291454
rect 544486 291218 544570 291454
rect 544806 291218 563930 291454
rect 564166 291218 564250 291454
rect 564486 291218 564570 291454
rect 564806 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 23930 291134
rect 24166 290898 24250 291134
rect 24486 290898 24570 291134
rect 24806 290898 43930 291134
rect 44166 290898 44250 291134
rect 44486 290898 44570 291134
rect 44806 290898 63930 291134
rect 64166 290898 64250 291134
rect 64486 290898 64570 291134
rect 64806 290898 83930 291134
rect 84166 290898 84250 291134
rect 84486 290898 84570 291134
rect 84806 290898 103930 291134
rect 104166 290898 104250 291134
rect 104486 290898 104570 291134
rect 104806 290898 123930 291134
rect 124166 290898 124250 291134
rect 124486 290898 124570 291134
rect 124806 290898 143930 291134
rect 144166 290898 144250 291134
rect 144486 290898 144570 291134
rect 144806 290898 163930 291134
rect 164166 290898 164250 291134
rect 164486 290898 164570 291134
rect 164806 290898 183930 291134
rect 184166 290898 184250 291134
rect 184486 290898 184570 291134
rect 184806 290898 203930 291134
rect 204166 290898 204250 291134
rect 204486 290898 204570 291134
rect 204806 290898 223930 291134
rect 224166 290898 224250 291134
rect 224486 290898 224570 291134
rect 224806 290898 243930 291134
rect 244166 290898 244250 291134
rect 244486 290898 244570 291134
rect 244806 290898 263930 291134
rect 264166 290898 264250 291134
rect 264486 290898 264570 291134
rect 264806 290898 283930 291134
rect 284166 290898 284250 291134
rect 284486 290898 284570 291134
rect 284806 290898 303930 291134
rect 304166 290898 304250 291134
rect 304486 290898 304570 291134
rect 304806 290898 323930 291134
rect 324166 290898 324250 291134
rect 324486 290898 324570 291134
rect 324806 290898 343930 291134
rect 344166 290898 344250 291134
rect 344486 290898 344570 291134
rect 344806 290898 363930 291134
rect 364166 290898 364250 291134
rect 364486 290898 364570 291134
rect 364806 290898 383930 291134
rect 384166 290898 384250 291134
rect 384486 290898 384570 291134
rect 384806 290898 403930 291134
rect 404166 290898 404250 291134
rect 404486 290898 404570 291134
rect 404806 290898 423930 291134
rect 424166 290898 424250 291134
rect 424486 290898 424570 291134
rect 424806 290898 443930 291134
rect 444166 290898 444250 291134
rect 444486 290898 444570 291134
rect 444806 290898 463930 291134
rect 464166 290898 464250 291134
rect 464486 290898 464570 291134
rect 464806 290898 483930 291134
rect 484166 290898 484250 291134
rect 484486 290898 484570 291134
rect 484806 290898 503930 291134
rect 504166 290898 504250 291134
rect 504486 290898 504570 291134
rect 504806 290898 523930 291134
rect 524166 290898 524250 291134
rect 524486 290898 524570 291134
rect 524806 290898 543930 291134
rect 544166 290898 544250 291134
rect 544486 290898 544570 291134
rect 544806 290898 563930 291134
rect 564166 290898 564250 291134
rect 564486 290898 564570 291134
rect 564806 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 33930 259954
rect 34166 259718 34250 259954
rect 34486 259718 34570 259954
rect 34806 259718 53930 259954
rect 54166 259718 54250 259954
rect 54486 259718 54570 259954
rect 54806 259718 73930 259954
rect 74166 259718 74250 259954
rect 74486 259718 74570 259954
rect 74806 259718 93930 259954
rect 94166 259718 94250 259954
rect 94486 259718 94570 259954
rect 94806 259718 113930 259954
rect 114166 259718 114250 259954
rect 114486 259718 114570 259954
rect 114806 259718 133930 259954
rect 134166 259718 134250 259954
rect 134486 259718 134570 259954
rect 134806 259718 153930 259954
rect 154166 259718 154250 259954
rect 154486 259718 154570 259954
rect 154806 259718 173930 259954
rect 174166 259718 174250 259954
rect 174486 259718 174570 259954
rect 174806 259718 193930 259954
rect 194166 259718 194250 259954
rect 194486 259718 194570 259954
rect 194806 259718 213930 259954
rect 214166 259718 214250 259954
rect 214486 259718 214570 259954
rect 214806 259718 233930 259954
rect 234166 259718 234250 259954
rect 234486 259718 234570 259954
rect 234806 259718 253930 259954
rect 254166 259718 254250 259954
rect 254486 259718 254570 259954
rect 254806 259718 273930 259954
rect 274166 259718 274250 259954
rect 274486 259718 274570 259954
rect 274806 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 313930 259954
rect 314166 259718 314250 259954
rect 314486 259718 314570 259954
rect 314806 259718 333930 259954
rect 334166 259718 334250 259954
rect 334486 259718 334570 259954
rect 334806 259718 353930 259954
rect 354166 259718 354250 259954
rect 354486 259718 354570 259954
rect 354806 259718 373930 259954
rect 374166 259718 374250 259954
rect 374486 259718 374570 259954
rect 374806 259718 393930 259954
rect 394166 259718 394250 259954
rect 394486 259718 394570 259954
rect 394806 259718 413930 259954
rect 414166 259718 414250 259954
rect 414486 259718 414570 259954
rect 414806 259718 433930 259954
rect 434166 259718 434250 259954
rect 434486 259718 434570 259954
rect 434806 259718 453930 259954
rect 454166 259718 454250 259954
rect 454486 259718 454570 259954
rect 454806 259718 473930 259954
rect 474166 259718 474250 259954
rect 474486 259718 474570 259954
rect 474806 259718 493930 259954
rect 494166 259718 494250 259954
rect 494486 259718 494570 259954
rect 494806 259718 513930 259954
rect 514166 259718 514250 259954
rect 514486 259718 514570 259954
rect 514806 259718 533930 259954
rect 534166 259718 534250 259954
rect 534486 259718 534570 259954
rect 534806 259718 553930 259954
rect 554166 259718 554250 259954
rect 554486 259718 554570 259954
rect 554806 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 33930 259634
rect 34166 259398 34250 259634
rect 34486 259398 34570 259634
rect 34806 259398 53930 259634
rect 54166 259398 54250 259634
rect 54486 259398 54570 259634
rect 54806 259398 73930 259634
rect 74166 259398 74250 259634
rect 74486 259398 74570 259634
rect 74806 259398 93930 259634
rect 94166 259398 94250 259634
rect 94486 259398 94570 259634
rect 94806 259398 113930 259634
rect 114166 259398 114250 259634
rect 114486 259398 114570 259634
rect 114806 259398 133930 259634
rect 134166 259398 134250 259634
rect 134486 259398 134570 259634
rect 134806 259398 153930 259634
rect 154166 259398 154250 259634
rect 154486 259398 154570 259634
rect 154806 259398 173930 259634
rect 174166 259398 174250 259634
rect 174486 259398 174570 259634
rect 174806 259398 193930 259634
rect 194166 259398 194250 259634
rect 194486 259398 194570 259634
rect 194806 259398 213930 259634
rect 214166 259398 214250 259634
rect 214486 259398 214570 259634
rect 214806 259398 233930 259634
rect 234166 259398 234250 259634
rect 234486 259398 234570 259634
rect 234806 259398 253930 259634
rect 254166 259398 254250 259634
rect 254486 259398 254570 259634
rect 254806 259398 273930 259634
rect 274166 259398 274250 259634
rect 274486 259398 274570 259634
rect 274806 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 313930 259634
rect 314166 259398 314250 259634
rect 314486 259398 314570 259634
rect 314806 259398 333930 259634
rect 334166 259398 334250 259634
rect 334486 259398 334570 259634
rect 334806 259398 353930 259634
rect 354166 259398 354250 259634
rect 354486 259398 354570 259634
rect 354806 259398 373930 259634
rect 374166 259398 374250 259634
rect 374486 259398 374570 259634
rect 374806 259398 393930 259634
rect 394166 259398 394250 259634
rect 394486 259398 394570 259634
rect 394806 259398 413930 259634
rect 414166 259398 414250 259634
rect 414486 259398 414570 259634
rect 414806 259398 433930 259634
rect 434166 259398 434250 259634
rect 434486 259398 434570 259634
rect 434806 259398 453930 259634
rect 454166 259398 454250 259634
rect 454486 259398 454570 259634
rect 454806 259398 473930 259634
rect 474166 259398 474250 259634
rect 474486 259398 474570 259634
rect 474806 259398 493930 259634
rect 494166 259398 494250 259634
rect 494486 259398 494570 259634
rect 494806 259398 513930 259634
rect 514166 259398 514250 259634
rect 514486 259398 514570 259634
rect 514806 259398 533930 259634
rect 534166 259398 534250 259634
rect 534486 259398 534570 259634
rect 534806 259398 553930 259634
rect 554166 259398 554250 259634
rect 554486 259398 554570 259634
rect 554806 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 23930 255454
rect 24166 255218 24250 255454
rect 24486 255218 24570 255454
rect 24806 255218 43930 255454
rect 44166 255218 44250 255454
rect 44486 255218 44570 255454
rect 44806 255218 63930 255454
rect 64166 255218 64250 255454
rect 64486 255218 64570 255454
rect 64806 255218 83930 255454
rect 84166 255218 84250 255454
rect 84486 255218 84570 255454
rect 84806 255218 103930 255454
rect 104166 255218 104250 255454
rect 104486 255218 104570 255454
rect 104806 255218 123930 255454
rect 124166 255218 124250 255454
rect 124486 255218 124570 255454
rect 124806 255218 143930 255454
rect 144166 255218 144250 255454
rect 144486 255218 144570 255454
rect 144806 255218 163930 255454
rect 164166 255218 164250 255454
rect 164486 255218 164570 255454
rect 164806 255218 183930 255454
rect 184166 255218 184250 255454
rect 184486 255218 184570 255454
rect 184806 255218 203930 255454
rect 204166 255218 204250 255454
rect 204486 255218 204570 255454
rect 204806 255218 223930 255454
rect 224166 255218 224250 255454
rect 224486 255218 224570 255454
rect 224806 255218 243930 255454
rect 244166 255218 244250 255454
rect 244486 255218 244570 255454
rect 244806 255218 263930 255454
rect 264166 255218 264250 255454
rect 264486 255218 264570 255454
rect 264806 255218 283930 255454
rect 284166 255218 284250 255454
rect 284486 255218 284570 255454
rect 284806 255218 303930 255454
rect 304166 255218 304250 255454
rect 304486 255218 304570 255454
rect 304806 255218 323930 255454
rect 324166 255218 324250 255454
rect 324486 255218 324570 255454
rect 324806 255218 343930 255454
rect 344166 255218 344250 255454
rect 344486 255218 344570 255454
rect 344806 255218 363930 255454
rect 364166 255218 364250 255454
rect 364486 255218 364570 255454
rect 364806 255218 383930 255454
rect 384166 255218 384250 255454
rect 384486 255218 384570 255454
rect 384806 255218 403930 255454
rect 404166 255218 404250 255454
rect 404486 255218 404570 255454
rect 404806 255218 423930 255454
rect 424166 255218 424250 255454
rect 424486 255218 424570 255454
rect 424806 255218 443930 255454
rect 444166 255218 444250 255454
rect 444486 255218 444570 255454
rect 444806 255218 463930 255454
rect 464166 255218 464250 255454
rect 464486 255218 464570 255454
rect 464806 255218 483930 255454
rect 484166 255218 484250 255454
rect 484486 255218 484570 255454
rect 484806 255218 503930 255454
rect 504166 255218 504250 255454
rect 504486 255218 504570 255454
rect 504806 255218 523930 255454
rect 524166 255218 524250 255454
rect 524486 255218 524570 255454
rect 524806 255218 543930 255454
rect 544166 255218 544250 255454
rect 544486 255218 544570 255454
rect 544806 255218 563930 255454
rect 564166 255218 564250 255454
rect 564486 255218 564570 255454
rect 564806 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 23930 255134
rect 24166 254898 24250 255134
rect 24486 254898 24570 255134
rect 24806 254898 43930 255134
rect 44166 254898 44250 255134
rect 44486 254898 44570 255134
rect 44806 254898 63930 255134
rect 64166 254898 64250 255134
rect 64486 254898 64570 255134
rect 64806 254898 83930 255134
rect 84166 254898 84250 255134
rect 84486 254898 84570 255134
rect 84806 254898 103930 255134
rect 104166 254898 104250 255134
rect 104486 254898 104570 255134
rect 104806 254898 123930 255134
rect 124166 254898 124250 255134
rect 124486 254898 124570 255134
rect 124806 254898 143930 255134
rect 144166 254898 144250 255134
rect 144486 254898 144570 255134
rect 144806 254898 163930 255134
rect 164166 254898 164250 255134
rect 164486 254898 164570 255134
rect 164806 254898 183930 255134
rect 184166 254898 184250 255134
rect 184486 254898 184570 255134
rect 184806 254898 203930 255134
rect 204166 254898 204250 255134
rect 204486 254898 204570 255134
rect 204806 254898 223930 255134
rect 224166 254898 224250 255134
rect 224486 254898 224570 255134
rect 224806 254898 243930 255134
rect 244166 254898 244250 255134
rect 244486 254898 244570 255134
rect 244806 254898 263930 255134
rect 264166 254898 264250 255134
rect 264486 254898 264570 255134
rect 264806 254898 283930 255134
rect 284166 254898 284250 255134
rect 284486 254898 284570 255134
rect 284806 254898 303930 255134
rect 304166 254898 304250 255134
rect 304486 254898 304570 255134
rect 304806 254898 323930 255134
rect 324166 254898 324250 255134
rect 324486 254898 324570 255134
rect 324806 254898 343930 255134
rect 344166 254898 344250 255134
rect 344486 254898 344570 255134
rect 344806 254898 363930 255134
rect 364166 254898 364250 255134
rect 364486 254898 364570 255134
rect 364806 254898 383930 255134
rect 384166 254898 384250 255134
rect 384486 254898 384570 255134
rect 384806 254898 403930 255134
rect 404166 254898 404250 255134
rect 404486 254898 404570 255134
rect 404806 254898 423930 255134
rect 424166 254898 424250 255134
rect 424486 254898 424570 255134
rect 424806 254898 443930 255134
rect 444166 254898 444250 255134
rect 444486 254898 444570 255134
rect 444806 254898 463930 255134
rect 464166 254898 464250 255134
rect 464486 254898 464570 255134
rect 464806 254898 483930 255134
rect 484166 254898 484250 255134
rect 484486 254898 484570 255134
rect 484806 254898 503930 255134
rect 504166 254898 504250 255134
rect 504486 254898 504570 255134
rect 504806 254898 523930 255134
rect 524166 254898 524250 255134
rect 524486 254898 524570 255134
rect 524806 254898 543930 255134
rect 544166 254898 544250 255134
rect 544486 254898 544570 255134
rect 544806 254898 563930 255134
rect 564166 254898 564250 255134
rect 564486 254898 564570 255134
rect 564806 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 33930 223954
rect 34166 223718 34250 223954
rect 34486 223718 34570 223954
rect 34806 223718 53930 223954
rect 54166 223718 54250 223954
rect 54486 223718 54570 223954
rect 54806 223718 73930 223954
rect 74166 223718 74250 223954
rect 74486 223718 74570 223954
rect 74806 223718 93930 223954
rect 94166 223718 94250 223954
rect 94486 223718 94570 223954
rect 94806 223718 113930 223954
rect 114166 223718 114250 223954
rect 114486 223718 114570 223954
rect 114806 223718 133930 223954
rect 134166 223718 134250 223954
rect 134486 223718 134570 223954
rect 134806 223718 153930 223954
rect 154166 223718 154250 223954
rect 154486 223718 154570 223954
rect 154806 223718 173930 223954
rect 174166 223718 174250 223954
rect 174486 223718 174570 223954
rect 174806 223718 193930 223954
rect 194166 223718 194250 223954
rect 194486 223718 194570 223954
rect 194806 223718 213930 223954
rect 214166 223718 214250 223954
rect 214486 223718 214570 223954
rect 214806 223718 233930 223954
rect 234166 223718 234250 223954
rect 234486 223718 234570 223954
rect 234806 223718 253930 223954
rect 254166 223718 254250 223954
rect 254486 223718 254570 223954
rect 254806 223718 273930 223954
rect 274166 223718 274250 223954
rect 274486 223718 274570 223954
rect 274806 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 313930 223954
rect 314166 223718 314250 223954
rect 314486 223718 314570 223954
rect 314806 223718 333930 223954
rect 334166 223718 334250 223954
rect 334486 223718 334570 223954
rect 334806 223718 353930 223954
rect 354166 223718 354250 223954
rect 354486 223718 354570 223954
rect 354806 223718 373930 223954
rect 374166 223718 374250 223954
rect 374486 223718 374570 223954
rect 374806 223718 393930 223954
rect 394166 223718 394250 223954
rect 394486 223718 394570 223954
rect 394806 223718 413930 223954
rect 414166 223718 414250 223954
rect 414486 223718 414570 223954
rect 414806 223718 433930 223954
rect 434166 223718 434250 223954
rect 434486 223718 434570 223954
rect 434806 223718 453930 223954
rect 454166 223718 454250 223954
rect 454486 223718 454570 223954
rect 454806 223718 473930 223954
rect 474166 223718 474250 223954
rect 474486 223718 474570 223954
rect 474806 223718 493930 223954
rect 494166 223718 494250 223954
rect 494486 223718 494570 223954
rect 494806 223718 513930 223954
rect 514166 223718 514250 223954
rect 514486 223718 514570 223954
rect 514806 223718 533930 223954
rect 534166 223718 534250 223954
rect 534486 223718 534570 223954
rect 534806 223718 553930 223954
rect 554166 223718 554250 223954
rect 554486 223718 554570 223954
rect 554806 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 33930 223634
rect 34166 223398 34250 223634
rect 34486 223398 34570 223634
rect 34806 223398 53930 223634
rect 54166 223398 54250 223634
rect 54486 223398 54570 223634
rect 54806 223398 73930 223634
rect 74166 223398 74250 223634
rect 74486 223398 74570 223634
rect 74806 223398 93930 223634
rect 94166 223398 94250 223634
rect 94486 223398 94570 223634
rect 94806 223398 113930 223634
rect 114166 223398 114250 223634
rect 114486 223398 114570 223634
rect 114806 223398 133930 223634
rect 134166 223398 134250 223634
rect 134486 223398 134570 223634
rect 134806 223398 153930 223634
rect 154166 223398 154250 223634
rect 154486 223398 154570 223634
rect 154806 223398 173930 223634
rect 174166 223398 174250 223634
rect 174486 223398 174570 223634
rect 174806 223398 193930 223634
rect 194166 223398 194250 223634
rect 194486 223398 194570 223634
rect 194806 223398 213930 223634
rect 214166 223398 214250 223634
rect 214486 223398 214570 223634
rect 214806 223398 233930 223634
rect 234166 223398 234250 223634
rect 234486 223398 234570 223634
rect 234806 223398 253930 223634
rect 254166 223398 254250 223634
rect 254486 223398 254570 223634
rect 254806 223398 273930 223634
rect 274166 223398 274250 223634
rect 274486 223398 274570 223634
rect 274806 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 313930 223634
rect 314166 223398 314250 223634
rect 314486 223398 314570 223634
rect 314806 223398 333930 223634
rect 334166 223398 334250 223634
rect 334486 223398 334570 223634
rect 334806 223398 353930 223634
rect 354166 223398 354250 223634
rect 354486 223398 354570 223634
rect 354806 223398 373930 223634
rect 374166 223398 374250 223634
rect 374486 223398 374570 223634
rect 374806 223398 393930 223634
rect 394166 223398 394250 223634
rect 394486 223398 394570 223634
rect 394806 223398 413930 223634
rect 414166 223398 414250 223634
rect 414486 223398 414570 223634
rect 414806 223398 433930 223634
rect 434166 223398 434250 223634
rect 434486 223398 434570 223634
rect 434806 223398 453930 223634
rect 454166 223398 454250 223634
rect 454486 223398 454570 223634
rect 454806 223398 473930 223634
rect 474166 223398 474250 223634
rect 474486 223398 474570 223634
rect 474806 223398 493930 223634
rect 494166 223398 494250 223634
rect 494486 223398 494570 223634
rect 494806 223398 513930 223634
rect 514166 223398 514250 223634
rect 514486 223398 514570 223634
rect 514806 223398 533930 223634
rect 534166 223398 534250 223634
rect 534486 223398 534570 223634
rect 534806 223398 553930 223634
rect 554166 223398 554250 223634
rect 554486 223398 554570 223634
rect 554806 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 23930 219454
rect 24166 219218 24250 219454
rect 24486 219218 24570 219454
rect 24806 219218 43930 219454
rect 44166 219218 44250 219454
rect 44486 219218 44570 219454
rect 44806 219218 63930 219454
rect 64166 219218 64250 219454
rect 64486 219218 64570 219454
rect 64806 219218 83930 219454
rect 84166 219218 84250 219454
rect 84486 219218 84570 219454
rect 84806 219218 103930 219454
rect 104166 219218 104250 219454
rect 104486 219218 104570 219454
rect 104806 219218 123930 219454
rect 124166 219218 124250 219454
rect 124486 219218 124570 219454
rect 124806 219218 143930 219454
rect 144166 219218 144250 219454
rect 144486 219218 144570 219454
rect 144806 219218 163930 219454
rect 164166 219218 164250 219454
rect 164486 219218 164570 219454
rect 164806 219218 183930 219454
rect 184166 219218 184250 219454
rect 184486 219218 184570 219454
rect 184806 219218 203930 219454
rect 204166 219218 204250 219454
rect 204486 219218 204570 219454
rect 204806 219218 223930 219454
rect 224166 219218 224250 219454
rect 224486 219218 224570 219454
rect 224806 219218 243930 219454
rect 244166 219218 244250 219454
rect 244486 219218 244570 219454
rect 244806 219218 263930 219454
rect 264166 219218 264250 219454
rect 264486 219218 264570 219454
rect 264806 219218 283930 219454
rect 284166 219218 284250 219454
rect 284486 219218 284570 219454
rect 284806 219218 303930 219454
rect 304166 219218 304250 219454
rect 304486 219218 304570 219454
rect 304806 219218 323930 219454
rect 324166 219218 324250 219454
rect 324486 219218 324570 219454
rect 324806 219218 343930 219454
rect 344166 219218 344250 219454
rect 344486 219218 344570 219454
rect 344806 219218 363930 219454
rect 364166 219218 364250 219454
rect 364486 219218 364570 219454
rect 364806 219218 383930 219454
rect 384166 219218 384250 219454
rect 384486 219218 384570 219454
rect 384806 219218 403930 219454
rect 404166 219218 404250 219454
rect 404486 219218 404570 219454
rect 404806 219218 423930 219454
rect 424166 219218 424250 219454
rect 424486 219218 424570 219454
rect 424806 219218 443930 219454
rect 444166 219218 444250 219454
rect 444486 219218 444570 219454
rect 444806 219218 463930 219454
rect 464166 219218 464250 219454
rect 464486 219218 464570 219454
rect 464806 219218 483930 219454
rect 484166 219218 484250 219454
rect 484486 219218 484570 219454
rect 484806 219218 503930 219454
rect 504166 219218 504250 219454
rect 504486 219218 504570 219454
rect 504806 219218 523930 219454
rect 524166 219218 524250 219454
rect 524486 219218 524570 219454
rect 524806 219218 543930 219454
rect 544166 219218 544250 219454
rect 544486 219218 544570 219454
rect 544806 219218 563930 219454
rect 564166 219218 564250 219454
rect 564486 219218 564570 219454
rect 564806 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 23930 219134
rect 24166 218898 24250 219134
rect 24486 218898 24570 219134
rect 24806 218898 43930 219134
rect 44166 218898 44250 219134
rect 44486 218898 44570 219134
rect 44806 218898 63930 219134
rect 64166 218898 64250 219134
rect 64486 218898 64570 219134
rect 64806 218898 83930 219134
rect 84166 218898 84250 219134
rect 84486 218898 84570 219134
rect 84806 218898 103930 219134
rect 104166 218898 104250 219134
rect 104486 218898 104570 219134
rect 104806 218898 123930 219134
rect 124166 218898 124250 219134
rect 124486 218898 124570 219134
rect 124806 218898 143930 219134
rect 144166 218898 144250 219134
rect 144486 218898 144570 219134
rect 144806 218898 163930 219134
rect 164166 218898 164250 219134
rect 164486 218898 164570 219134
rect 164806 218898 183930 219134
rect 184166 218898 184250 219134
rect 184486 218898 184570 219134
rect 184806 218898 203930 219134
rect 204166 218898 204250 219134
rect 204486 218898 204570 219134
rect 204806 218898 223930 219134
rect 224166 218898 224250 219134
rect 224486 218898 224570 219134
rect 224806 218898 243930 219134
rect 244166 218898 244250 219134
rect 244486 218898 244570 219134
rect 244806 218898 263930 219134
rect 264166 218898 264250 219134
rect 264486 218898 264570 219134
rect 264806 218898 283930 219134
rect 284166 218898 284250 219134
rect 284486 218898 284570 219134
rect 284806 218898 303930 219134
rect 304166 218898 304250 219134
rect 304486 218898 304570 219134
rect 304806 218898 323930 219134
rect 324166 218898 324250 219134
rect 324486 218898 324570 219134
rect 324806 218898 343930 219134
rect 344166 218898 344250 219134
rect 344486 218898 344570 219134
rect 344806 218898 363930 219134
rect 364166 218898 364250 219134
rect 364486 218898 364570 219134
rect 364806 218898 383930 219134
rect 384166 218898 384250 219134
rect 384486 218898 384570 219134
rect 384806 218898 403930 219134
rect 404166 218898 404250 219134
rect 404486 218898 404570 219134
rect 404806 218898 423930 219134
rect 424166 218898 424250 219134
rect 424486 218898 424570 219134
rect 424806 218898 443930 219134
rect 444166 218898 444250 219134
rect 444486 218898 444570 219134
rect 444806 218898 463930 219134
rect 464166 218898 464250 219134
rect 464486 218898 464570 219134
rect 464806 218898 483930 219134
rect 484166 218898 484250 219134
rect 484486 218898 484570 219134
rect 484806 218898 503930 219134
rect 504166 218898 504250 219134
rect 504486 218898 504570 219134
rect 504806 218898 523930 219134
rect 524166 218898 524250 219134
rect 524486 218898 524570 219134
rect 524806 218898 543930 219134
rect 544166 218898 544250 219134
rect 544486 218898 544570 219134
rect 544806 218898 563930 219134
rect 564166 218898 564250 219134
rect 564486 218898 564570 219134
rect 564806 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 23930 183454
rect 24166 183218 24250 183454
rect 24486 183218 24570 183454
rect 24806 183218 43930 183454
rect 44166 183218 44250 183454
rect 44486 183218 44570 183454
rect 44806 183218 63930 183454
rect 64166 183218 64250 183454
rect 64486 183218 64570 183454
rect 64806 183218 83930 183454
rect 84166 183218 84250 183454
rect 84486 183218 84570 183454
rect 84806 183218 103930 183454
rect 104166 183218 104250 183454
rect 104486 183218 104570 183454
rect 104806 183218 123930 183454
rect 124166 183218 124250 183454
rect 124486 183218 124570 183454
rect 124806 183218 143930 183454
rect 144166 183218 144250 183454
rect 144486 183218 144570 183454
rect 144806 183218 163930 183454
rect 164166 183218 164250 183454
rect 164486 183218 164570 183454
rect 164806 183218 183930 183454
rect 184166 183218 184250 183454
rect 184486 183218 184570 183454
rect 184806 183218 203930 183454
rect 204166 183218 204250 183454
rect 204486 183218 204570 183454
rect 204806 183218 223930 183454
rect 224166 183218 224250 183454
rect 224486 183218 224570 183454
rect 224806 183218 243930 183454
rect 244166 183218 244250 183454
rect 244486 183218 244570 183454
rect 244806 183218 263930 183454
rect 264166 183218 264250 183454
rect 264486 183218 264570 183454
rect 264806 183218 283930 183454
rect 284166 183218 284250 183454
rect 284486 183218 284570 183454
rect 284806 183218 303930 183454
rect 304166 183218 304250 183454
rect 304486 183218 304570 183454
rect 304806 183218 323930 183454
rect 324166 183218 324250 183454
rect 324486 183218 324570 183454
rect 324806 183218 343930 183454
rect 344166 183218 344250 183454
rect 344486 183218 344570 183454
rect 344806 183218 363930 183454
rect 364166 183218 364250 183454
rect 364486 183218 364570 183454
rect 364806 183218 383930 183454
rect 384166 183218 384250 183454
rect 384486 183218 384570 183454
rect 384806 183218 403930 183454
rect 404166 183218 404250 183454
rect 404486 183218 404570 183454
rect 404806 183218 423930 183454
rect 424166 183218 424250 183454
rect 424486 183218 424570 183454
rect 424806 183218 443930 183454
rect 444166 183218 444250 183454
rect 444486 183218 444570 183454
rect 444806 183218 463930 183454
rect 464166 183218 464250 183454
rect 464486 183218 464570 183454
rect 464806 183218 483930 183454
rect 484166 183218 484250 183454
rect 484486 183218 484570 183454
rect 484806 183218 503930 183454
rect 504166 183218 504250 183454
rect 504486 183218 504570 183454
rect 504806 183218 523930 183454
rect 524166 183218 524250 183454
rect 524486 183218 524570 183454
rect 524806 183218 543930 183454
rect 544166 183218 544250 183454
rect 544486 183218 544570 183454
rect 544806 183218 563930 183454
rect 564166 183218 564250 183454
rect 564486 183218 564570 183454
rect 564806 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 23930 183134
rect 24166 182898 24250 183134
rect 24486 182898 24570 183134
rect 24806 182898 43930 183134
rect 44166 182898 44250 183134
rect 44486 182898 44570 183134
rect 44806 182898 63930 183134
rect 64166 182898 64250 183134
rect 64486 182898 64570 183134
rect 64806 182898 83930 183134
rect 84166 182898 84250 183134
rect 84486 182898 84570 183134
rect 84806 182898 103930 183134
rect 104166 182898 104250 183134
rect 104486 182898 104570 183134
rect 104806 182898 123930 183134
rect 124166 182898 124250 183134
rect 124486 182898 124570 183134
rect 124806 182898 143930 183134
rect 144166 182898 144250 183134
rect 144486 182898 144570 183134
rect 144806 182898 163930 183134
rect 164166 182898 164250 183134
rect 164486 182898 164570 183134
rect 164806 182898 183930 183134
rect 184166 182898 184250 183134
rect 184486 182898 184570 183134
rect 184806 182898 203930 183134
rect 204166 182898 204250 183134
rect 204486 182898 204570 183134
rect 204806 182898 223930 183134
rect 224166 182898 224250 183134
rect 224486 182898 224570 183134
rect 224806 182898 243930 183134
rect 244166 182898 244250 183134
rect 244486 182898 244570 183134
rect 244806 182898 263930 183134
rect 264166 182898 264250 183134
rect 264486 182898 264570 183134
rect 264806 182898 283930 183134
rect 284166 182898 284250 183134
rect 284486 182898 284570 183134
rect 284806 182898 303930 183134
rect 304166 182898 304250 183134
rect 304486 182898 304570 183134
rect 304806 182898 323930 183134
rect 324166 182898 324250 183134
rect 324486 182898 324570 183134
rect 324806 182898 343930 183134
rect 344166 182898 344250 183134
rect 344486 182898 344570 183134
rect 344806 182898 363930 183134
rect 364166 182898 364250 183134
rect 364486 182898 364570 183134
rect 364806 182898 383930 183134
rect 384166 182898 384250 183134
rect 384486 182898 384570 183134
rect 384806 182898 403930 183134
rect 404166 182898 404250 183134
rect 404486 182898 404570 183134
rect 404806 182898 423930 183134
rect 424166 182898 424250 183134
rect 424486 182898 424570 183134
rect 424806 182898 443930 183134
rect 444166 182898 444250 183134
rect 444486 182898 444570 183134
rect 444806 182898 463930 183134
rect 464166 182898 464250 183134
rect 464486 182898 464570 183134
rect 464806 182898 483930 183134
rect 484166 182898 484250 183134
rect 484486 182898 484570 183134
rect 484806 182898 503930 183134
rect 504166 182898 504250 183134
rect 504486 182898 504570 183134
rect 504806 182898 523930 183134
rect 524166 182898 524250 183134
rect 524486 182898 524570 183134
rect 524806 182898 543930 183134
rect 544166 182898 544250 183134
rect 544486 182898 544570 183134
rect 544806 182898 563930 183134
rect 564166 182898 564250 183134
rect 564486 182898 564570 183134
rect 564806 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 33930 151954
rect 34166 151718 34250 151954
rect 34486 151718 34570 151954
rect 34806 151718 53930 151954
rect 54166 151718 54250 151954
rect 54486 151718 54570 151954
rect 54806 151718 73930 151954
rect 74166 151718 74250 151954
rect 74486 151718 74570 151954
rect 74806 151718 93930 151954
rect 94166 151718 94250 151954
rect 94486 151718 94570 151954
rect 94806 151718 113930 151954
rect 114166 151718 114250 151954
rect 114486 151718 114570 151954
rect 114806 151718 133930 151954
rect 134166 151718 134250 151954
rect 134486 151718 134570 151954
rect 134806 151718 153930 151954
rect 154166 151718 154250 151954
rect 154486 151718 154570 151954
rect 154806 151718 173930 151954
rect 174166 151718 174250 151954
rect 174486 151718 174570 151954
rect 174806 151718 193930 151954
rect 194166 151718 194250 151954
rect 194486 151718 194570 151954
rect 194806 151718 213930 151954
rect 214166 151718 214250 151954
rect 214486 151718 214570 151954
rect 214806 151718 233930 151954
rect 234166 151718 234250 151954
rect 234486 151718 234570 151954
rect 234806 151718 253930 151954
rect 254166 151718 254250 151954
rect 254486 151718 254570 151954
rect 254806 151718 273930 151954
rect 274166 151718 274250 151954
rect 274486 151718 274570 151954
rect 274806 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 313930 151954
rect 314166 151718 314250 151954
rect 314486 151718 314570 151954
rect 314806 151718 333930 151954
rect 334166 151718 334250 151954
rect 334486 151718 334570 151954
rect 334806 151718 353930 151954
rect 354166 151718 354250 151954
rect 354486 151718 354570 151954
rect 354806 151718 373930 151954
rect 374166 151718 374250 151954
rect 374486 151718 374570 151954
rect 374806 151718 393930 151954
rect 394166 151718 394250 151954
rect 394486 151718 394570 151954
rect 394806 151718 413930 151954
rect 414166 151718 414250 151954
rect 414486 151718 414570 151954
rect 414806 151718 433930 151954
rect 434166 151718 434250 151954
rect 434486 151718 434570 151954
rect 434806 151718 453930 151954
rect 454166 151718 454250 151954
rect 454486 151718 454570 151954
rect 454806 151718 473930 151954
rect 474166 151718 474250 151954
rect 474486 151718 474570 151954
rect 474806 151718 493930 151954
rect 494166 151718 494250 151954
rect 494486 151718 494570 151954
rect 494806 151718 513930 151954
rect 514166 151718 514250 151954
rect 514486 151718 514570 151954
rect 514806 151718 533930 151954
rect 534166 151718 534250 151954
rect 534486 151718 534570 151954
rect 534806 151718 553930 151954
rect 554166 151718 554250 151954
rect 554486 151718 554570 151954
rect 554806 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 33930 151634
rect 34166 151398 34250 151634
rect 34486 151398 34570 151634
rect 34806 151398 53930 151634
rect 54166 151398 54250 151634
rect 54486 151398 54570 151634
rect 54806 151398 73930 151634
rect 74166 151398 74250 151634
rect 74486 151398 74570 151634
rect 74806 151398 93930 151634
rect 94166 151398 94250 151634
rect 94486 151398 94570 151634
rect 94806 151398 113930 151634
rect 114166 151398 114250 151634
rect 114486 151398 114570 151634
rect 114806 151398 133930 151634
rect 134166 151398 134250 151634
rect 134486 151398 134570 151634
rect 134806 151398 153930 151634
rect 154166 151398 154250 151634
rect 154486 151398 154570 151634
rect 154806 151398 173930 151634
rect 174166 151398 174250 151634
rect 174486 151398 174570 151634
rect 174806 151398 193930 151634
rect 194166 151398 194250 151634
rect 194486 151398 194570 151634
rect 194806 151398 213930 151634
rect 214166 151398 214250 151634
rect 214486 151398 214570 151634
rect 214806 151398 233930 151634
rect 234166 151398 234250 151634
rect 234486 151398 234570 151634
rect 234806 151398 253930 151634
rect 254166 151398 254250 151634
rect 254486 151398 254570 151634
rect 254806 151398 273930 151634
rect 274166 151398 274250 151634
rect 274486 151398 274570 151634
rect 274806 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 313930 151634
rect 314166 151398 314250 151634
rect 314486 151398 314570 151634
rect 314806 151398 333930 151634
rect 334166 151398 334250 151634
rect 334486 151398 334570 151634
rect 334806 151398 353930 151634
rect 354166 151398 354250 151634
rect 354486 151398 354570 151634
rect 354806 151398 373930 151634
rect 374166 151398 374250 151634
rect 374486 151398 374570 151634
rect 374806 151398 393930 151634
rect 394166 151398 394250 151634
rect 394486 151398 394570 151634
rect 394806 151398 413930 151634
rect 414166 151398 414250 151634
rect 414486 151398 414570 151634
rect 414806 151398 433930 151634
rect 434166 151398 434250 151634
rect 434486 151398 434570 151634
rect 434806 151398 453930 151634
rect 454166 151398 454250 151634
rect 454486 151398 454570 151634
rect 454806 151398 473930 151634
rect 474166 151398 474250 151634
rect 474486 151398 474570 151634
rect 474806 151398 493930 151634
rect 494166 151398 494250 151634
rect 494486 151398 494570 151634
rect 494806 151398 513930 151634
rect 514166 151398 514250 151634
rect 514486 151398 514570 151634
rect 514806 151398 533930 151634
rect 534166 151398 534250 151634
rect 534486 151398 534570 151634
rect 534806 151398 553930 151634
rect 554166 151398 554250 151634
rect 554486 151398 554570 151634
rect 554806 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 23930 147454
rect 24166 147218 24250 147454
rect 24486 147218 24570 147454
rect 24806 147218 43930 147454
rect 44166 147218 44250 147454
rect 44486 147218 44570 147454
rect 44806 147218 63930 147454
rect 64166 147218 64250 147454
rect 64486 147218 64570 147454
rect 64806 147218 83930 147454
rect 84166 147218 84250 147454
rect 84486 147218 84570 147454
rect 84806 147218 103930 147454
rect 104166 147218 104250 147454
rect 104486 147218 104570 147454
rect 104806 147218 123930 147454
rect 124166 147218 124250 147454
rect 124486 147218 124570 147454
rect 124806 147218 143930 147454
rect 144166 147218 144250 147454
rect 144486 147218 144570 147454
rect 144806 147218 163930 147454
rect 164166 147218 164250 147454
rect 164486 147218 164570 147454
rect 164806 147218 183930 147454
rect 184166 147218 184250 147454
rect 184486 147218 184570 147454
rect 184806 147218 203930 147454
rect 204166 147218 204250 147454
rect 204486 147218 204570 147454
rect 204806 147218 223930 147454
rect 224166 147218 224250 147454
rect 224486 147218 224570 147454
rect 224806 147218 243930 147454
rect 244166 147218 244250 147454
rect 244486 147218 244570 147454
rect 244806 147218 263930 147454
rect 264166 147218 264250 147454
rect 264486 147218 264570 147454
rect 264806 147218 283930 147454
rect 284166 147218 284250 147454
rect 284486 147218 284570 147454
rect 284806 147218 303930 147454
rect 304166 147218 304250 147454
rect 304486 147218 304570 147454
rect 304806 147218 323930 147454
rect 324166 147218 324250 147454
rect 324486 147218 324570 147454
rect 324806 147218 343930 147454
rect 344166 147218 344250 147454
rect 344486 147218 344570 147454
rect 344806 147218 363930 147454
rect 364166 147218 364250 147454
rect 364486 147218 364570 147454
rect 364806 147218 383930 147454
rect 384166 147218 384250 147454
rect 384486 147218 384570 147454
rect 384806 147218 403930 147454
rect 404166 147218 404250 147454
rect 404486 147218 404570 147454
rect 404806 147218 423930 147454
rect 424166 147218 424250 147454
rect 424486 147218 424570 147454
rect 424806 147218 443930 147454
rect 444166 147218 444250 147454
rect 444486 147218 444570 147454
rect 444806 147218 463930 147454
rect 464166 147218 464250 147454
rect 464486 147218 464570 147454
rect 464806 147218 483930 147454
rect 484166 147218 484250 147454
rect 484486 147218 484570 147454
rect 484806 147218 503930 147454
rect 504166 147218 504250 147454
rect 504486 147218 504570 147454
rect 504806 147218 523930 147454
rect 524166 147218 524250 147454
rect 524486 147218 524570 147454
rect 524806 147218 543930 147454
rect 544166 147218 544250 147454
rect 544486 147218 544570 147454
rect 544806 147218 563930 147454
rect 564166 147218 564250 147454
rect 564486 147218 564570 147454
rect 564806 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 23930 147134
rect 24166 146898 24250 147134
rect 24486 146898 24570 147134
rect 24806 146898 43930 147134
rect 44166 146898 44250 147134
rect 44486 146898 44570 147134
rect 44806 146898 63930 147134
rect 64166 146898 64250 147134
rect 64486 146898 64570 147134
rect 64806 146898 83930 147134
rect 84166 146898 84250 147134
rect 84486 146898 84570 147134
rect 84806 146898 103930 147134
rect 104166 146898 104250 147134
rect 104486 146898 104570 147134
rect 104806 146898 123930 147134
rect 124166 146898 124250 147134
rect 124486 146898 124570 147134
rect 124806 146898 143930 147134
rect 144166 146898 144250 147134
rect 144486 146898 144570 147134
rect 144806 146898 163930 147134
rect 164166 146898 164250 147134
rect 164486 146898 164570 147134
rect 164806 146898 183930 147134
rect 184166 146898 184250 147134
rect 184486 146898 184570 147134
rect 184806 146898 203930 147134
rect 204166 146898 204250 147134
rect 204486 146898 204570 147134
rect 204806 146898 223930 147134
rect 224166 146898 224250 147134
rect 224486 146898 224570 147134
rect 224806 146898 243930 147134
rect 244166 146898 244250 147134
rect 244486 146898 244570 147134
rect 244806 146898 263930 147134
rect 264166 146898 264250 147134
rect 264486 146898 264570 147134
rect 264806 146898 283930 147134
rect 284166 146898 284250 147134
rect 284486 146898 284570 147134
rect 284806 146898 303930 147134
rect 304166 146898 304250 147134
rect 304486 146898 304570 147134
rect 304806 146898 323930 147134
rect 324166 146898 324250 147134
rect 324486 146898 324570 147134
rect 324806 146898 343930 147134
rect 344166 146898 344250 147134
rect 344486 146898 344570 147134
rect 344806 146898 363930 147134
rect 364166 146898 364250 147134
rect 364486 146898 364570 147134
rect 364806 146898 383930 147134
rect 384166 146898 384250 147134
rect 384486 146898 384570 147134
rect 384806 146898 403930 147134
rect 404166 146898 404250 147134
rect 404486 146898 404570 147134
rect 404806 146898 423930 147134
rect 424166 146898 424250 147134
rect 424486 146898 424570 147134
rect 424806 146898 443930 147134
rect 444166 146898 444250 147134
rect 444486 146898 444570 147134
rect 444806 146898 463930 147134
rect 464166 146898 464250 147134
rect 464486 146898 464570 147134
rect 464806 146898 483930 147134
rect 484166 146898 484250 147134
rect 484486 146898 484570 147134
rect 484806 146898 503930 147134
rect 504166 146898 504250 147134
rect 504486 146898 504570 147134
rect 504806 146898 523930 147134
rect 524166 146898 524250 147134
rect 524486 146898 524570 147134
rect 524806 146898 543930 147134
rect 544166 146898 544250 147134
rect 544486 146898 544570 147134
rect 544806 146898 563930 147134
rect 564166 146898 564250 147134
rect 564486 146898 564570 147134
rect 564806 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 33930 115954
rect 34166 115718 34250 115954
rect 34486 115718 34570 115954
rect 34806 115718 53930 115954
rect 54166 115718 54250 115954
rect 54486 115718 54570 115954
rect 54806 115718 73930 115954
rect 74166 115718 74250 115954
rect 74486 115718 74570 115954
rect 74806 115718 93930 115954
rect 94166 115718 94250 115954
rect 94486 115718 94570 115954
rect 94806 115718 113930 115954
rect 114166 115718 114250 115954
rect 114486 115718 114570 115954
rect 114806 115718 133930 115954
rect 134166 115718 134250 115954
rect 134486 115718 134570 115954
rect 134806 115718 153930 115954
rect 154166 115718 154250 115954
rect 154486 115718 154570 115954
rect 154806 115718 173930 115954
rect 174166 115718 174250 115954
rect 174486 115718 174570 115954
rect 174806 115718 193930 115954
rect 194166 115718 194250 115954
rect 194486 115718 194570 115954
rect 194806 115718 213930 115954
rect 214166 115718 214250 115954
rect 214486 115718 214570 115954
rect 214806 115718 233930 115954
rect 234166 115718 234250 115954
rect 234486 115718 234570 115954
rect 234806 115718 253930 115954
rect 254166 115718 254250 115954
rect 254486 115718 254570 115954
rect 254806 115718 273930 115954
rect 274166 115718 274250 115954
rect 274486 115718 274570 115954
rect 274806 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 313930 115954
rect 314166 115718 314250 115954
rect 314486 115718 314570 115954
rect 314806 115718 333930 115954
rect 334166 115718 334250 115954
rect 334486 115718 334570 115954
rect 334806 115718 353930 115954
rect 354166 115718 354250 115954
rect 354486 115718 354570 115954
rect 354806 115718 373930 115954
rect 374166 115718 374250 115954
rect 374486 115718 374570 115954
rect 374806 115718 393930 115954
rect 394166 115718 394250 115954
rect 394486 115718 394570 115954
rect 394806 115718 413930 115954
rect 414166 115718 414250 115954
rect 414486 115718 414570 115954
rect 414806 115718 433930 115954
rect 434166 115718 434250 115954
rect 434486 115718 434570 115954
rect 434806 115718 453930 115954
rect 454166 115718 454250 115954
rect 454486 115718 454570 115954
rect 454806 115718 473930 115954
rect 474166 115718 474250 115954
rect 474486 115718 474570 115954
rect 474806 115718 493930 115954
rect 494166 115718 494250 115954
rect 494486 115718 494570 115954
rect 494806 115718 513930 115954
rect 514166 115718 514250 115954
rect 514486 115718 514570 115954
rect 514806 115718 533930 115954
rect 534166 115718 534250 115954
rect 534486 115718 534570 115954
rect 534806 115718 553930 115954
rect 554166 115718 554250 115954
rect 554486 115718 554570 115954
rect 554806 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 33930 115634
rect 34166 115398 34250 115634
rect 34486 115398 34570 115634
rect 34806 115398 53930 115634
rect 54166 115398 54250 115634
rect 54486 115398 54570 115634
rect 54806 115398 73930 115634
rect 74166 115398 74250 115634
rect 74486 115398 74570 115634
rect 74806 115398 93930 115634
rect 94166 115398 94250 115634
rect 94486 115398 94570 115634
rect 94806 115398 113930 115634
rect 114166 115398 114250 115634
rect 114486 115398 114570 115634
rect 114806 115398 133930 115634
rect 134166 115398 134250 115634
rect 134486 115398 134570 115634
rect 134806 115398 153930 115634
rect 154166 115398 154250 115634
rect 154486 115398 154570 115634
rect 154806 115398 173930 115634
rect 174166 115398 174250 115634
rect 174486 115398 174570 115634
rect 174806 115398 193930 115634
rect 194166 115398 194250 115634
rect 194486 115398 194570 115634
rect 194806 115398 213930 115634
rect 214166 115398 214250 115634
rect 214486 115398 214570 115634
rect 214806 115398 233930 115634
rect 234166 115398 234250 115634
rect 234486 115398 234570 115634
rect 234806 115398 253930 115634
rect 254166 115398 254250 115634
rect 254486 115398 254570 115634
rect 254806 115398 273930 115634
rect 274166 115398 274250 115634
rect 274486 115398 274570 115634
rect 274806 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 313930 115634
rect 314166 115398 314250 115634
rect 314486 115398 314570 115634
rect 314806 115398 333930 115634
rect 334166 115398 334250 115634
rect 334486 115398 334570 115634
rect 334806 115398 353930 115634
rect 354166 115398 354250 115634
rect 354486 115398 354570 115634
rect 354806 115398 373930 115634
rect 374166 115398 374250 115634
rect 374486 115398 374570 115634
rect 374806 115398 393930 115634
rect 394166 115398 394250 115634
rect 394486 115398 394570 115634
rect 394806 115398 413930 115634
rect 414166 115398 414250 115634
rect 414486 115398 414570 115634
rect 414806 115398 433930 115634
rect 434166 115398 434250 115634
rect 434486 115398 434570 115634
rect 434806 115398 453930 115634
rect 454166 115398 454250 115634
rect 454486 115398 454570 115634
rect 454806 115398 473930 115634
rect 474166 115398 474250 115634
rect 474486 115398 474570 115634
rect 474806 115398 493930 115634
rect 494166 115398 494250 115634
rect 494486 115398 494570 115634
rect 494806 115398 513930 115634
rect 514166 115398 514250 115634
rect 514486 115398 514570 115634
rect 514806 115398 533930 115634
rect 534166 115398 534250 115634
rect 534486 115398 534570 115634
rect 534806 115398 553930 115634
rect 554166 115398 554250 115634
rect 554486 115398 554570 115634
rect 554806 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 23930 111454
rect 24166 111218 24250 111454
rect 24486 111218 24570 111454
rect 24806 111218 43930 111454
rect 44166 111218 44250 111454
rect 44486 111218 44570 111454
rect 44806 111218 63930 111454
rect 64166 111218 64250 111454
rect 64486 111218 64570 111454
rect 64806 111218 83930 111454
rect 84166 111218 84250 111454
rect 84486 111218 84570 111454
rect 84806 111218 103930 111454
rect 104166 111218 104250 111454
rect 104486 111218 104570 111454
rect 104806 111218 123930 111454
rect 124166 111218 124250 111454
rect 124486 111218 124570 111454
rect 124806 111218 143930 111454
rect 144166 111218 144250 111454
rect 144486 111218 144570 111454
rect 144806 111218 163930 111454
rect 164166 111218 164250 111454
rect 164486 111218 164570 111454
rect 164806 111218 183930 111454
rect 184166 111218 184250 111454
rect 184486 111218 184570 111454
rect 184806 111218 203930 111454
rect 204166 111218 204250 111454
rect 204486 111218 204570 111454
rect 204806 111218 223930 111454
rect 224166 111218 224250 111454
rect 224486 111218 224570 111454
rect 224806 111218 243930 111454
rect 244166 111218 244250 111454
rect 244486 111218 244570 111454
rect 244806 111218 263930 111454
rect 264166 111218 264250 111454
rect 264486 111218 264570 111454
rect 264806 111218 283930 111454
rect 284166 111218 284250 111454
rect 284486 111218 284570 111454
rect 284806 111218 303930 111454
rect 304166 111218 304250 111454
rect 304486 111218 304570 111454
rect 304806 111218 323930 111454
rect 324166 111218 324250 111454
rect 324486 111218 324570 111454
rect 324806 111218 343930 111454
rect 344166 111218 344250 111454
rect 344486 111218 344570 111454
rect 344806 111218 363930 111454
rect 364166 111218 364250 111454
rect 364486 111218 364570 111454
rect 364806 111218 383930 111454
rect 384166 111218 384250 111454
rect 384486 111218 384570 111454
rect 384806 111218 403930 111454
rect 404166 111218 404250 111454
rect 404486 111218 404570 111454
rect 404806 111218 423930 111454
rect 424166 111218 424250 111454
rect 424486 111218 424570 111454
rect 424806 111218 443930 111454
rect 444166 111218 444250 111454
rect 444486 111218 444570 111454
rect 444806 111218 463930 111454
rect 464166 111218 464250 111454
rect 464486 111218 464570 111454
rect 464806 111218 483930 111454
rect 484166 111218 484250 111454
rect 484486 111218 484570 111454
rect 484806 111218 503930 111454
rect 504166 111218 504250 111454
rect 504486 111218 504570 111454
rect 504806 111218 523930 111454
rect 524166 111218 524250 111454
rect 524486 111218 524570 111454
rect 524806 111218 543930 111454
rect 544166 111218 544250 111454
rect 544486 111218 544570 111454
rect 544806 111218 563930 111454
rect 564166 111218 564250 111454
rect 564486 111218 564570 111454
rect 564806 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 23930 111134
rect 24166 110898 24250 111134
rect 24486 110898 24570 111134
rect 24806 110898 43930 111134
rect 44166 110898 44250 111134
rect 44486 110898 44570 111134
rect 44806 110898 63930 111134
rect 64166 110898 64250 111134
rect 64486 110898 64570 111134
rect 64806 110898 83930 111134
rect 84166 110898 84250 111134
rect 84486 110898 84570 111134
rect 84806 110898 103930 111134
rect 104166 110898 104250 111134
rect 104486 110898 104570 111134
rect 104806 110898 123930 111134
rect 124166 110898 124250 111134
rect 124486 110898 124570 111134
rect 124806 110898 143930 111134
rect 144166 110898 144250 111134
rect 144486 110898 144570 111134
rect 144806 110898 163930 111134
rect 164166 110898 164250 111134
rect 164486 110898 164570 111134
rect 164806 110898 183930 111134
rect 184166 110898 184250 111134
rect 184486 110898 184570 111134
rect 184806 110898 203930 111134
rect 204166 110898 204250 111134
rect 204486 110898 204570 111134
rect 204806 110898 223930 111134
rect 224166 110898 224250 111134
rect 224486 110898 224570 111134
rect 224806 110898 243930 111134
rect 244166 110898 244250 111134
rect 244486 110898 244570 111134
rect 244806 110898 263930 111134
rect 264166 110898 264250 111134
rect 264486 110898 264570 111134
rect 264806 110898 283930 111134
rect 284166 110898 284250 111134
rect 284486 110898 284570 111134
rect 284806 110898 303930 111134
rect 304166 110898 304250 111134
rect 304486 110898 304570 111134
rect 304806 110898 323930 111134
rect 324166 110898 324250 111134
rect 324486 110898 324570 111134
rect 324806 110898 343930 111134
rect 344166 110898 344250 111134
rect 344486 110898 344570 111134
rect 344806 110898 363930 111134
rect 364166 110898 364250 111134
rect 364486 110898 364570 111134
rect 364806 110898 383930 111134
rect 384166 110898 384250 111134
rect 384486 110898 384570 111134
rect 384806 110898 403930 111134
rect 404166 110898 404250 111134
rect 404486 110898 404570 111134
rect 404806 110898 423930 111134
rect 424166 110898 424250 111134
rect 424486 110898 424570 111134
rect 424806 110898 443930 111134
rect 444166 110898 444250 111134
rect 444486 110898 444570 111134
rect 444806 110898 463930 111134
rect 464166 110898 464250 111134
rect 464486 110898 464570 111134
rect 464806 110898 483930 111134
rect 484166 110898 484250 111134
rect 484486 110898 484570 111134
rect 484806 110898 503930 111134
rect 504166 110898 504250 111134
rect 504486 110898 504570 111134
rect 504806 110898 523930 111134
rect 524166 110898 524250 111134
rect 524486 110898 524570 111134
rect 524806 110898 543930 111134
rect 544166 110898 544250 111134
rect 544486 110898 544570 111134
rect 544806 110898 563930 111134
rect 564166 110898 564250 111134
rect 564486 110898 564570 111134
rect 564806 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 79610 43954
rect 79846 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 213930 43954
rect 214166 43718 214250 43954
rect 214486 43718 214570 43954
rect 214806 43718 233930 43954
rect 234166 43718 234250 43954
rect 234486 43718 234570 43954
rect 234806 43718 253930 43954
rect 254166 43718 254250 43954
rect 254486 43718 254570 43954
rect 254806 43718 273930 43954
rect 274166 43718 274250 43954
rect 274486 43718 274570 43954
rect 274806 43718 293930 43954
rect 294166 43718 294250 43954
rect 294486 43718 294570 43954
rect 294806 43718 313930 43954
rect 314166 43718 314250 43954
rect 314486 43718 314570 43954
rect 314806 43718 333930 43954
rect 334166 43718 334250 43954
rect 334486 43718 334570 43954
rect 334806 43718 353930 43954
rect 354166 43718 354250 43954
rect 354486 43718 354570 43954
rect 354806 43718 373930 43954
rect 374166 43718 374250 43954
rect 374486 43718 374570 43954
rect 374806 43718 393930 43954
rect 394166 43718 394250 43954
rect 394486 43718 394570 43954
rect 394806 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 79610 43634
rect 79846 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 213930 43634
rect 214166 43398 214250 43634
rect 214486 43398 214570 43634
rect 214806 43398 233930 43634
rect 234166 43398 234250 43634
rect 234486 43398 234570 43634
rect 234806 43398 253930 43634
rect 254166 43398 254250 43634
rect 254486 43398 254570 43634
rect 254806 43398 273930 43634
rect 274166 43398 274250 43634
rect 274486 43398 274570 43634
rect 274806 43398 293930 43634
rect 294166 43398 294250 43634
rect 294486 43398 294570 43634
rect 294806 43398 313930 43634
rect 314166 43398 314250 43634
rect 314486 43398 314570 43634
rect 314806 43398 333930 43634
rect 334166 43398 334250 43634
rect 334486 43398 334570 43634
rect 334806 43398 353930 43634
rect 354166 43398 354250 43634
rect 354486 43398 354570 43634
rect 354806 43398 373930 43634
rect 374166 43398 374250 43634
rect 374486 43398 374570 43634
rect 374806 43398 393930 43634
rect 394166 43398 394250 43634
rect 394486 43398 394570 43634
rect 394806 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 64250 39454
rect 64486 39218 94970 39454
rect 95206 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 203930 39454
rect 204166 39218 204250 39454
rect 204486 39218 204570 39454
rect 204806 39218 223930 39454
rect 224166 39218 224250 39454
rect 224486 39218 224570 39454
rect 224806 39218 243930 39454
rect 244166 39218 244250 39454
rect 244486 39218 244570 39454
rect 244806 39218 263930 39454
rect 264166 39218 264250 39454
rect 264486 39218 264570 39454
rect 264806 39218 283930 39454
rect 284166 39218 284250 39454
rect 284486 39218 284570 39454
rect 284806 39218 303930 39454
rect 304166 39218 304250 39454
rect 304486 39218 304570 39454
rect 304806 39218 323930 39454
rect 324166 39218 324250 39454
rect 324486 39218 324570 39454
rect 324806 39218 343930 39454
rect 344166 39218 344250 39454
rect 344486 39218 344570 39454
rect 344806 39218 363930 39454
rect 364166 39218 364250 39454
rect 364486 39218 364570 39454
rect 364806 39218 383930 39454
rect 384166 39218 384250 39454
rect 384486 39218 384570 39454
rect 384806 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 64250 39134
rect 64486 38898 94970 39134
rect 95206 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 203930 39134
rect 204166 38898 204250 39134
rect 204486 38898 204570 39134
rect 204806 38898 223930 39134
rect 224166 38898 224250 39134
rect 224486 38898 224570 39134
rect 224806 38898 243930 39134
rect 244166 38898 244250 39134
rect 244486 38898 244570 39134
rect 244806 38898 263930 39134
rect 264166 38898 264250 39134
rect 264486 38898 264570 39134
rect 264806 38898 283930 39134
rect 284166 38898 284250 39134
rect 284486 38898 284570 39134
rect 284806 38898 303930 39134
rect 304166 38898 304250 39134
rect 304486 38898 304570 39134
rect 304806 38898 323930 39134
rect 324166 38898 324250 39134
rect 324486 38898 324570 39134
rect 324806 38898 343930 39134
rect 344166 38898 344250 39134
rect 344486 38898 344570 39134
rect 344806 38898 363930 39134
rect 364166 38898 364250 39134
rect 364486 38898 364570 39134
rect 364806 38898 383930 39134
rect 384166 38898 384250 39134
rect 384486 38898 384570 39134
rect 384806 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use controller_core  controller_core_mod
timestamp 0
transform 1 0 200000 0 1 24000
box -800 -800 198812 30800
use driver_core  driver_core_0
timestamp 0
transform 1 0 20000 0 1 78000
box 1066 -800 268862 107760
use driver_core  driver_core_1
timestamp 0
transform 1 0 20000 0 1 206000
box 1066 -800 268862 107760
use driver_core  driver_core_2
timestamp 0
transform 1 0 20000 0 1 334000
box 1066 -800 268862 107760
use driver_core  driver_core_3
timestamp 0
transform 1 0 20000 0 1 462000
box 1066 -800 268862 107760
use driver_core  driver_core_4
timestamp 0
transform 1 0 20000 0 1 588000
box 1066 -800 268862 107760
use driver_core  driver_core_5
timestamp 0
transform 1 0 300000 0 1 588000
box 1066 -800 268862 107760
use driver_core  driver_core_6
timestamp 0
transform 1 0 300000 0 1 462000
box 1066 -800 268862 107760
use driver_core  driver_core_7
timestamp 0
transform 1 0 300000 0 1 334000
box 1066 -800 268862 107760
use driver_core  driver_core_8
timestamp 0
transform 1 0 300000 0 1 206000
box 1066 -800 268862 107760
use driver_core  driver_core_9
timestamp 0
transform 1 0 300000 0 1 78000
box 1066 -800 268862 107760
use spi_controller  spi_controller_mod
timestamp 0
transform 1 0 60000 0 1 24000
box 0 0 40000 37584
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 22000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 22000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 22000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 56000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 22000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 700000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 700000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 700000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 700000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 700000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 700000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 700000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 700000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 700000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 22000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 700000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 700000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 700000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 700000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 700000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 700000 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
