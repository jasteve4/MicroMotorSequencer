VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO driver_core
  CLASS BLOCK ;
  FOREIGN driver_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1350.000 BY 550.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 -4.000 573.530 4.000 ;
    END
  END clock
  PIN clock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 -4.000 544.550 4.000 ;
    END
  END clock_a
  PIN col_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 -4.000 1095.170 4.000 ;
    END
  END col_select_a[0]
  PIN col_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 -4.000 1124.150 4.000 ;
    END
  END col_select_a[1]
  PIN col_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 -4.000 1153.130 4.000 ;
    END
  END col_select_a[2]
  PIN col_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 -4.000 1182.110 4.000 ;
    END
  END col_select_a[3]
  PIN col_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 -4.000 1211.090 4.000 ;
    END
  END col_select_a[4]
  PIN col_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 -4.000 1240.070 4.000 ;
    END
  END col_select_a[5]
  PIN data_in_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END data_in_a[0]
  PIN data_in_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 -4.000 370.670 4.000 ;
    END
  END data_in_a[10]
  PIN data_in_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 -4.000 399.650 4.000 ;
    END
  END data_in_a[11]
  PIN data_in_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 -4.000 428.630 4.000 ;
    END
  END data_in_a[12]
  PIN data_in_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 -4.000 457.610 4.000 ;
    END
  END data_in_a[13]
  PIN data_in_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 -4.000 486.590 4.000 ;
    END
  END data_in_a[14]
  PIN data_in_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 -4.000 515.570 4.000 ;
    END
  END data_in_a[15]
  PIN data_in_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 -4.000 109.850 4.000 ;
    END
  END data_in_a[1]
  PIN data_in_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 -4.000 138.830 4.000 ;
    END
  END data_in_a[2]
  PIN data_in_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 -4.000 167.810 4.000 ;
    END
  END data_in_a[3]
  PIN data_in_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 -4.000 196.790 4.000 ;
    END
  END data_in_a[4]
  PIN data_in_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 -4.000 225.770 4.000 ;
    END
  END data_in_a[5]
  PIN data_in_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 -4.000 254.750 4.000 ;
    END
  END data_in_a[6]
  PIN data_in_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 -4.000 283.730 4.000 ;
    END
  END data_in_a[7]
  PIN data_in_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -4.000 312.710 4.000 ;
    END
  END data_in_a[8]
  PIN data_in_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 -4.000 341.690 4.000 ;
    END
  END data_in_a[9]
  PIN driver_io[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 -4.000 22.910 4.000 ;
    END
  END driver_io[0]
  PIN driver_io[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 -4.000 51.890 4.000 ;
    END
  END driver_io[1]
  PIN inverter_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 -4.000 1327.010 4.000 ;
    END
  END inverter_select_a
  PIN mem_address_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 -4.000 602.510 4.000 ;
    END
  END mem_address_a[0]
  PIN mem_address_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 -4.000 631.490 4.000 ;
    END
  END mem_address_a[1]
  PIN mem_address_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 -4.000 660.470 4.000 ;
    END
  END mem_address_a[2]
  PIN mem_address_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 -4.000 689.450 4.000 ;
    END
  END mem_address_a[3]
  PIN mem_address_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 -4.000 718.430 4.000 ;
    END
  END mem_address_a[4]
  PIN mem_address_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 -4.000 747.410 4.000 ;
    END
  END mem_address_a[5]
  PIN mem_address_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 -4.000 776.390 4.000 ;
    END
  END mem_address_a[6]
  PIN mem_address_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 -4.000 805.370 4.000 ;
    END
  END mem_address_a[7]
  PIN mem_address_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 -4.000 834.350 4.000 ;
    END
  END mem_address_a[8]
  PIN mem_address_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 -4.000 863.330 4.000 ;
    END
  END mem_address_a[9]
  PIN mem_write_n_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 -4.000 892.310 4.000 ;
    END
  END mem_write_n_a
  PIN output_active_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 -4.000 1298.030 4.000 ;
    END
  END output_active_a
  PIN row_col_select_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 -4.000 1269.050 4.000 ;
    END
  END row_col_select_a
  PIN row_select_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 -4.000 921.290 4.000 ;
    END
  END row_select_a[0]
  PIN row_select_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 -4.000 950.270 4.000 ;
    END
  END row_select_a[1]
  PIN row_select_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 -4.000 979.250 4.000 ;
    END
  END row_select_a[2]
  PIN row_select_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 -4.000 1008.230 4.000 ;
    END
  END row_select_a[3]
  PIN row_select_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 -4.000 1037.210 4.000 ;
    END
  END row_select_a[4]
  PIN row_select_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 -4.000 1066.190 4.000 ;
    END
  END row_select_a[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.340 10.640 24.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.340 10.640 124.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.340 10.640 224.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.340 10.640 324.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.340 10.640 424.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 519.340 10.640 524.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.340 10.640 624.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.340 10.640 724.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.340 10.640 824.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 919.340 10.640 924.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.340 10.640 1024.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1119.340 10.640 1124.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1219.340 10.640 1224.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1319.340 10.640 1324.340 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 69.340 10.640 74.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.340 10.640 174.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.340 10.640 274.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.340 10.640 374.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.340 10.640 474.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.340 10.640 574.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 669.340 10.640 674.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 769.340 10.640 774.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 869.340 10.640 874.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 969.340 10.640 974.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1069.340 10.640 1074.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1169.340 10.640 1174.340 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.340 10.640 1274.340 538.800 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 534.425 1344.310 537.255 ;
        RECT 5.330 528.985 1344.310 531.815 ;
        RECT 5.330 523.545 1344.310 526.375 ;
        RECT 5.330 518.105 1344.310 520.935 ;
        RECT 5.330 512.665 1344.310 515.495 ;
        RECT 5.330 507.225 1344.310 510.055 ;
        RECT 5.330 501.785 1344.310 504.615 ;
        RECT 5.330 496.345 1344.310 499.175 ;
        RECT 5.330 490.905 1344.310 493.735 ;
        RECT 5.330 485.465 1344.310 488.295 ;
        RECT 5.330 480.025 1344.310 482.855 ;
        RECT 5.330 474.585 1344.310 477.415 ;
        RECT 5.330 469.145 1344.310 471.975 ;
        RECT 5.330 463.705 1344.310 466.535 ;
        RECT 5.330 458.265 1344.310 461.095 ;
        RECT 5.330 452.825 1344.310 455.655 ;
        RECT 5.330 447.385 1344.310 450.215 ;
        RECT 5.330 441.945 1344.310 444.775 ;
        RECT 5.330 436.505 1344.310 439.335 ;
        RECT 5.330 431.065 1344.310 433.895 ;
        RECT 5.330 425.625 1344.310 428.455 ;
        RECT 5.330 420.185 1344.310 423.015 ;
        RECT 5.330 414.745 1344.310 417.575 ;
        RECT 5.330 409.305 1344.310 412.135 ;
        RECT 5.330 403.865 1344.310 406.695 ;
        RECT 5.330 398.425 1344.310 401.255 ;
        RECT 5.330 392.985 1344.310 395.815 ;
        RECT 5.330 387.545 1344.310 390.375 ;
        RECT 5.330 382.105 1344.310 384.935 ;
        RECT 5.330 376.665 1344.310 379.495 ;
        RECT 5.330 371.225 1344.310 374.055 ;
        RECT 5.330 365.785 1344.310 368.615 ;
        RECT 5.330 360.345 1344.310 363.175 ;
        RECT 5.330 354.905 1344.310 357.735 ;
        RECT 5.330 349.465 1344.310 352.295 ;
        RECT 5.330 344.025 1344.310 346.855 ;
        RECT 5.330 338.585 1344.310 341.415 ;
        RECT 5.330 333.145 1344.310 335.975 ;
        RECT 5.330 327.705 1344.310 330.535 ;
        RECT 5.330 322.265 1344.310 325.095 ;
        RECT 5.330 316.825 1344.310 319.655 ;
        RECT 5.330 311.385 1344.310 314.215 ;
        RECT 5.330 305.945 1344.310 308.775 ;
        RECT 5.330 300.505 1344.310 303.335 ;
        RECT 5.330 295.065 1344.310 297.895 ;
        RECT 5.330 289.625 1344.310 292.455 ;
        RECT 5.330 284.185 1344.310 287.015 ;
        RECT 5.330 278.745 1344.310 281.575 ;
        RECT 5.330 273.305 1344.310 276.135 ;
        RECT 5.330 267.865 1344.310 270.695 ;
        RECT 5.330 262.425 1344.310 265.255 ;
        RECT 5.330 256.985 1344.310 259.815 ;
        RECT 5.330 251.545 1344.310 254.375 ;
        RECT 5.330 246.105 1344.310 248.935 ;
        RECT 5.330 240.665 1344.310 243.495 ;
        RECT 5.330 235.225 1344.310 238.055 ;
        RECT 5.330 229.785 1344.310 232.615 ;
        RECT 5.330 224.345 1344.310 227.175 ;
        RECT 5.330 218.905 1344.310 221.735 ;
        RECT 5.330 213.465 1344.310 216.295 ;
        RECT 5.330 208.025 1344.310 210.855 ;
        RECT 5.330 202.585 1344.310 205.415 ;
        RECT 5.330 197.145 1344.310 199.975 ;
        RECT 5.330 191.705 1344.310 194.535 ;
        RECT 5.330 186.265 1344.310 189.095 ;
        RECT 5.330 180.825 1344.310 183.655 ;
        RECT 5.330 175.385 1344.310 178.215 ;
        RECT 5.330 169.945 1344.310 172.775 ;
        RECT 5.330 164.505 1344.310 167.335 ;
        RECT 5.330 159.065 1344.310 161.895 ;
        RECT 5.330 153.625 1344.310 156.455 ;
        RECT 5.330 148.185 1344.310 151.015 ;
        RECT 5.330 142.745 1344.310 145.575 ;
        RECT 5.330 137.305 1344.310 140.135 ;
        RECT 5.330 131.865 1344.310 134.695 ;
        RECT 5.330 126.425 1344.310 129.255 ;
        RECT 5.330 120.985 1344.310 123.815 ;
        RECT 5.330 115.545 1344.310 118.375 ;
        RECT 5.330 110.105 1344.310 112.935 ;
        RECT 5.330 104.665 1344.310 107.495 ;
        RECT 5.330 99.225 1344.310 102.055 ;
        RECT 5.330 93.785 1344.310 96.615 ;
        RECT 5.330 88.345 1344.310 91.175 ;
        RECT 5.330 82.905 1344.310 85.735 ;
        RECT 5.330 77.465 1344.310 80.295 ;
        RECT 5.330 72.025 1344.310 74.855 ;
        RECT 5.330 66.585 1344.310 69.415 ;
        RECT 5.330 61.145 1344.310 63.975 ;
        RECT 5.330 55.705 1344.310 58.535 ;
        RECT 5.330 50.265 1344.310 53.095 ;
        RECT 5.330 44.825 1344.310 47.655 ;
        RECT 5.330 39.385 1344.310 42.215 ;
        RECT 5.330 33.945 1344.310 36.775 ;
        RECT 5.330 28.505 1344.310 31.335 ;
        RECT 5.330 23.065 1344.310 25.895 ;
        RECT 5.330 17.625 1344.310 20.455 ;
        RECT 5.330 12.185 1344.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1344.120 538.645 ;
      LAYER met1 ;
        RECT 5.520 7.520 1344.120 538.800 ;
      LAYER met2 ;
        RECT 19.470 4.280 1329.300 538.745 ;
        RECT 19.470 3.670 22.350 4.280 ;
        RECT 23.190 3.670 51.330 4.280 ;
        RECT 52.170 3.670 80.310 4.280 ;
        RECT 81.150 3.670 109.290 4.280 ;
        RECT 110.130 3.670 138.270 4.280 ;
        RECT 139.110 3.670 167.250 4.280 ;
        RECT 168.090 3.670 196.230 4.280 ;
        RECT 197.070 3.670 225.210 4.280 ;
        RECT 226.050 3.670 254.190 4.280 ;
        RECT 255.030 3.670 283.170 4.280 ;
        RECT 284.010 3.670 312.150 4.280 ;
        RECT 312.990 3.670 341.130 4.280 ;
        RECT 341.970 3.670 370.110 4.280 ;
        RECT 370.950 3.670 399.090 4.280 ;
        RECT 399.930 3.670 428.070 4.280 ;
        RECT 428.910 3.670 457.050 4.280 ;
        RECT 457.890 3.670 486.030 4.280 ;
        RECT 486.870 3.670 515.010 4.280 ;
        RECT 515.850 3.670 543.990 4.280 ;
        RECT 544.830 3.670 572.970 4.280 ;
        RECT 573.810 3.670 601.950 4.280 ;
        RECT 602.790 3.670 630.930 4.280 ;
        RECT 631.770 3.670 659.910 4.280 ;
        RECT 660.750 3.670 688.890 4.280 ;
        RECT 689.730 3.670 717.870 4.280 ;
        RECT 718.710 3.670 746.850 4.280 ;
        RECT 747.690 3.670 775.830 4.280 ;
        RECT 776.670 3.670 804.810 4.280 ;
        RECT 805.650 3.670 833.790 4.280 ;
        RECT 834.630 3.670 862.770 4.280 ;
        RECT 863.610 3.670 891.750 4.280 ;
        RECT 892.590 3.670 920.730 4.280 ;
        RECT 921.570 3.670 949.710 4.280 ;
        RECT 950.550 3.670 978.690 4.280 ;
        RECT 979.530 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1036.650 4.280 ;
        RECT 1037.490 3.670 1065.630 4.280 ;
        RECT 1066.470 3.670 1094.610 4.280 ;
        RECT 1095.450 3.670 1123.590 4.280 ;
        RECT 1124.430 3.670 1152.570 4.280 ;
        RECT 1153.410 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1210.530 4.280 ;
        RECT 1211.370 3.670 1239.510 4.280 ;
        RECT 1240.350 3.670 1268.490 4.280 ;
        RECT 1269.330 3.670 1297.470 4.280 ;
        RECT 1298.310 3.670 1326.450 4.280 ;
        RECT 1327.290 3.670 1329.300 4.280 ;
      LAYER met3 ;
        RECT 19.450 8.335 1328.415 538.725 ;
      LAYER met4 ;
        RECT 562.415 14.455 568.940 282.025 ;
        RECT 574.740 14.455 618.940 282.025 ;
        RECT 624.740 14.455 668.940 282.025 ;
        RECT 674.740 14.455 718.940 282.025 ;
        RECT 724.740 14.455 768.940 282.025 ;
        RECT 774.740 14.455 818.940 282.025 ;
        RECT 824.740 14.455 868.940 282.025 ;
        RECT 874.740 14.455 918.940 282.025 ;
        RECT 924.740 14.455 968.940 282.025 ;
        RECT 974.740 14.455 1018.940 282.025 ;
        RECT 1024.740 14.455 1068.940 282.025 ;
        RECT 1074.740 14.455 1118.425 282.025 ;
  END
END driver_core
END LIBRARY

